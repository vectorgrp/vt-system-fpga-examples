��/  !5ц��Fc=���F�jgg�.!l=l%!�uN��S^�6�)�Kgn���H8�`�BH��RXMTl#�4N�3����;p�)o���;�Xu^�V"΍I%���V���G��!��g� ����A=������4��Ó;
����6F{į��0Ѵu�;o��g�-ͨ́!	=�dMz��p��q�� � 2��#�D�1�)�RB�p�bg3;�}�a�=D/])�t<��QTӂ7B�ܙ�NC�����;����B��3O�G]��(x�Ng
����������x3�X�����_qz���9��@�G 3�������FeS��h�I/�N����(z�����{�''���Z��b\g��j�;�,��� \��+2��N��F�T+�iK��W.1��M��П/��q��ѻ&��Q��I�B���ɮ����G~Y���	���Y���/7�P��E�I%n/��N��@���	�
b��uc��=�n5�f���;��kk�����@�Z�t��['.>8���^�r�UsT�m��|B�ƅ�W�9�i��E<�Bnwo4�**´�:�mw��?d�gom�ud�LS:�r�n�%�J�2���H#>���)�A�շ�caE��:���q��i�CH�� �),G�N��m�v��>Q��5=T���;	���_��\�@(jF�EJ����@��!:H�Z��=v�;�uAZ,H���&�_�3�uw�����۝ֵjd��L]P��'&$O� ��T��)�tY��8M\���1:�nDou1.�QV��������g^3��eN)��k���A�q���R�6�(ޡ�iZ.�
 ~lXƽKY��ؤAI� MC�����Jk��[�����w��Lߑ	�������6<k��gs�fr���Aٷ�Ƀv��3bX�#\�hC��a=�.�f	@���`��D��دdM���_+KrEܼ���, ��tl�s�R��2m	�@Y�������X{&�jA���iU3i��C������I��>:l���y�g�,?,aA-Z�q�
���L�e�,ʲ�.�(��(��x�n�=é�;O�}d�f�2�H��r"�07��`&b��j�k#�*��w�#��7(6&�(����F�C�|�֏�6쨫�;l�B�Ǘ�/���?܋z�Ӊ��=ZL���ه�¡f�1�f�X)���eǫǡiZ�=��=������r�m	�w٬s���M���6���"cV��S�2�\&^mkdl<n��D���ޅE�2�2��L%Q�̰��H"h�����^�ƁR3�'+hi����1h�� ��;�X�㦔^x$=�>T�����̺9p]U���.��N]����)�3`"���9V2���C��4���㠳�B�f��G�#C4� ��sD�x��|�I�6B��^=��i�w��s�~&A����5�ZM����Xp�ȇ�4�Yf�M�8��MO�6V�ȍrV�<Ă{�?Q�g���b=��v{�*���h�l��Y]��I�ʅʆ�*.�po�<�H|z���@�V)��ѯY@�-h+e�sPkZIջ��vo��N��f����h��.��S4�����<�D��诌ޏ��K��T��t��b���$��95�ޒ9-��$L�_�ʮ����+������D-���&��t���?v9����a[�(�\�m�L��ik��6|�6�Rn[A���f��J����g�Yi��T�vG�'�O�M���,�[��%;ʢF���)^
�A 4�l���1l8l���}y�ڔZ��\��F`�\
�:=~zJ�*|G�l���%��ze��4�U5�y����y������	\fETYF<?�ۭ��
:a;#����ߪ�+}G�|��z����)��)���4Uxc�t���E{�O��,]�Y2�e��H@3z^�r)
����;p�� �c����"�r7Thzc����szyJ�C�,��r�Z�ؗߵ�F��M�p�����J��f�IF�sJ`¼��)�Qdl�Wt�zC���o���\J+_F�*�'���{�	�=�%�����l�D��	PN��t#��8�ޤB����dZ}^�W20�L�a��d���X���t]�7�ώ����'��k;y�Ѕ^B���B��U%�s�кnY��I���W��+�Vc�� �7@�K��d��8',�fQʋv�)�.�e?���V������~�{.?����ſB�0�+c�ÀC=M�ۍ��=���T0f�9� ����%��[R��XS�|:�`3oTA���E����������i"�]9�T�-	17k�>��=]Yl�G�_=��L�B�q�UC2<-H8O.�d�|KL�����U������=X���1����ry���䳃��d��(W!�_�.��+���L�0D�C�� ���<��l����ֺ���+䯳i����II�����I���A�ʄ���Q�gv8�Fs�d1�$�6TxN�/O�k3@�r���xH�W�V�#�*nu1��d�"�e��D_��VY�����Eǩ}h`BO��$�6x
~�X�� .��6��f'c�ĭ�U����F;���?A�=�Um�y~L��<.Q��|Z���:�v����o��o���]���}�����������D�Ж�Ae'Ҿ���X��[���Еs�}���" [���B\7q��v�W�����V�Q�/�9�S�vB8����{�E�'���eT������C(�׿E1s�,P[R5��Nf���/���<��4z��<�Z�7I^	x�B�G�q#�abnw���]z�x�q����X�!=Wڇ�Q캭cG�80 .Ŕ/of���7�/EW�(�,��N�I[ ]�t>�a��!�-�7���u���'�qO3�G��K�mֽp�ޫ�=�dͿ��~��f[����[k�1�c+[��b�t�Ӝ)k��Y�Ȫ(hf�UИʢ��G��&7B� �KR��o+�yyWˣ���G�TU3�lU��~���b>�E��ҷo`�l��e�_è�P�Wi�D:����k������(/��z�6*	�v��Q����.��#���\�|���=Yɡ��]Q��E�h��R��݅ɗ^�%v�[h��7�d�ϸ�H��b��\��U�\`��pmDS1�f|�z3v��*��$¬�j�lw1��i�4��zl�����cצvj�ڢƩ��ۺX�&�T�6i���U87'���4�l���E���%V����fM�ϧ��.}�.|vĹ
?^:_�L����R;
���a�c�Á#U���S��|X\��#�殈rȃ>8���ab(P��ʴ�bl���SQ�GQB�}#cv�0s��w�z�b8p�xW�Zg���3�64J�A�Mە&�	�aя��q�P�l��r�*0�DC.�0�}D�i�0)��jZ{�c�Ƹqݰpy*p%Q��?fF�ej�h:�Q������Q��׶l���vX���'N��ȉ;�g'/7���x: �U�B��}��
�q��V3�U64�Zim���nNtm^�zu�)c�͕)���`_֮�6Sy�9�`zЋ�Q!���RQ��s.��j�w��:�Y~���t��;*l�����l��GB��,�U'�^�s�lb�l�c'����p��殯ƶ�LDZ����#�.X��zC��+��t����d�W!�(�]�N�f�KH��UVv&�`A�.���!�iQ>��l��Fju�H��l$���N<a[]�v2�����T�I�G߃\�Y��F��A��ƫ8\�'ؘc�!�?ת�N.�Rs5 �&붨-��V\T�O4��HyxX�b�URA@":w�.��N2�WC���Q���� ̸�p�of����p!�q�2�ƀC�^ԊK���S����=�I�;Yt��vzbv�	g"��t�~�<�����N��z�/D��KHq�(r ����'u4*o'�j?�[B8�<�>X��By6�]�F��9;B,1�c�rzb�C�C�o���姊���!��r��n1�4���5�yb���t>R�.[m��$4H�������͛wl�켛ƴvj���H�^��a��ɇ��t�Yrb�7a�i�eZ�r8(����s�WxGj#s7��A�qذ`��7v�ڹ�$�vd���N^|k���/��٪��� �C/�Q�Z�
A~*�q�Կ��u�K��ɏk���l��[���,���a'�R��2l��ݓx+,@�5�l�S���� �$'x���k�&|?h"�����y�J=�C�ʰ�IK$�jPş_Ѡ�PΓr�Y�d4�7�-�4����l��J�������""KgJ�)�x����b��b�8l���*�$�(���'4�e�RR�+M�Z;l��3.  �/�@Q9�k��1���*� �+��z��"ؠ�/Z�BgQ�:��65���i�Y�&���U�C�/ΰ"��
B�.�W��8�2Zl���WC��K<�Li�օ�u~[]@�jw����ܦb|O�i8O�
�N9�7�g7e��S�W �Z/u�k��c��$��83-��������+���ą�/p_��r��U��Yb�9�Y�b(���P֕3q��q�#�T���~T�X5k�{q_a�D�1��?���0y�HЫlq��u��9���7\�̄��a�>>�^�]}��]�#�s-@rQ*'?��-p�]:�����4K-}T��oRU:o�(9ruKzK��h��'�TzKy�������%���C�.`��ms�%�� ~�.�UU_�O^9���F�sr5�X�d��$T�`)�.%%H���O'|��#p�q���F���w���uE#�IvW.��K������4�����sI��C��i�PO�-�x�5��(��c̛�0��@.qH/*�H�ց��t�
��F������`�"�VX+�<9�'�t�]�. ���vd% �JfE-��Z�5K�fŚ��Kןb#�J�%�}�\���Tw앶�d���OW�y����U�4�]z���y9 ��.U$8_l�A���Đ-'k ��Oe {�(��q)y�wV�O ʙmyf�g�;�%���+�,Exe�9�V�V?d�X��゠>�+���W��!Kt�CDmυ���g��'r�AΫI ���,�U�7+���&�[��t�nŴ�����������KO�q�x���XZpR̸x�$�	-���)#����^8LV^��ޘW>NXNK:��P�P�I�a�,�p��ġ��ݒ;��.�����(oy��1orV;�� 3.tQ4�w�cB�7
����)�X@F�M���A�ں�B̻�����d�l���i��(!j~ب�.M~\�^��x��%'�+x5�t��4���Ж���j,���{TG_
]��f��QF��#�HE�aD2� ����B\�(�Ih��fg��ep�	�m(�%T�2��?,8sXt ����sq�a��&�S7[����d��S\��єx$:C�i��K�̜*���zĖ�� Yc?�eG#q����� �����5��HiBq��hW�iL�
K�iW?�8E��]98�l>�:�F��\S��	ĺ���~
�f-���	g�눧o�u����r�$�g��Ӻ�Ue��
�#H*��>=e�h�|�x���!��7+ [_������"�b���}�9`(�7c�Z(-ǄT���R���c�{���V��8���'���MkX;.��B�R�[<��92ũG�u�rW��Gá@v�9�ۗ`�Otd��~}&��T�&��T�྘��oy��`�]c��j�an�8��55"�V�-e[f�u]�ց�(�A<Tq�MцQ��i3�C�jA����Z#�1����EX"?JF�OhB	a�#~���2'�8���1(��S3T�8���,����<�S�_�i7�%�k\�Ѝ�l�99b���T�T/���>P��������v%�;!p�@���_	���f�->�u�W�d��:*f��m�_����C��}�Z�-	�bP���$ˎ�����Mv��է��7 5�������UC�>�9|�$+J�Ѿ�v3���p��d�#�r`T�+��3&�?]���~�"�0*7�/§6��+���%ܹ��	JB�s�)��6�=iT+2Z~?j/:̂f��?�l �@��JbU��N�&F��$��?�D돔*g	g�d��:~��׭a^(�}�J�/.�b��	��)6��vwV �w��ޚd�-S�+���2`t�@�ɤBq���y� z��Z�����Yx��J�\����{}P�Bc�J(��4��O��)�K'>���7o�ۅ2R����C`�}K��U��c�=�N��~��{���,,���_��0^���㚃ܞ)��e�zj�M�]}����6�8�6�n]f9d��0M��eX��r+O������j�oM��N!�t˪��:�`I�\x�[{DQh�?8���#8�pr4�؊(��>)%��F�=f�.�^z�I�:�p�����`Ix�����G��W��LF-���=����Jr��r!C��Y���È�iX�-o�� ��;Y[hz1(��Y�Ą��<"=�¨�ks���"L�Ps��9Ŋ�f����4�e�{� _~�s�?�k�^�0�/�z��,��Ѯ �^ep9�,�{�(��c����T��N$���2���Y�tN�m	�}9�M]�����*�Pay�O�>���9�2�~�=!�5���!��`��s�p�����<��$�*����TY��V-���)͖�6���o����\}���cx�[�������#5�eP1�-��pk����aJ���tL��в�A�H�)�������6�Zo��c/�����c�6��f��SN�Cx�g1���4��p!��1��V��u��'�p��E�I���x'��yYc}cYf1r�����DR�&5�W���ˣ��~,���|����oK�x���Z�5-n��7��Y�%�Ok�s���܃|%(�����>x�-�~4��%#$�)u����I��H�O�'��T�k���b�ޓ˅�*l�]/�~dgtbL\ƕT kh��vA��t
�����a��GÅ!�t	֏6���`J����&�s���Z��}q[�4/�oI:�g�y��l��N��b��{:*34s*0�P`�ԫ* Q���S��u.),�����!ci7��6yT��Z���>�!�
`�o9�U����#����{	t���4{���2�������g"jԟ��0�Њ���)��q?�L�S�1xE�W!��\��ȯ��ɆD��.�71CW�Ǩn�hTП��]�bnl2�/:���e]I.G�c�:�������[�@�p^�{0��
K$��.q)�͖e˝x�t���ϟ�d�08��UW6/5ۦR9�D�
x�PO�w�b�SΡ�j3^�S�Ppr�qCO�i�z��,�q�6�}��S�;�[��8d��X�BS�.�8��2,������v�B)T4��u��V�����%!D���L/eC6I__yo@�Ӭn ˲HB��<֋�R~�jy�	q��O�x���@�|���	V���v�No��}�ˎ�(���Qh��N�T�J���1L�hm��	�oYY�ߣ:u;v���b�e	�H��Wr�U�u�՛�UK~ L�o�a<4Q��U8zɔ��� ��P�P4��ߤ���3��u3�>&ʾX�>7��'��	R�lAD4���v�D���p�r� �W�`�n/�����K	!��`1�u��˔r��΢ad��q�8#�L��wM��	�xڨ���;�>$��"������|+RWAx_�9�������]�'K�TC��~WO�������\�`u
J���hnӔ4l���ֽ�Zo��~G�	��-;�������+�Ǹ|��2�Y�\��J�k�F��UJ��m�$�O���F�0
c�lE��L~	�����!^w�o��k��K����:U��B�Ma��e��jPe���_��tm;+W p��� �7}�ub�SgTh��E�ȓ�
�>]T#Y�i����s��J�!�������n)1@���)��NF"��Y�W� ���^��4��ê�C7���Y��Ub��^(�yi�a�h��!K�FOw[�ȉ��v���y ;��9U���-�vK�t��Z�f�V�aI���+݌H}򹷈EܾI*��A����zpx�g��ǾE!� 0�n�cPL���^�;�2�X�+�R7
��ö����s�$�F_�
3�]%�Q?}�����jl��;6���\�}�QL�_��3��떆�A(*pl����q��R4�P-���K�0;���Q����w�r���r�G���]�j���8��jJ��q�D��:B]�h.`��q�j��eN6��t/1����=J]��Z���3����A[U]f��K>8����=L�F~��)��l�\U	#�*��l���R�F{��]r�YׯyD%�?��u�*#5��َ��*��m�n���Sr%s����BD�_� ["�6�l�OR�;nLʘjw���S�'%� ��۞|ݵ��7-����-�5虶���@`�A���U�.xk{�Z���|k�b�9ݳgu d�e� ;�j���O��v�8�W�����l��[��O2��g�g�y3?G������-w��U!���y�ۙ�<���F�y�N8{uQ����P��y�kc>-e���b
K�tW[��N�}���ޚ�1�QC��jdԘ�	����q���_�^�KQ�3}��9����"�/Զ�FYK��G�)�G���z	�ں����h��Q&r�[v�`��u@l��4 ֻ�pxG���r�,��V*y�vLѹq�l[��I�'�z������ˣ���H06<��x��6�E
�`���%�m.ָ.��7 ���D�
����]{烣�X�_$a�R.4Ό����N޾����
ˆ�P���7���|���~�K6���F�M�C��
�*�l�b����f@�i^��tj7z->�������_)�00m�z^��mNӿ�#�����Kͫ��l�f���J?y�j���}:
��Q��>j�-j/�C�O���@��n-*��C,Pw��|���`�Mr2Ԅ�iN6#�J�4�+��}lT?���:�95'ʀ�{E��6^S��Y�J��
��ہ �'��h9Z:��ȴ�$�Q�s:����ΉW��Q߻Z�Df�x��`]@s)ۮH{�c삕>o���E�QW�հE�geD�,T����B���R��tg%�"h��3ټ�h�$��:M���6�(�t�ƎD2qU���0=�b0N��p�.}�z����p-4Z�h����t�;��{���y�8��@}Z������R*�	�]cB�ǦM��<��Rʝ"�{<L����7��E��C��`�l--��Cn�=.�O��R�ǻV��/�:v>��>޳�Y�TȗIZ@�s��1U}�@:fP�9���3_�������|�$��Y����ك~��W��PR%wz����8UB�j�<�N���� ��B�%<�<R����+�C�Am�yD;��,c��9b3�i�f��|�(F2�\~u��+R%���-�Zrf�E��7�\��7�o�+;
��+�P�A��a�2z�)�/]>!�����*#����d�����RxR���jte�����p8��k�C%>`�j��ݐ��ڄ�����Y!�����<�������l<�raT;t�!���kNjƀ�%IY��<N+�Kp0%�|���;�Y�!��ӑ�6#��EeIN��Y�F���:���v��I�݂�_{�@�0O$N���3�����x*� ??�S$�Hͬ��V�!�a�>����)�l��pV������J��V�A�RA=K]����)U���՜|/x�@	=a[p������jҐ���ŷp,��R�ֱ��+��PՋ^�Eh����d<�JQc�m�Ϋ�?��j�)]t� Q:�;+���.�YC8�Y�"x��0����u_��~(�}쑼B�ǧ;�-O\�̂7N�Q������Yh"�\�`�׆�����ID��$�I!5_����C7W�Z�9�;�M!���d+2u؍���PpOæ�SP\v�wj6R�����F�g�|'�4�J(�Ʉ]v����4��"��/6by��t"�3kx�~N�X,��u�]�amN������C"U���I{�{���i��(N��ס$��S3q�e\߿4�L���HؒΩ��Enqg��r���Y���X^�1G)�H�9�IPઓ���~ ��G�C?��lO����Q�M�l��d,,�Ym�����Tm�ᾃ>�͠ �x{���dD!�q��\M�N������}�و��{�O��3��-X���,����"K��?�4�lDKd�U���g��'�@�b�\����.Ơ��F���ã�-����n�)B���h-H�ND��7�N���OUf�=����$��A���Y��� )g��,2_�yT�޷,pd�u&�NQ*� ��؃z(���J�k[�����#h}ךld��^�O;T�ƩR�N���YBc[��V�ޫK<
i|�<�?z�')���-�Kt��
U�G��N|_@A*��)��6���B*��Gŧր�Y?}��WOTd>�Z��N��ד`�ˬ4�v�e�����:
��/�2���z������#Ւ���̸	��T��J�<wP��������-�ܾ[���������9E�ڪ�,�4m����.7����cJ��I���޼�^ę3!;:ă؃�$D�r�'>�ʉnp�� �[�% R>��P�%��ST���w�� aqv66�G�ʊ�#I�\r��A������(�ND��C���������g^Q=�ʷ�nX�6��$&㊈Ɂ���=��JX�n�g��)dIWD���~�65+#F�������u����T�1\�j��<>0o=�B�uɂ��:7o�΃�\���`�=Dƍ=I�{T~����f>�(�����Q�W�h���Js' �9;����<�o��A�E$kRA�(�P�s��F\C�%ۺ)Dw�eڗ��`I9�T�E��d�:x蟽2�p�j�T@���GSj����{-{��Yj���%��j(Cw�	�vD�LH|�G=�l���Ƨ0"�&�G��<�ƚ�Z&,>]�#>|A���C�8ՙ�n%]�ܡ�4A����t�ߦy��� �]WXX{�L.�L����,DY���I��8�;���Y�x��3Kd)�y1�IX�7)'[Fb\�nV����k����q�>wh(�l�6�o_0˾��sK�����8y*�x<$���R$�﷕EC��7�����ُo�.ѫ3r��&�֥��|+�o{�@��{������"/�ҽH6���F��Gj�E�4�ƾ��:������(5���B��Qk��b���y{굝X��f�cI:�ה�`Ύޅ7遨��RǄ�K󣈼q��69��S�5,u��Rd��ϲ�B���f�E����i�w;�?iy���G�ڬ$��+=7��w	P���EL���q�����:6@,[����`��CL�[��4�%FA�����e��b�`��̊�4ꭊ�EH��p���:�zJ���;�Q9.�bN�=��-��
��]s�Q������)uH;�@U�,�jP�S/2*~T�z�8�r���p�Pass���~τ���YN�e��F���&cp>��8a<_�q�t�>��V�}��r���pF0��W�w_�@uQ~��O��}ńI@|���=+�lQ�~�3�7��;��D����h�s����_x6�%@�}��H�f.����k�P�	|c��.h�������Bj�R���2�s	�u�q�	&?[�0���@��Tu~}����F#D��F�Y�4��*{�)�B\'���.��O���> ^�����w���\ٚe f��J��٪�� �����6D\�1ȳ;]��*��2�ʿ[�@CT�����2>lP������n�`࿴`��[im\h���4����V�e4_$�ct�ÕuY��FAC�0���UѮ��� G������^ tW�E36��������'� 
�������gc-/ vX����D�3.�El9b9��^v��d�:	@]O4a&�j�)�u��x������Ԝ��@i�t�F��%�y
ow��XcK��<�J 4�wQ�#Jw�0�d֘P� 蝆� 	:E.�x�,���Kgf� zWNfӠ1Ax�G��1�\o��%��"B&ms�ܝ�3��	��jؘU�伆�%"0Y��1��V,�Qh�w１Y��	Y�^=P2��ܑ́���!���=Mɺ�bA��,ᮦ�j6���fl<������:�u�3��dnx���������u�<l�nqf����0/��wլ�saÇ���t���)r�s�ʖ��j;㱸�����+�c�쿈n�8ao��� c2��L�j�K�����f�ؿgo�r@���(i��m��m����n��n��~���t�.��a9J��Y�l�|�� *�f/r&]:�}���Q'XG��0���'�iQ¸��_�bY`
Ia<P%b ��p�4
�#���[Q���-�z�u�@o�0c���է�^�W��:��]:��Z���M����I�� Y�wJ��Rq�S�	=΅�|���@���w�e8�CK�z������L���jNzF�����|ӑl���q�+R�	�^\�{��vY/��ߨ& 'Nw������_�V�nAE���jx���=Qﺸ��(n�0����U,��t���lJ߅mj�[��i�$�+�����΃�ORw �|k��k��i��~��%d)T�9C���g���"�+��ch������	�/��<�!�uKX��o�\%�U"/8μ>7�/)���V?1^�|&��Ty�o��u��\� �����N;>}񌠨�Q$� �)Zl�>}� �н��dd���!���N��*���Q�g�Φ��^��ث�-k!�]�\�}�8D�ò!cNUnynX�gN����en-��X��*G�{̰�t9��I�4$]�l��IW�S��mm��34
᧥~4�����@�Es���KD�p������tnд*g���y1�m��)�K;���4�}����F��Ei�aO��A@�:��_���z��w��E+��&!(���Оf���#dC�A9�5*�Ti��{��D���� �?1]y�!�QJz����)m�ٻ~�J�}k���l��jZ��;9"�bA�sh�X(ڞ�ݼL����6�d�m�A�{��BI�4Ղc�����(&7�DFQ�L��x@�R<"x�ó��%B���A�3�ndu:�z��%�m0%�փ�bH�Xs�0`^�ڞПI�1����p�{%{���;�ĀȾ�"�k\X���qD��BG�Ҕe�yuVO�e�:�����߇��Ȃ��Q}��cbi�e�|)�@h��/ɖ
r�{�ҁiV[Y5�_'� �(�&�a�Sm�+u O�Yo!-N�)����</��ys�:��%����������}·3�S䱀�S�QҞ�P"�Sd��KY�!zn�z��Fd��r:J�å�;֭^�:CXd�Ȭ#�Dr���,(%����*�W� ��&ܪs�	�.�nt�X�`�+f�Ib���Dp�.P�T���9�]m3��Ṗ�T	׀�2V�5�o�ma�U/�ޯ��FW�L�����+��b����M'B���J��C���J�~�"K�(�i|�戚�tK����cy2r����RS4AAQ�K���������4��jxdH��_��SDXG�՜����JB����E&, 8�f#������9�̤��uhS���E�%u%}K�ӿ}�A�*��	��W��R���\3ٮ&Z�e�a+���z�ꕡvm}g^�|x�S�k�4����l��^"�0�潃U��0�݀fS��dV6J�.7:'���y��eX���b��}8V����X��w�n%c��T!>пC_	�$Q����|��"f��Ir2Y��D���VZd�z�?[bN�ֆ쒖��2��S�l�����������SX��:S�p�G(�,.�����$k��{W�0���vJi�vDjf=x��!�`�`�3�� R�r=�O0;�8L��N����[T�1R KG5�G����׷��b��l��%��T]򳜒8�|�ԙ��FR�0�����Q
O�s�~���� �H�.���< ,"���u'�!�.�.����ŃZQ��j��T�μ�dL�ԍ��a�Qӝ����G�4L^�|�v�i5���#�����{V��9�|9�	��uϩ�/�-���Q!.Y�$��^I������g
7�[�/��ȁ�����򪔕�5�%U��k��!d�)���VM��l�˸Ź]�3� mԜΩ_���ڎ��ߍ�j�ƦS���?���2��o��
m�'Y�<U��]q�SD�j�*����f�Ȣ*����"��i��&cB����ɧW���o�r�_��{�R�"|�^<@s�Xs�Х����R�߄ZE�\-�������o/�R.@������_VQu�6+.��h��I&�Y"�Xln[���Ŗl�ʓ�_�N�M��G�˰[��d7dX@�H�٣f�XI!��&?�*:si=���M�ڌ���n_��B�\�H���6�z�Bj5q �8��@��4&:�^�U�� `\�-}7��s�D�o_�Z�o��ز?�qub�@�?~�V̥<E�����}�/"�|�Q��&���5A�d9��l����������D<�b��ۈ
��6��/ ��s�I�EZP�O8ٰ�?�0h�X���VM&�!em���l����G"NE�@�j����3 |�INy�J)�^}��T�	k�5��ɣel���%] ��)P�+ГAl+����'Xq�9(�=�m9�`����N��1!͡�K�_R�[j�ʕ��T�T�~�0{י G�t-��������i�� 1j���������T�6=�q�_�)߈<֩��<`�u�g/�N���$��ikht>O�L�aQO��,v2��N�;��mF=��� �i%S�D1��Km�{�V"|�ʠ;�8���	���g~<���K�X|�q 4iA��::���?q�x��#8��I��b�Ʒ�.���e�+�$̨ȕ %1���	�{���| "k&1�e�DW����>�[�T-/�@w�P�'�it�s�8�m��C�$_.��n���h��Y^�i��^룡*������� x�_+���({ήzP��.)�-�!��D';�Оm��Y�l�����=sQ� �{�9[>�xx}�e��h�6ǆ��[t�0��*�-*�O�L�tF�;f&M�h���������a��ߠ�X����G,�b<(�7a���J�lN&-�p�u�^���7� {p�0~Wa�f��گ�h� Z�o��� ���v�+��0��]�-����޼�9�:<pዮ���V���6�8Q�+Y�2F5H�m��'�g)S;T&����]�.��bDҎ7|[)���%��ia���=D��h���<D��p�=A�9��#�-r�&Z��T (�P^���D߅�ӏ*��N�)�}��lH��rap"�I!�[l��6J�xu8��+2v��ïw+���O���b�5���+5m����y�3������,�����lU��;�āK뽺�-æ�M+�����ȷ�@�;�G�+����>��g.B��F��]�..Ρr� 9u���s?����w3���b|7������(��b��=
�`��P��wj:����T-Z�U�A��D�'���s�qUGuZ�?�n���T�a7���4���Ux��]��6?��p�y�#���tTQ��㱃�ئ�<�Z��&-?�M]#5����^[VFE����g _�>'&���Ԓ����?���<j�+L�@r��y:��Hk��6&�<=fY���v�j�D�u��x����G�>�8���?��J�q�
��x���6�}�8?GrY!.Cxت�!أ���m��y��F�&����JJ�w�+2�U^�;)�Jp?��2��ǧ��@7�sX]��G�Q�p�X������X7�$I9g˧���lC���5iR ��"ܝ��Qӣ� ���Oi*����`}65�.(�7:� &����P%�a��=J�AN܏�(��vT��HZ!>��޾5�WV2�űs�w�'�$�aS 9L�qz��& �8��y˩�Y���O@�S��D�e��A��c^~����Kb�)�P\��|�#����r�8wU ���������Z����/�O��n��<4n�cn�8_��,�|���9�_$I��W����>�B
�b�n)l���S��v���[�5
����l��A�.%�
�옺�b ��$߲���F������31^��>-lV�
�Ov�X�Q>
t쟜?��6��b9�[E�����ʋ	�>Q���sҦ�`�P��!(���pc�<�G�5�>'0��O�\	G��:��f����,7]w �G4OR�p�0���b\�5���;	~��:\l�U���/�.���>��� ��i�0R� ����8��AK����4��w����D��?�Z�.��p���MŋB5���;,�D��2t�#,8�U(���c��n.wa�Ԟ��+��╭׾D��`R|.��q�q�I*rT���f���m�d\?�	�9ŇG��|���L��dTp���L��	7a2�y����j00��7�H�� )֮�!�9�E���>8�m����;��#d?�Эث���%�cF��E�񣥵Y��\���y���	�8S�Ҥ~o�.Uk�kM/�$���	�u�ݾ�!��*ݱ��(b^�(f�@�OQH��ĳ�:��=���e�-A���Q\Z�Fd'�C!�����=c-1����New\��>=�|�~N}&3��h� -5��;�Mh ��$ �gbؠ�-u�0S~����껛@��>-E6X���LIH+��2�,6 �w.6�(�2Cg��T��5rk"f�۳���.C�{�9���Ը3�3��i8��㲜�
{��7;c ;N���3WL�J��/N�����_��jT�V%1��2��	������+ɷ��,T��F6(X�q⮑��k��8sK�P�=�Đu�o&gj��Z�n����IF��,K����20/T��N��|��b�Q�J�#S^~��"�k��%��4?�p�w�w�Pp�]�>�.�hn0,=�d�dT[n!�U�#b(�jNf�`C,�)S����8j@k⒨f�.��E�#�NR���4����9c� 1E3+�S�sף�̠�b�w>����ty�b��X«��f,��l#(a�ˤ)׵�/Y�T�L JG;�O��q�W���ݓddzw~V"�ͲGV�VZ0-��^K�4u��+���B�a��&Ӗ������H��E�"�U�#�I��S7F�����#n�������\|G$~W[��k�M,��U9\���U�����H�?��;F|��ج�Xxz����(p�Ah[>�<�����M�$�U!f��vTO����G+��̒�U1�������G�g-���P���wu\z�lh���b��ڻ�6���B��B�J�sy8]�h����1HN�;G�Ղ�~���ɏ#���~����Fj�K���4䋵ޭ�=!�󊖘��+Wg�r�E�
m=8؅�0�e@R,=�7��Cӕ^�B���C���Ԓ��e���4e�|��K��$/(�)��M����˼,u"��ݗ�.����W��pm���L�Vi�hZX�RWv�������e,�O{��YI����;������h�J�w}����(�����f�>��w.H�����u��/��x�,-gBC�,i��}��Px����W��B�#c�w�jQ�h���#���C �]ʱ0�rI]̣��q�Σ[�U%�dKj�]�(����oCz�밧�)��\so,��9�\��0׀4��7����So3�TCW*�F[S2Ϩ��xG��K�PL���^�b���-"��9Fqp=�ٝ��^ ��&4΃�ñ�VA�%n�
eӖ�����T�c�ޱ�K�|�����¢)���݃����8�
EV������J��T9�ë��zWƧ\�Sj���e	�>a-�\@�����N���K���O�4{�����X�H���z��
p�Z�ȍ#'+�]�i̠���٨�x�4�$BCt�+!�E���>tX C
�l1���*v�m	*b���_������G*F����&�oEe�T'b��������L&��Gc��@ꕔL��|&N%�Է%B�`K�W ���.F�OJ�#���3�W]��k�Kc'���=$��!O4��r�Zz7Da�f��Ĳ�L6�=�3�� ʂ�ـwI8�Þ�m9�����
4���J��K�^�����S��z
��U�1>��G��ak�a��,{�u/�݁%�n��T��:
���嶀��e�,4�&�Uo�%2��?_���:J���|�At��R:�:��C��e���1���+�W�ʹ�1�����v�B��ٱ	;�TB���v����:$�$Bi���N� 
l�u�U�������L��!|v�Mt.5 g-��E������A�Ry%�y%��q}q�j*$#����^��x��PM(g*�+!3�c�;�"aaĔq�����z1�9b�L��3���n���,B'��T��+�^�2�с�G������eYQ�qT����aVc-p#f��d+�Q��*�Ui��'���t'��a�d�ۘo���e��b9}���/6����h����v��3?4���R��E`���m��ж����6mO�Ó���ļ�8CO�s��3_ �]G��9��ΓYF�$��X�p�8t&�r���'���	2����us���֓�6l<�B9�wx���c�����=��b,��/���$r��8'��-g�b+���e��V,�D��+�
x{pU�1EY�8�K�_ꅢ�~���^�Kq��NbErTubb�&�1�=���B�6'�W�v$���H�y3�O��`�}�e����ƇL�v�.��s�(��zY�`�lI}~��U{aO��e�Pn l��N��*�{'~��q轃���.��m$��#�<��q��){�u����A-�)��#�P%�nm,�&|(]0�Ξ���6Eo}jq�w�8p�5�t&Ϯ2|����e�\剛�'r�zѷ�h��'/�1�(�4݆2�wU��˳,�Fg&�E���B�4��8���kg�|�������O� ����ܺ�֝Z[r�]�,�̾�/�謕_�ؤ9+����E�,k�L��>��?��b1]����Z>ut��������,]݅�����Ue���r	>�:���iI��lE�*	P@�Q��2�H��jy�5�E��U����{��p��҂bmїiD����F%�JL��iXv`x��Đ�x��#x�_������;�n=����GQG�osGBw�%�6FmyTDpA�S\0+�	m����bu�����ȥ%�DT�O:z�+�KU�$��h]9�F��6�M�.w�ϋ�}[�l�9˱f�Z�����LbS���H�8<k�%���u~�>L0&`#������A9�Է�2f�`��^�l��<�{O�Q9A����"��R�)-�c0`�6QY�ڍ��)b ��m8$P�G�j5rj�����`�n�V�+�y�,u�U�,~kqy��++[���d�Jw�|�M0V��׎й_�^�)�NA���XD<}���ţ�|U|;��O��X^��:�:�(�����z5�.95>�{��=n����f��mO���e�PU�+��֊����IZ�q5����T*̓s��ұ�Y��a�1�Rc"�e�#�Vϵ��D[ ��|L���@�1�q�%���z�]$��⋓��*�hL�pY��ܜ��5�U��`R�����D�TDh����t��):�1��ܺ&�6A*o��>ߨ�&ƚ���Q-�� ��/۲䢺syq/�$��r�E ��-g�I��:j��Y�� ѮtyÐf�v�Č���AM�n{��3[��1�פּ��s��į�xw˞_`��n1�h՞2��A�o(m��R���:crr<�V�k-��:c=������]U��Z�D�I�Л٩�Q4��t�b��E9R�S�NA��>� �v��d/�%$�U��1S%:���(��M�{�T� S-wt'�
/\�/!h�<�k@��|[Ra��.�O, �J�%�`�+�6KENJ�" ��I�۸�mx��	7]��@x�X����:��I�5G|['(ˀ4(�:� $]�,,L�2�O|ԇ�E;�N��:��ίX���d�Zu�������qp{�������{I��u"��	��*1JZ���o�>wiS�e%ӫK�V)qڨ�wY~Ó�Uaք'� �C�D)�Xl�S�}���@wn�օ��Jzl5�|v��`���ON�a�Ɓ��.�pY(�I[WN��.?�f��[��4ΐ%G��!��ߝUȺW�ꣿ�U���p���6���e万Jύ�;��K��lv6�hޝHw��:t��1p ���*_V��X����0��\�n�N�f��,���>e7�y�-�NKf�m�����ڀ��$���V�J^�ST�|�����PG�h�2�eb�RӚ'N�_A{�Y�@�2?���d���푣�oFҁ��Q4���w�����dl�9�{�1^�n������5~�"�:.b^�aCD`��׺
 ��4�����c�C���/�%ºe�\� ��D-Eq�R��d�#��1H~�
����/Ը��x��t�\����s>�S�*��^=Fm�)}7�� ���Ê�q⤟���T�� ]��U�8��;��aԩ$���p�E�*�����^���Gs)r@��^y#Э3�z�*�TJ�ڇ6��<Xc�|&恃F�կȃ�6�D��|/��
Q��juN,��)?��]mn��1w~J��0�F�R��5�������Mp�1M;�e�R*��J�oP�!��H�k�m̲6�C��9�yMhy]G=��k1y�a�*�&��_�?u�[ޤ��[.h��f���������������uI갷��[ɤ�%�-�?e������Ylș�q����f�=�3��	��w��]C����!����E�詤�d�C���30�?��dU�t�a�T�������Zt���D7���t�q|K�A},�6���ǽS֘P�c�㶜�d��~f���R�lLtѐ���<�0�O8����rhxS<e�M�Ơ?��"\�^I�88趸c^���V�4;��j�cз-I'r�����F'�\ID��N�����:w���M�})b�{��S��Bn��j6c,	��7o���)%�P���� r�ba\��"������!V(x���l�
۷�#䟺�Nm���x�ժ;�2s0P����=-�nL[�ϟ��m�-C����*��|+[��Mލ�������Z_���*@�Y��is.Bt+��w�:|{�/���S�	�R�`N��͖��VC�u<��i�Y��|�j�'ⲨK�[�z5���2���A�,�t�Zq!��l����"��4�M�7`'����a|J��~�q��t� ��4�V=aQ_��d�"^�j��u�c4�T;�y%7���s��b�-�hNE�����@�n���'��MRG2������A^3�1H�����u"�#��"�+��e)���m�8���q
j�5�.��p�� ��Z�E��w��,rp���}J���~������G;�K�����&X
�/f&�Ƥf�w�!�-��H�,�rĭ�xt���+p��$����Ǡ�:�j�d~�MRLeR�q��WސM�9�H�W�/
 �l�Y-%w ;ď��rJ����fEˇ�XI�_Q�1�:F2Af�t���SFx^T��d��gX��k���_~le!�3`d����h2N#@�s���r�|;k�I\�Ah�ҽ��jc�\(�-����h7x9T@8yc��e	m���Ϥ=��i���hD"`�TM�X��=y��c�7�X��΄9zn�����0X�����5TƠ�}�ܔ#_'�۫BIm�l�k�~@ʄ-S{���!�w�r��%|w2�\�z�]��<�w�4h2�j��e@��כ��"E[0��H~��ɧ��&��Z���������*��\Z���EC����IvL=f��4��#sQ�;�������	�H�ф����YR_3�z|�e�%0�j��kMˆ\�j!�z�˜�b�1�!e����u)�e֗!�_ܦ�*SQ��@�tq�r>��Zp]X��g�;�H�P"3=��uN��G�8E{��f.���_Ϧ;�?Z/��ɢp�^_ �|8�S[�uA���r㟁:�9M7�;�^[�>fr��Y���g(�1
J�l���|��ux��>^��԰N=P_n�d����3c]��,��A$Q��~��*�O�֯;�O;�6=�4ړ�[����hY aCoR2��Q;Ę��D�jk�?��%���|I��.�FL����V��;	_i n��PN\,�3c&����������M�6s�i�V��QɈߊas]*��0[E~B�T� ��E��G��7�o�P�N�Y9?d'������8��ԄZ;���S~����չIK`�\l���'�S0K79ه��B��!��z�Se�P�}PRPV`��N��W�2/��W��ˉ.�tN�*����86�/���<)�l`���]_;���ؙ&�^�/�O�-+���{�����cO��h�TJ�Z%	��h
�7���!�ߢ(c��
�;�>��(9��t����b,�a�Ë6l��UO�n!W�F�_sNc���]7�S`����P-w\$�9l�Li�Mi/�d�]��Ϸ1��y�����k���G��+ף�C�Ur���<Pf�0�W��6�h]l����ہ��b�ӛDt���j5t[����8@��u4[��:�)�-��g����>U�L�E���L����5q�.'N�\�����pyҞ�/W=�&���[�
��Jc�u�_���i�M�t������+D*�<{�<������]1_G�T8�M�����g.|-TW�Z҇�/ǧ蝿4{��h�ύ�VxT�Uݍ�NdHm��vƦd=N�z�aO�,���ϥ�\u�쯔p�Έ�E�"�m58����k̾�6|�O�秆�a�94�1�z��7��q�5�aƠ��!N^�X�<��Z^�a ?���eBO���\~RJ�	5��4��C��]%��Y7�kc�7�����'-�oU��,�m>�YY�L�'�K�
T^����R��D7�/�˙uR7�j/�
ݟ��p[k�١G�ͫ�C2��p@����e\�E�����5w�M�6����n߬�f���A3U����P�yv���ƛ$��o��������˓���0�5��Tɏ��2r@�u����:M�Cm��r.�fv��f�3ʇ�h�5�́F7W.o��R�v`�j���f����=Ù�k�^�M����R>o�	67���ː����!B��-[���>��+�6ʯ��@�<R'���Ԁz�pJ9�jMk%W&�V[]��>j����Xž�)zz���1�6��w�X�v��X�_��D.2�D�v��ۏ�:'�ew�Zs�q%׭}xԯ�Z�Y���F|���2DڎD�צ\�x�/�Y��O�b�'vD�m5x��}O/��Q�Hs�m��|��e���ttp��)��ujn�5�� 
�	��eXݫsr�!�'��2��g�PՊ��1��B@b�k������p��`���p��H@�t�g���=�"�KL�/��f��=
��Lh�#��1����'�ꂤI���k����G����ݵ�%} w�D��n��{�:�T;������0�?f��OL+�r���b��!|����o�{	_��|��]�E3%��[;Ϊ��$��I��!�~�X,񻠡Ȉ�+�I��4'���Pi��nD78�!ZI�b��=��fU�#�1��7/���ϝ�y�/}�oKt�uWN!�ќ���4����M�ٴ;d�ey���Q��e{U��ΈGd�M��-�!�+q�'�뎕E�R��58Q ��z�?҂R�����t��N�3ÂJ��@���%:1]�e.P����p��Uqp繰#V�)�����xL��)Y�u緔:�TK_�P�x�����;����g2�Ji5= O�=����M3�@1]��T!��Hl���<�}�8��h�&���H�MO��R�ˣ�;���/ѩ8ԅY�l�e��/$��As�#�/��n�D�NJ��B�����!#܄��qn�Fk�T�3�8ܾ�pz��g	˼��$t�Q ~o������8P?A��N�O�6���~=�P��C4S�a!�]t�I�{��)V1���t9�4��	��si&��ı��sv$��]�s&j���O�x'U���Q���ђ��Ӷ9�|��~Ж��o!��iB>�Zȹ�<0l��hkn���,��2l�ƶ��Q����D�zuk8�J�����YQ�6.�Dag�2*!���iJ}���N�C�*!т����x����c�qIڙ�`�N7tw���\��OI%o�W��ɊD��`�D@�j�De��F��gG��$�@�T���Nd�pcvKYy�Х�f����SSu;��*o�Wʟ/)㞦U��Msc����y���z����^������d��:QqC+�G�a����z,����ҹ��	���bc<*K]A�N��[e�3¾�YC��j��n��B��$�d�w�����X�zLq]�Y�FO�/�{�)ƤP]zh6�S-���ʲ� [���kfɴ?P��d%/L�h�ɨ�4��-f�	V�i��t��&˔tug�'_Z��Qy7�|YOVͰ��^�jJ��oz���l�Џ�$�>�F���6|��S��&��P�S��Ju���aYK�CB�* N˫U_�9�6�N��4W6ߏ��	J+�K��a{��A�}�>�ZE���.�w�Ѡ5��&֐�Y]L��e{*D)O�����CW�.��;�k�����r,����ϓ��b��L��׋�mWM���)����u������ә�wqL��/�=�xI�U絨͈R�c'Os��KG��bGk�s[����2DK}�w'?y�?4�:���r��B�������T1;�"��D�w	NɌ�O���V��;�{�|W�V`iw)�,S�>���i	��״��d$�V��	��F h�*�e��� �M��Ĭ�1�9�4�;� ������O,Q��5bH[��a��}[Z��۴�yA�L���v7�W�/�w�i��ށ׺_�5�5$�;44VO�d� �p=�y��:;�nU��z*��KX��A��n^#m����7M��Zs�gk���"��I�J�}�:���]�-��ɫ���w��3��
�@��Y�5���Q�9<�r� �K���<X�si���r�DM��BCޫV��|�=G�;�����i2֘���$e~���4�C�O�]��薨��{zf�Uc���;0�T�:R�eL��� 6�@Z�����1�R���I��#�O�}13-�tQ�Z� ��rf�ң�Z�a��������h/������r�k��E}ڙ_�Ŵ�ؼ�q��Taxm��ds=7�dn���L��-�l�\���B^��7�eJ@j;�c~$���ڄ6�e�Ӂ�|) �0�<�߀�r՟Lͅ��`+�"j���?�+��5r�"]̰���%�HVV�z�\́�����E���:�A���&@aQ���(���`?���\��[f.��Y4�{8��x"����"��Ľ�g#��s�����HQ���4<���"�ec��UWN�j����9@ڏ���q�_rQ�@{E:�AW첃!l�2�Kjz²�ơ_٪Q�7��$�,ji�3�x��K��L�X�c�a��!� ）�U��S b�4��b�w�7�2���]���8$�ܠ��ضG�OJ���2�R}-h3�u*a �(����$�Àt�0ߟ�1�W���bO���)n�$j�$��'����L�{�@%e}���o���z1�U��$e��_�0I5����Q���W�����l6$�/[O�-�Zs�������E� ���ʧ�C�E��a�M�5�x�X�O-�b_�S�I��!
6`;ajr,��9�S5�;m��I�eh���Vb4hH���jЬ��~�z��!:�l��r��і׫����j7�Ԭ2M1V
�B�U[��arY���F0ء'�:B�0���tT�T�ם[$�MdyY�%8w�71���'I����q�1[��S�YU+7w���vuS�/���ąѬ���5ܸFR�1����F���EA�F�,�F�i�7Aw�Uf�ϢNOI��:MP�{���_�c�������T&#X�Y�+�$윑Z���Ċ	_1!�"UA�C%�w(i�e<qy�T7t/a���y���W߁AnŬ�e(��Z���#��>���EA~����Z�W_5�$pH��^�@q�>Fo���YNM�ö��5p�c
uۦ鿉�(���G�vg�����=�������Z�xl��fA�X8��+(�o�.��ϙ8rVP_�� O�����t�7=5����<bO�4�2�*�  &����j_Z��1W�\Τ��Ji{�	/z�l/k�H>�e0>��řa�UO�R)��,�°�c뫾��R-�h�j��8G}�,���P]WgN8>gr�W��󲶺�:���Boy�C�`O��.= �����#�U�3�m���Is��|`��2����P�#,Xq�'�B�7��2ᗾqSUr��|af�����.�VM:��vC�T�_�j���h���CC�L��L�pZ����cN��h�b�� �
�zȑy�&�+f� ��%��C����~~��?�䏯�����SKD�͌��䂨j�ڐY7h�Ko�-�������F��V�I�sU��nk�l�}n�\���B�Т*����K�CeB��\�C��'ѯ+�9���������O��]�g�XwY�/�^�;�cӵ�-Ayl��AKY��@��m.�>��֮x�o�S(�S)��ER�����J5�ɢ51��|��Y/�P?^c��[Um�t��۽���/<S�=4��}:�sK�ɸA0^��N	����NY��})n�K���>��sʸ4+�1�ao��t9�}�X�)��{�%X��CLݗ�CR>�[�ݓ�Y�5�-[�g�F%-�Ɛ�dŗ��/�~�D&���
L���ѓ;G��-y�KG����մ+[9iCo�b5�'
�L��Fd'=W�A�7�c_�Z��'�[�m��\u� �6�� ����P�rYڦj���~y.��J��_J�cM�P�f�j�^�?�͍���2��"lK[b�B����1/��8;���o�#�k������*f�aZ��S����{)�������f�B1Ǻ ��V���F�a���`k�؍��J�,�	I�7Ρ�-A&c���:/
���]�����~[�,/ ^#N�����r$a_�G!#�]<a$�x����d��T#��F�菶<Qm�=���jq|�|���3�-Ӌ����˝�"p��� X��n�=|����)ˇ�l�\���e�S�&�r�X�q;�i���r�<L�7N.�-�c�������$g��ck��G�ǡ���6!5����k,x�y�=�R����D�pq�h��6�K��	5|�����U�v�V�p^��\���h����-v��s�ij%P�l�I쉶V}�0H^�B-�Ki�-��6+���ć��=n p�K���BH��{�P���Bϖ�i{H>P�-ŉ�����p-��I�J"1�RM���+�SK.I��I�U#.!���j�EU͛���_����P�,��e�>d���.�1��1lNܭ �yY-������8'{��֨ �3����6�W���k#W��ئ�R5UyX�N\�w�&wAr�} -_����d�=���v�Hn��9����/s���Eѣ���@�4�m.<�$Lz�ES��o��>R�9��8õ��)s����,�xJ�wB�(A���>��[.ր)��xp~��I����"U�YE��K�K(I#��� y!��#�HY���d�N���H1<o� ���G�:��(�h��C�-�*���S߀�q�lU��L�|宋e/�e�V��DS^����YL
?݊��Yr���V�-/jsR�����J�Ήއ���sI-Z#75Kp�-n$��	"���2&.�j= �A��I���o`�����S
"8�d'�]≺�c|90[���?%�ݯ��橏�������؉ 
G�]�F,}�rա��7Eɠ�n�AZ�"����AqpO�����9L���a݈���+C{��u���O\; ��U�n7��K��}�Ê��/mV}oI1���	�L��&�M�F&���P�B|��śCM%$W�.���,��i�F�n�#�]]��2��Y=�fL3�|�u�iZ��s/n� ��o��Օ�+�$4�Sc/X��&i`vHj$n�Ld����ً�dZ[��X�Dg]Pe]��"��[����+�^K�֧JO�}�3��.��u�oZ�j�J%/0��ı�x����(n�
�׋7��� v��ZuU��=2k�
�_^��A�J��N���x�e
�"s�,�1�J#hb�+~a�Ӈ�^sFB�/�0 ��������k�� 5�{-;��m�Ɔ��1����E�/����P3�����
ҫ16��f�@L>PB�c�#�U��F��t�p�����lC�~��)��,|.����tR�'m�:{�g�,���z�x�Ę�O��v�Ai�{����p{u��K���+>K�E����(����i�s�jM�җ@�n�Y�F6|p!�T�q�i���8�$�
����.gE��%4����o4Ώ�+��c(�r�# ��X���>>L��~Qb��Ȑ?a�t��ªܘ�s�A^�}!87��lx��55%T�22ۅ�[��]�]�*��$,q�<�鲑���c��/^����?d=S��F��Q�2��\�u�����,�+�;q��7����!VXa�.a���/��$�k?�*&���+ɺ�����;܅�ZwLک]z�������tRꤦ2�9��8��r@���$ON��h�^�۷<����p
,�nF��K��ަ�0�k���Nn��T@��"U���D��*�
cY	t%��[�Q��p�A�%��;kC?�(�)����J���{j�V,��lw{���*ߗ&c~�̛)����|�82L"m�Ff�\̚<�:4��L��x4_�]�H�#o����0e^�5���NQe��̐�$}r���OQ:1����L��5r~����g�J����l�>`�%%����2����o�)�@��iq0�{��!e�,.�a^�C����خ����<0_���F���'�V�E���;
�qw�Mq�J�ę4������3��H��<�XO?nAZ{�N�ԛ�e2������^��Ap���e��ݳ�l�
K>���p���Ԕi��� h�Q@���u�e�+���t]�W�d�)J<�}{�� 	�$��v�2?�pၽh�-�U�p�z�ЧS�uLo ]e�PzH�M����R޽���zv_�%�r漇��>^��	�|�>A֤l�[#"vd������~�R�<�}\Qlh�#_88�3�����jw}:���0��C��p0E狉��v�aZ<�����op���j�0��=EmfwP�
��*�%zO�u�XNgd@o@0����r��J�y*U�) Y ���QY���#8:�7��3�)-���+{zϞn�6)��.��H-V�sN����3H��?��X�� �,��w�߬".P�B�A�l#���NS+�e]�&���[�{��.�GGۡ_{�>wsd��u@|!�P.{u��d�n���z\�;r/��c �i��<T=ʥ����f��htjF5^G��4��ru����	 �x����R����̑^�x�G����@��$��~fF(*����P�c{�K��J��<J�g�� �Eg~��Wj~�)�2"������m�F�!!�tu����F��-ruɊy���9��T����~��"���\9ua��`�0N���#�i��ݕ�}ľ��bRgi�m�>ً�U���(HĪ8���Z^5�����1�E)�u��0��q����q�@?�֖9��(_�};��|�ry��6)����ʄ(I"�:�6�Y�6��JH�����W���!.q��T��6_2��}��f��L@��Ֆ��J��.��I_��3�8�1COF��J
��(#�:��B ����Ǔ�OQŧb�=Di(���9C�1+	V�t��J�B�W+B��
C�z���?'���Ӭ�Kh�6�?�X�\�`�M�V;ɺ[�D@�P��;�@3ayK~ޘ���]?oȌ�hk�]-M,�/RS�432@.a��=�PY2�Ex�����Q�l�w+aY��m:F�)s�+��%:����^|�j��,�)�OM��+AΎ]���{���m� �����0��]�t���R~p��[MG�hD����f��S7����7��h�,/b|��a&kө
M��m��j$)�(3�HE�>n��qS�8A�E,�Y�-5�X����M��Ѓ��}C1E�<˒�w(.U����!��v��c0��7��Uۚ�H������F�w��$"��t�R�L���/�>=V��$'����Vյ��8�����s~s�|��I��T���=���bp���J0���73m���G���̜�`FUR ���5�]��ߡAT
�?M<Q���K���.8�
�tsM@̮ǵ�q��d��®�Lq�TQ�� �����ȰK�	�ujP$�%�(��e�=e�9���}j��bxN  �����+i6�tz�<���%J9Ρ�q���5-�:�U�fĽ�������:[l��6��ې�}�T�!�t���>�ߐɦ؁��C�a'-+�n�y=b�{W�Sq�R3M��_o�uo"�%Z��L�i>^gI�kF�Fy�G���[��#�f�W#�r�
��J��*����x=�{#��l�l,7k��^���!�(�eӗT��c�O0�!�iAF����z�C>����]G���.�H�� ��R��?g^���9>b}L�e�g^l�癦[qV�?���֎Z{�E�c��������@�y��}!�U���ƅ������1�7W��N`�=���F�J�O|� �Ưkv���u��C舂U�PdS�՜����Cc��.MTĈC'�bP��Y��������l�E�;i��N�1d-�;�=E�2���`�E�f���&R��ra�s�;O!��2�ǌ�J����O���O��p�G?
�lf-�#a%�*�g�_�+����&�&i�+`��c=�=p�X�x��P S����7!�:i|ƨ
'}cߪb�j�Q�6o�j7��y�ʈ�d�Y�V|F��%���~.��o�u����=ݓH�]�$�q�,��w�Aq� �	�r�N�˻�n����_,@+�������C/E�!�X��5CY��9���L@���P[<K��GV�)��{��,���M�e��f7c4��V4#�gT��	lHC���)�D���͈m��
5*O]���z�qC8�E�nՔS1�v(�L(�OK�S}ƚ�d�XM�tl(������1�f�O+BBH��j^�D�C(���3\�H�j~pL�ANkD�F�HT�uش��s�d�]O�"A0?i��O`��1�F�v�v5j�CB�^�1u;&8���T����m�)l�'"9�2Ǔ�����j�n9��Ӥ
�(&�bw1	U�Nަ|���e�*�g�92D{���PRʝ���F�2z*�y{'�X�P��*��N���J9���wEW�Ѫ�hy�RփN�G�jl����u�"<�W�e4(g��R�1�/�U��b1��N(�o�{��vP��vZl(���g��:��E?�t�D�n��11�r�R�7}cV��.H��0����ȂS�1�t0�	����%ap��9��L삫UEd��3O���Nv�u��ܷK�����Ia�d8� }!��$��VXʠ�nm�JMHl��@f�i�ئ�����c���$�F�i[8��I+�л�¢��VG��	���0���ۢ_���D8ޥ.���x����㏹\�>��������ͭ�p�U:�:껰��6�;1`��\d�Po]g���>|k���QA%C�[K�E���Ѡw8�-��)�@��������b��$(��оh�t��  �" �e� �g��12&��{�&Q�`�K�Ⱥz�K��T����j�U�sC�]��j����.c���G.ۥ�:��7�P.�P�g��d�fu�1�#x��J��5��#��j�`��YY�Jݮf�nB`��{#nS�!�lM%�7��vc�<�5��^xf��Q�Z�;��%_\��n�������78##TwГS,�I��c��г�k�k��۬��Ve��N�v�Y)z��*��Tg,�lh9��)�i��q��!��"�Ŧs5����zU&f�_�?��Zkl0b7d��Wε���IM���ϖKQv��Mn�\ʀ���@�ǻ��$�Ʒ�P ����`��[��3���7�%���Z<�~u9=��9p�`"�E��V�B+�.]n��N"&� :M��^T[W,���L�i�J��$�u���\ BU^o �NJ&���~[��h�	{������6���`VYĝBǥ0�dAe�m��&�P��[	"#�ǆ���g�	PK)+ӡ���}!*���&���[��G?R�@���k��A8��Q��C�P-��h��oP�%�d�� �5ӭOPВ
���U��9R�P�Ʋg�Ù�u�fv��09�N�
߰�d4�;�ٹ@���[6�T(IG���6��}D8������Y�Gh�aA9���5���H�cvD��˽O:�.�ɔ��Y�.!6���R��Yx�8�S�V!r�N���u�e�GD G���!�=~�lI�n��������@8�Ld�t�+..T����e�"Q�t�u�˭(���N�d/�~>᪍���2^����R�p~y/&�^7���ma�I�ed����*_�~k~0�n1�`o��E?$m�;4�~ލI5K���
�kQ�^�`�hV[���*i		��6	W`�Z �������I��,7�2~12%��jY3��ɷ�v'��nu�u P㽜&D&�� ������xX��|�x�٨W5��@Ά�	wKg�0��J>�$J_��a<}�U+/H�wmD�]�6�O�)��M���� A��=���]$�_��E�u't��o�?����VY��V�8u.ᤞ���K�\/10����K&"��P��p,�W`a����E���i>���~�ʑ���nW�$��q���{��Җ�Z�x�n*�m9�����d�gŃ�,��A��̛J�A���qH.Sq����Q$[oB���G��Ih�8�#�o�5�;Ni������qWA������vV��Y���fG�8�}�J�X�e�cN~�zx#��t(���W|wbͅp׆o��ϐl�\��y]�sӹV\�ws�����ղ����o�׀��ǳiVS�^�fJC�h�����*'.��� F�޷��a��R�� ��ԧ��>�½����k��l%�s.2_UV���
��}���şb���hG� 	�O�K��0���UU^׋�����$ݼB&st��,ip�%Nk}�3���Wᙛ��y���sϥ���@�5HdǛ�d4D���9�@&L�������=���~�7
/սU�-��jY�w�����%�o3�1����g�wN���p%�V��sk���/��"���`����Bz&���V� �+�+!�]ʊ�+�BHl��Mç@7�Ew���B�y�r�6,`!p �Y���a)ռ�Y���Ӿ��"�.}5֠�'�N=���L����W+닁zzK1��H��5�m[lx\�H���ё]s�#n;�4"nE�NZɆ�jy�6N�n	/IE�Rrq50NW�ɰY
�s:no�H"]9��f ;�x����ޥ��d�J����`�;>6�,�$a��c��c�<�N�s�*�ѡߏ_��6�X��1����G���OE��V���pf��j$���6�]	����;�M<]�nAb�+��X�����$K&z7�8O����e�%Ok�{���vT��h��7�w=0^�^ʘ��d���,خ�,k7���8��r	($lJq%͟o�[h� c��W(�N�@ϒ�Yh)��ۇpU2��_O3!�t�[�B�Tm��� "X�S�V�cA���[�l�̩����p��e�j��@q�=��Ta��4]ZKb����T@�j(��H�O��0�6����+Yԟ����A>�.W�Tlp�H�O1�*�U��\_|��nd8.>��W[�ѸN�a���h/4������<��zW�M�:�0�f�^w&̾�(x�
�� -��s @{�����^���fOl��S�J����,4�U]�<̄���9Z���G{+�k�HHq� �����-j�K�1���c	.��u#cg��J@��(�`Y8F)R�e��]��N�kt�<��P0���.�T���̸t@��2h���h[fWl%� �\ħ|�<���#�BpC�B�3m{����o_��lE$<�!҆��iD\��H�bϗ��ݐW��]���#1������0O|;Z
S���!~M\o�0n ���D�J��m&������v"W�?ƻ��x�+/��g�Z=�U���X�U�թya��K�A`��v�k��݀�ND�UXU���{29��.���Lp��K���e@�Oj���T����ĚL�|�_��z�T�qc� v�_�V/庌���l3zYGc�^��F�K����e9��iT2kP0h.e�����)�*5X�㐦T^$���č#n�#l&Ж�Ck@¸E=��Ӑ��G�A9�gs"��H��Y�I���l���F��R�+�L��Kڿw��S�U�p�/
iD����8o-j�%��!� ����k�U0�_Lןq�u�0xl�ɔ��`Q2`�):s���l-%��;���_��.���p�� ��X��Go:�<|׷+�:Ğ�ag��}�'G�aɀR�m�C'��c�������H�],��������ٻ�A�[���|�`�T����@"o�dl��@�ت*�I���TX�sr7���Ze�3e?ަɁx�j�*B�Vi`%�h.�.����'�e�2��0���3���r\z��jL*#8}�eH��X�6��2Y b[��j΂0R��E�,z���-&�˖\٠
0� �0�jlD��kI�D�����)�oW�U��2��Ul���/ �[�r�}�ĝQD�b,��<"�n�h��n���~�=_@�	���᳇,ѷ�Uy)Tk�ۚ�U3��67iJ�Q^ȫ�;�q}��7�*��Wj��������Eۗ�&&�HC�%�ϊb�z�O?ƪ^����6�z�R���y0��!�X�(G�Cgl|�DIT���.1�Ԙ�4�L%�������>�k����;��A�9��)�c;����0x|E�l
}좢��&o;�O���D<`b���@�D�0��h��gl4��3���N��u��*����8�l�T3�%"�vZ�.�~�-<�[��uh�#�+R�\�$;��ʜ	�|���}���/|�6tJ1	��H�6��D��D=�������� ���Q���@4��oد�t���t�t��7�)� �H��1\��������a�7�Ӆ��E֤� ���X��):�a7�8RK��;�� �F�{���a�Z�) 
=^���cx��v"��{��h�sH��r /q]|�x�Vf#-�xk&�G3l~l��IJ�!{��)���=虯���è�#���ܲ�*�د�1�k��(������R��o���Kv���܋�f�)�v��s��8%�]��M
:�s�,�d�[��i3�dY6z�N�WwS�fj���$_m��~�<f�?i"ג^�]7����%vxj1@�_
*���;!�|��{�DYQ�֝ ��+r�ì�%�-ޛn��HK2��<�Yv����la�V��H�����u0H̪t��
*�H�9uðF��{��	��ٕųD�ͧ-���k�����N��d��#���IV���Y	��R��Rq�O&zex���������]�엷M'��uϸ!��2���mv�$6�v*!4�Pk�v�jmb�A|��!���
g2�.��'�տF�F0�DR�dC��MR����>�t�mI��]��s�h�����p˕�r�21r��Y�)ΰ4L7��=�,x�99����>����M�?<2yRU_��v�x��F��6�_A���Ў��A��}W-�m�1mNy��'����.6RA��*���B������ұ#��%��\.	�(w\���_9�\�'2���N.��&�n�n$�T&)3����7�%EM��x�j��U����5��!�P<,���ы�a>���j"˫^9g"�K��=tJ���-t3R��k�헂I��Q��&A)��� A*<h���&!�K���k�k��V��5
:�����C��EdN�WؚT �����'屽��!T�w�_�R�q��d
�  �n�gp�"'ѝ�Td�L��Y�����MA����t�"a��l}U�!"�(�]|�U��@�;���e�//����d�v��_ȣh�P̤�Hϒz��?��R��2�N���T�:R�3^���;��>Gx�
������>ۀKV{�P�.��Jqm�s�J��!i'�5?,
�듼��~A�Q�HUP�^f1�vqPd(�}RH�1�a}H�R$�x�������S<��Յ]�t��B�����HQ�!t����+eh��@)WCW����n�p�
��`>�"�EXTQ.]�e���$��JMS�uP���pT/�j�&����V2
y#�<mcg�D�r���J<k����;ɶ�\��Y��(����Q2� �Z���#��᎗9�Y���ۖd}B'���S��`��.y��m��f�i����A\�_F#֤+�&�'�]bDJ;ʋ�示��(�Į35��WX����i���b~zh�Ʒ���&Z:�h]�1��/X�x�X�\V��Ï���4d+�D�\�S�Y���
�3��>�+������9�Q5�P�0�����#�{�V�i/���TmZ�]�Q@R*~�}	M:����x�f��bņ�@�v�I���ñ�32�*������G�s���e}�7-���t,�G�K�� ���Az�_�F��8hd1�e�3�(��7�BىG�n�Lx���-�!BR
ɺ�й1�[�Pn�n�]r����K�܉ �v�7+�s�ˤ���l�-�swٍ9��`��̍#�w%��0��g�|ub�]ӭ�܇>��A_i�?�>�~,!���%�g����X����w9��5D�z����ҍ�����mc����"��@�e��<#d���뾹	�+	4"��-{,���c���g�.�#�Vb��W)k��PƳx�����B������<��L�^<F���'�ϓ�:U�"��vzP�As�4�h��E��V�y2�.3�K��H�M�/n����A���p�+آi�-�%�".XĞ<ڇv��鼬-��>���!�`d${�^1; ��OX��\·X�H��Ti��+j�Z��y~%�I5B$x�@7Q�� o�(I�Ź��s#�fc��ϔ�A���Jh�F���fHWLnJ�I��`E����{���)P������O�=�öK��U�>�Ѐ��r<���[�R��+3���t�PC�-V!J�#�lɊ���e�B�l����k����,� �e����F�צ��*d�[ә r�Ѓ�~�j�8)���h��œ���7�Ų�)ˑծe@�]�8Z�F�"M>ӊ��ݫ˩����ξ�h��#r�W�*�`�dU�����yS$�}�i���{#_��xc7"n+^�x��$ިo�5y��}� �,NT��9�&���f}�4%�jh��6{��c�[	uU��ז��.9�Cd�<�O�k3� .�o^�d]�-UI��1GƸ�<�HZ@��m�W�0ew��U�&��#zN��\��t�t9�q���������0�ϧN��{-�;D⁛�)�#�䩡m�k���.�bCW/��S�u�I/���M/�_ �}c��S.�B���W��H@ ��'�FN*8`-v��[���6W�����|,�G�IT���m��� ���ۈ�24�
�tk�r�b�h?7��P
I���/n�(2B/�k� �9+�q���	svc�\.��Sdf7�q����W����~T�?mF&B�lɕ����n�Q�����fv���V�.n	��h\�H]��hد=Jb���(��Q1T!/����T=�_l�h�}��i�W����K�Ǥ�g��my)m,���"S> ����̖��k*�@�m�=�!��z(&6GG��>�z�85�,�<��ٶ%��0Bz�D�K��1<s�yc�0�Cr�~(e��D_B?�t\����T깲���;�ȕ�@��w�˰�Cd �-;���1�-0�	J_���ߔ}z��\%������ ��:�QM�D�6/S���ݵ�B�^�1�I�����1t�oS(�V���WW=�����C§��֭ �]q �/�0}�w��
;�#��5��^���V�Kvf54>�/�v�9�O�ى���;���J�W�y �_�\���NQR
S�f"#��+-�PH4��^�8�zEX������=g&�_0�b��=1_x�>�e�K{�وj$?й�W���c��o�ލ����,%7���:E����i�r.�;c�r�Qw� n�qk��m��A6�
�
#)ܡJs��a�"��ZFק��⩻S&�
���#U�����Jq��B��<��".H�E|��Н_:$�ꚟ�r���bحl;/D}�w9 �{��Fͩ�)0�g(&�}�m�z����R�$-P?�d�2��1l�W��������Uېa�k<������h}X�LC��U\0�T����Hj����K�3�a(ͿK�k$�A[�v�AI�����N"��Q!�&�B~s!�ML6Y��\Zo�J}�r�зQ9$N����z����>!.�# ��&��K�o8�]�^!DD���o�wWB�.�Z�n
o�[T���K	�3�]R:/%x���,=g�;1�1F����������,vʺ��J�9L��Ϗ ��ooc���Y�.�Zs-��e����|W��ۈD�ڏ�>�g�D�\ՙJp\�Ą��Xq*�љ[rs���'s���(@p����适�Wb	�l[�'�f�s��.���C�Շ�:!�atn���Yt�*a���-p�[��Q�A��v��:��<��q�b�̀�wf �0���}�;����pG}�Vj-���s	��?���nL���٤�����Xl�B�r�7֡QxW2�p��.�b�P8�AN���uo���3�%W��r1 t� ��p |1�;L��S�_�-���'�fn=�0���[?�qm+P� �s}qK��KJ��)���(�P��iұ��D�=��\�9J��rz�(E;���X��[!����J��*0�\[��O�Lm�?�]6@���J�*O��>W��	R�4���w���y��чJZL�W-z�i���镴a�y�5R�c+��xL�����ɼj��T��u_U\�q���sL���#1�'��j��r�/'F^��w bL��*yo��1�SD��J/�k��b�@-K�)x� u���N�K~��4D�����M�O��Vk���?&z��λ��x�	V2fg�b�}��|$١��9��o��	c~Al�_��QV�6^=��(g��#v ��v`�P����x�ο}���g����_�ߟ�P(�%�������G7�V����7���O�S���齿�:�M���J~_�zWcqUm�	�]�
?:��J�Y�)w��5u�������;'�z�+���O�#F������;A�~���(�����?Z���l9��*�v���X���F5cpq���@l�c��!�$�,|}b4w8,oY�d~���-w4��+S�ǉ���wD4�Y��1/1e�9�����4�z��s�d�8��Ԟr�8�ZZ�-��?|}?�Z� =��n�ɐ����̵ٗp��X���`y��e=U�Lv�;�`��P3a����me;,�5��ڡ�u���/��!<g�[���5��g[x��Ȧ�m/� a�@����)\�x�s���mJ�u�Ą�^�bӣ�,�M9'��& ���f���Hu��}�ڿ��w�X�Bic�����a�&����(Eu���������c� ���2�x�v�J�F�Ş�h�3EW�{�r G����9Hu;YU�k ��rȍ��w +�Q�"R!o:��H�vv2��|�-L�K�SЏդPlQ��}T�Z����W�AӅ9���i�Fd�o'Y|<<�F����H!�nL�%7��X���P���a�9��5�C��|bT�j�<�*tҷl��g�v$�w.R�&C�R\���f�d�Jt���M4�NE���9I���S1zO��K���A/PTI0�ؔzF����@D>�T=���ȨU�j�߶Pa����V� @V�K� 7���v@�X=��b���A��x�5�we	E|R��&��3~�Oj�/e��V��jM�inޤ��@#�
C���5c`g����Y���I�\�6�=���W���j���[!MW�7,��i���Z_�{7#pD��p^:�;�GҸG��7pE������������Q���i���P���]=���ڼ�k�9���;�ZlO��c����4(A���k
�B��;�l;Pvk�Ye�5;���xm�I~��D�D�q��O���\����!��s�^(�6�f��΍��2��Px�'�9�֧������v��W	us�����Uv�c,ŕ>�H�/N8�l�;�E�哘�u���a]��i �sCn��/�C�OZNEM%^�9��������3��w����/I��YO�)�&�[��S'oc����F����{��9v���Jx`Ί\M��ES�K�V9�Sd�7��$M��1����E�4:��t����3�B�kO/���Q���>�����d�xɢ� ��&��>[y>�wҌ.a��ip�}q+��]�_�F�!�;,z��n��M�"��~��amCa+Q�������hS�uz��Ua��6��$e��E贩O-�q%Ȓ6�K�Xc�F���d��OC��хF�.HG���6�[���������؊�h��`���x6!����馿0���"�m�D��_LW_S�뚽�N}�B p�9�{��ƈ�L�����[�M�Ż�b� 5�~�����6k�RV$���ca�Y�ZL]N�;�{�"i���с�WY������[$�
-0�SH ����'��a���B0C���s��@�H7V��D�Lǯ�͋�/�8h��S�8�C/�����7�nX���g�w����i��1�Sd�1X���۽;���c1O]�V��O��(pur�!�|�0���{���[�H$�Q	Ma9�iͺDzFx}����r��l��V�@R^/g~�-p�FV�\��4e)UIL���S��C���(���	�� oC^�wx�g�0����K"bж���P���u�����.;u�m`J!R7�o!����*���d����e����7��@]���	a�'k��+����m�]�"����Qi$c����`��-)E�a�V�5߼D2~��$�?a$8�Ø!��b�e�E�!�D�PX��Iޓ����<Ӛ��1ľЃ�ɜ�:,.+�JpD�[0�R�?�NJ�Y�b�����b�S�X;lI�����+����Y�[���lW3˱SO��A��m��2�A9d�����q��`5�	i�[n�e��1IjP��A"�J��]p(N�-�����sPo�m"Ѱ��{"�AQ�$f�I @\��<��&ߐ1Sż��sC��<��,,��ݯ9�v�bh)�VE3���Ok�4)N��È9�
4��Q�2��QZ���8a0x�ml2X4ч-͒ }*�c��!�a��,n���pT��������rG��C�E$Fm������]��2�m�tW���\���v-�`� �7�(l���-�P)��:[�I|ߒ���bZK*A�9�m��t]X�y"�A� C��9�v:�ġ����8���~O��k5�v~�w��w�����8���y���qD��~������M���(��稊3���i:���7�o����W=hC����٩��J��W������@��I�b�$��S�f
`�Q&ΉZ!r@�zVb����Z���Xƌ�*B,�而b,��l~�O5�����Ҭ��A� Q[9���4k	v��я����ɡ޶�b?�c�Cʶ��e�_5	�^�V�hg�hk�=��,��H�W��7�PO^���?�
6�V�u2����q����3�Qr�_ec�Tń�
���q.9�ͽcG��i\�Y��5�O(p��`9�w��Y�\ד��T,��G{Б�c������;T�	�s�b=r�jS��Y�\v�����<ǳ�%���o����r(�H拁e���u84��//�tC�}�l}��*�44ps�5�#�^w��[��������Ųh8�Lb�=h�-"�_5玴u�)��F	�h ��_�� ,��i��|ƞ8����VP���(}1b�q�W�0|����`pЄ�� ��DײB`�[qePS1SցWկc��w\wq����8���J�(棛��(fF�9w:0�¹c�1�7�=�>x�v�dM��l���OZ:��Ŧ��#�b�wI�K&��C�����_
��zO�(�4孂�߸y1����"e8�z���HIoux�c�k��`PMXC�L:s���x	*pϟ-ѓ�?��ߕ�`C�;T�\J{,�������},2v��R��.�Å|zU���7�=؂�?�{��(��������g��ķ)
���t���h���OW�rR�hQ����l�N��DS]��Q���l�/}��K����/\�v�mUR��LY`xO6v�ᯏ"���lp�CA�}b2pѦtu���Ñq�����_���G�E�L����Z�r����d%�h+b�m�wyH�����j:)��4��1�8KqRuiGm��iU8���&v�M;��^`��,+vMP�I7b�]&^��\�Xd�,�z�|r;����m7]W��>��F*���[�h�{n������<Q8I�m!J��X�6�i�
X�q�>c�u��y���:E�Qذ��*�8��o��:�˿�pw;k@��k���.xM�Nbf�aҌZ<��;h�炶;�O���B�\��r`bÍ�-�M�
�|�������&�W��;s���ǆ�ǝ\��ͭ�0�
T}Q�����2wy'����ݘ��͚��̀-H>}kѹ%F�B��3��;!x��5r���9�@�W0@:q:��hF���q�%VT�h�����6�/#B9xU�q<Ǐ,�/�d�7��P^ͫWŭ)�Z���o�
J�M��.��,�
\ �_�s�c��_m�$����麿�����B�����l�(:4�֩}.H��b���X� ���Zd�[��n���%0��� $]���p�S"T	�I� 7�]p�-!ss����O�A��a3��B��ȕ�tdY�ә��(�Cu�/v�:�J[�/�! I�ծ\|�
M�{��~��B=� Q ��酠���/U�4��Ol�GO�yCX!��&[U�5TJ��}�%���n���O3���|��'z��tQ����<tE�R�
�	�7��P\�-�MW��\V���!^�ў�Q�<�j�������ƘN�^i�?Q�4���K�]�1����{	����!��NG��ç)ʞ���1�����*uļ�)��m�ױ'�gQǒ�;�r����b�ml�C�4��TT��}l�e���tdY3h#�Kud9ؒ}�����uZ�5����|�ER�~�|�
)����#LY2w�E0����{7�O&õi>:Խ�NPT7tXߠq������@'Gʎ�"N�+���5	��?S���GCZ1Gj9o�ͪ�)A� ��)��s /�5��K�����
y,���7ت'g� %�)�=h�v.9tB��q��ﲦ�Q=ީ���'~(ѮF�?��l'w�%��`ΏI��J�B-e��U+���7�K@��Y�۶�Nw*R�,�N��I��t��i���x��5��!�����g�����"o��E�+
��t1��b��'e	�t�U���t��H\�k�T�q֫%AF���3K�K��Û,�����)�!����MR}gBT�ݖH���G���Po�)��	�{PG��S���[Rͺ�ڶ$�M�d��IO�D������:5���R�B�������,�]Ʉ�������8�q.�b��7����k��Yyr�,���d�Gi]L�O�4�[8�~����$�������t:7���A��U����o�` +T�MK-��L^u�f�Vh�f�3���Y��e��r׌j��'#�n��ʜ�����oԾ��5����.Y�Z-ǲ���>�FH�1�B��"|oI��$���G¤�ͺ�u#NEU>�K5Q��dhM�=F�l�U%v�=��Og�cN�lY�\E"KʥYv�D��ţ�XJ<����k��I�����3A�ŪHܜ���3�&���
��i�)��A^!}�o� -�k�`C�qy�	�37�iS�ω�8�	�����2T�.ZN8��vG����X+D��X;%�1(��p�	|	��y�����.�mvX���.�=�qs6u%x�H��S��R�@qFQ���'�X2��nB��Y�z�+z��q��k�`(z�BB��dH��ϾA(=��+4���҇�����R*Q�$�� �b��Q��;(�]|��O�!G�D�=fF&[��¦2b�D>�����"�J`�(�0K5��vW�ȥ`W�1���T�>����Dn���a�a��w�6	�l �,PL�;�ʟiKԼ�J:�u�����-�܍A��H*g����k��l2��F�mc�D�$�?�}TR;i�	θo^��1R���G�|#�C>fa���,0'�����������@d���G�`�#C��k�����i��s����ʤ��E�;�j�ei;B%M�nL�t��>ĸqM�+��lP >����Gd�x�> ��8�K���"�:L�MU�o�Pڥ�=wb��:�&xo���_C7�?fN:p~%������>�g�Q�x�J�����&�O��
����}��6��岥sH��&��z� ��j�&��.�|��*ւl�q��{!߈,�Ь�#�^N۬$e��u|��Uq�-��#3�.n�g=��}g��x�2]�Y�9r�Q�S���bj~�;�]eиR(z:!#�@)!Dł|��Z�!S���ʫu_�U�C) 걍5��мϩr1�"l1��⧂
}��yi�7�/���"��z�N��p7gIN��у�N\�	Ӫ0bD�C�]����F��2p�����z�y_��q4[�e[��a?����!���w�nP����Y)Bu����b�щ�nÊw-[{��p3<oj�=̓ �53H�}o˓VwZa�h�,Yv؊!�䐳�1���qP̧C�4�|ε�0Y�h�%ѷ���~'�w�z ��
�uݞ�9(EϩNI順s�O+K�`�:2�N�K�M�@J��A�,˔6kCw��أ�(>�yB����ߛ���z���v����n�9zu�q�b��ql�ͻ"�k���m�ЌoO��z�#��Q�"<� 6l�/tQMd���7_�EX	�y�sx�WF%�2s���3��u.7|ڠ��'�����4����nd����0�<��t�6���|/4����	��q�.�l�w����xҒ,ўڋ��`S�nS�/`����~yL���L���Y369Ro���0Zt״����7�fP�<K�.֪OJ8��t,�̋�G3fK�|&n3�wZ-T�հ:����h�=db��:TI�o;��eoZ�en0˳�KΑ�r�X��nѳ�?�;/qy���S�a1�I�:Uf����~^Yd �LSL��	/�����.A� �(9j��@��j�	H��r6����G��P���L���.=0_�y
�_�#��jC���v�C��Z���U	�*V{c���o/)�iyD	�1p��e@�]��a�� ٤�����45��`G��K�'҃�!6�S�Ȯ�q"�&�Цv��J�r�o���D�96H�{�yd�g=�(�K�$U_-v
���q;GL]G��Q�)2��>ӫ%��2�4%�^9��3�5%­�+���xpf�$$i��k4J����Y�2v(�%˭���&H�eV�(�7�t9O�(�L�Zi��r.�>���&�c�a�X��+�_Qs�.c���}<L$�%/e���pQW��y�T��;�N�	S����Q���q�U�S��Z-�qW�g#�L���� �3]����Ϊ��Mb�5铎���^Me�r�h�24%�5e������~�Z>���1O����,b�X��y��7o�'��Yݨ�#��u򱇶�0,}\.��Ks�6��+qo�E�;��U�'��̮�|��07��5Wy<!��1}�I����7�4�Z���Xr���ח�ˤl��s֢c���d�]vɎ�{�q �.(�������厺�4̯�*C��6��>8G�d���I�(�nk�/Eo	IlW����l��f�W U	@�	#P�P�c�^�WbR$'^�&��F��Q&�tx��1�dޤy�6S ;���FB���ɇ���t�m��ܱ����v==z������oe��8}Ġ3ы-{K�<�e�9��^�MK��w��y�xٞ�YA��q`W&��˛1�����Zݘ��������,���&�T4�k�Ž_g���KYz��TK�E_%�0}�v�-�t�W}����kHq$xv\�ϭ��a��M,�C�ġ�
@ne"�Z������e�B,�0�AT�J'!S�l��5'9�q\�i<���ot4��y�����Mg��d�v���F�A��$BBӇlo��&K�7�`�r�ڮt�������0���P��9����-��xӁ����5ecr���� K���4a��a1�����@%FVd�@N�:w�����u.�1ko�sx�\RZ����N����L:֘S��,_���o0���8S�7�O>��踹����qH[�=]��H;�g,�N�n&�Lo
�/��]�6_H8���Z����lyP��l���-�-������w��(�����*
bR��'?ǩ�^�� �m�B���\S}S��G�ig�¥؆�^�R.�D�f��CL�.!�*��y�/H�13Ǹ$�҆u-��ᘉ:ILqT��Q�Be9�cDg&N�aBSMƀs�$�k�.��;iӅ��V=� x�Ӝ�3FkorͿ�N�ʉRr�n=�T���=��~>u���Ql7'*���) �H4V��[���
�E��\ޤ����y�b�����>jN2���*H�"x��a9ûs�3�zf����lж��ZC?�½|_�ؐKr�=?��/yfL�o}����Ck2�?�ʸ3(<ϗc�{|R�i��a��}��:�����ZZ�MSA��{��D3ă�{Zb@Aj���	�%�I��=�l$� �+<X-w/�{�l���Ι���*8�Bg�^w��6�Z�	��Ҥ�s�2�S�E�!o����Y&",��zW�y0�c���a�1�e�*S��H���F6��(�w��*xS��dw���`����.�W�ྡ����̋:lC��` 2���6��9�F�I����v�u á&)D�ǀEϗ��-���h#0�>�oI-����������w?`ݝb����DT� '��ü.<���}@+|��z*^�~!W�-v�@\>?X�s��_``�q�M�ܠ{����w��1FO�2/�ʙ�'�Y�W��T�5Z�5�ye���{2 �[U�������V$Zï��ѥ.D�L�+q��8
-k��椤���@c��R�13X���/-��޳�(
������
�.�n��R�Z���3���*1S#�L���Q���<�$�v��o�Ґ��T{��턍~-���|�pIҏsk��:iUl�W�ÍS��S�F�;u��a��{��P�n|����1����\�Ko~	�0��9u�ј�"�Tݤ;����H�æ��/=I.��a�	�oܜ��x������L\hVI;H)������>%V���T���/���Q$�@	-
���P=H[K{gJGF�.�V�'���9$���.c��*�ێ���v!�h��$_�^X� ��p
R��q{@�e^���~由��U�ӇߓOmT���͚ڼ0G��qj0��i��Yi�;�j�gW���R��jOM�9�84��x�" �Ƣ��~���ߐ��Q��0�E�_޲��JJc\.�N�|����I����t���d������� ^�:��%�!I޶���M�:��6ݪ��3: ��[@LV�X*V��_��G��뀶5/Ƌ�>��N*}�
��=44~c��l�gS�"���9�eِ��h0hgt����-A�󺠡�ʡ<����	֘�ϛe���K���i9���L��a���AhxRwa��)����C&�Ag(4Czt��ָ�ς�Y�2<i6+��-k��-�eKΖ�����!i}�OO��.^��+T���#�O�Ep�V-��E��$�x�L0.�>f�(I��E�l��5BH����p���tʠ7R�*�>�[���`�/�#5��npo�I�#ͪ��\VV��������ٿ�=cu�h�FXb��y?���Lr���y�ѭ�P��Ł���vc���[,�VS�مr�"G���=ָ�_M[�����e1G�޹�T�1��h�_�� ��w.����=8W��k�	�d�D��w6�
�������ئl������y Kd���ǔb�r�Zٔ���WT�]3$�7��`��e��m	���k�fj�v�ˈ�ػɚ�$l��l6#��+K�F��n�z�Ec���~t��@i)�G�Li�4�\mA�C�1:�Nl��'$�� ODĩBW��D���\A�`����m�$�PB�{���OM]�2m4�w-R���۲p�,v��z�ͭ~�H��9��W���O�}�.�����;���ԉ�|\@[\�;�wL��	}������ly�>}� �4w��g��^*f�H���������S��wY�����Fh~K���y>\� ��h����j�O	�;��Naҗ�zFMRhv�лÞ@����'�w���V$�ν�T�s�V��?I�M!���л�k��<!�#�rt����0Ħ��-��r@o9���l��4��8{3,�������;��h�=߅Y �Hu&�����FO�
�	��	���J�0	���2L,x�3��<����9�h	���5��}N`��o�g�	V��("v�/�Ԇ5���E��O�4IH^B�#�h����RޟK|�~m��}΢獘�s�h䝏§���yDFb�� +�f4���cm���p�q���}���E�{�K���h'	��E$O�T����"4tt��C�P��;��+��I��!Z�񶆡�֛)�PȻ!y��.�X��W̞�R������03��Yף�FW���֢L��~�c��v,�LQ@��!i�.����S)@i�3��]q��tJ����l�w=�{���a�Wl�� J,t����(&Σ#��L�x��GH7���"0_Hmw*�|�&����7��[�	��9\�D��{��u��;E����M@~o���4y��Ɯ�t��R���� /�ؿ�T����m����}!�h��T��������I@ 4ߥ{��S��z@�H��~(l�e���`N@=���(@6�|L@2:s��wh�	�D^**/m���CX�S؆��1.dsa_!!���<iUX\]����u�4�Nڠ�01��Ձ�b=�E-35}�e}���/S�C����\&��!�s[��z�[�Q�g�@ �t�3&�9DØ=�?eO�!�r�9]� (�E�!1~Jy�No�ٸc`KeAh�̓J*U2��M���,+�i4��z悴%u������\}���ե�ق��Ӄ��E�:z��a��;#��h��;e�����;+G�t7�4���j>���U�A�߈|�ǗH�����"9�Q�q0笋�}+���v��i��`�E$j��QA�Y��IB���o��^�	dWSg���0Li�h�rw��M���!�2Cg+�7Ct'JQ�����C᝙�m'Ћ)]�kt~�0h��Z�x^�>�Go��d!V7�W�g��v����
瀨s '!��1����ErHVq*�!l���N"�_D��G�j2���	��!�la�'���ql)H��=
�f�=��@�	�����r]o}���Ǐ�[��l��B����ओN���ܾw��s�4$U_����l ��{W�����<O����UG����'��xj[mޯy�e�I���^{�L��P����y��i�paa��_��j��\���Z�z1��V�X]W�iF\/��|�_g�!|6 L�<���P]W�����p�ᦎC�������^��3�m	�-���ps`2�R�n����1'��F_��Khko�l��i�D���Yu\R��+{�D05\�[&g*��v�����pӊ;��1&M/1q��*�u��k��Ș�v�N)�?���5񄞿)B��4F��\��c����w��
�������7K�V����_���y�y�Bg�������c����U���G�#����w�������w��V$�*���.h�[�N�޿/����؏g�3_KmS��x�6�vūG4�9�SP��HnF���z��?=K�ؼ�W� ���ڗ�G")��xZ]?���3u�o��Ո�z��Ž�l�t`cT�/jE�Ԙ�5��$@�v,-����I�Ms��t��9瓼���`���{�g�o�����*��'>��d�5���3���Wv��J����i��=R7��)��eH`1`��q�+��������<$�	��t���EQca�n��c�Ej�;�����|�*�)m(�k��>���&2rK�.0���˟#��(7�.V-qz����Dg��[t�R�wP{I�`5������ŭDK��c���Cݪ�zk��A��h�\8�NY ��{lw$�ԘP����i5��%|�p�H@�FH��vo5{'|R!�[I��V(�]�e#{�GMe�>��� �����a���ja	
2�AJ�67��eW(H��t� .~NӁ���Zu�gĿ��C\���)�3�/P٠>A�=����9��ܥ��!)PB"��&�u�Zq��7�r2Κ���Y�6m�;B�"pe%�l�o�2k��>9|�1�r7���Śa�1��bb�O�Z���	��|�(*n�5;`�`���ܴ�@K���Ax̞ue�e�X��i7��,1�-$S%ƕ�ĭ9�T)�*�mwy���:��p�)�?B��l�Wo��l��N�G���1�0%oD!��r��(gj�P�/�����K�A�v
�˭��π�U�F��-�z�"��+Y>�d����E��	�?�����b�J���qџ�����o�jH��ͷ���p�IvŰb�ͻ�^L`�0a�%��z]�'jV$��t�n>Ѡ��=Ѵ����6?\��u��{�O�n�����ꙛŔt����0a߿Np�P��a����_�R�{��p�'���'~/�6��u�C���I��n�z�ʐ��dY�?�UI������[�m뉿�P��1��0Ic ��7��(Na���GN��9i�2:̰�z/H�ڬ\  ��hP"r2�
��\��F5�`K�+W[��J��Q���(��W4���o���7�w��U���i�q����=�����"e�
� ߏ?���Iu�z/��[p�,����8��F@�~+��%jz���������ڎÖ���h�����n<$���h'�N�L�oq�r��@�N�p��5�?&l#�ͫ$&?oj@G4<|f7����EB�N��i��g��k]��f�Y��ڢ'"��} �/�>���֦��#�^�|@�˭忞���L�$ʃZc�������HQ������]@ލ(���1�d����r�Yc�zA�u�~݇r�L�;Y��0�0.�u��к�SӎD�x�����u������� f�ah�e!aM�R;�:����#��؝b!�����C$"�jn���ꆅ_�7D�l���*f��f��M8�Pj�Q�wT�����5ͻR����-o:���)�FL�!�]�C�6l�x$yqC@�6�qW0�R8�'�GZ��z?B��֎�S��2�>
�� kbk�`��pi��$�"~|%�Mb�+�8?�kԮj�KTc����	ͱ�tD}��k>�{��A���ܽ|.�,�U��ě8"���uqH3����˃�-5.W�WYν�`p�#�s?��%	Ss��+���H[�8Q���W~	2ɛ�M��U����b	�	
.�+'�a���!!�A|4�/��I�d��y=�4��tx(�0�
h�tj�t엽1f�H�:�C�u�����`����^��c�k"����Р�vْ4z[���]�>@����'�:�q�ۀ�s��ӳ�oװ:te�Ao���v��ź&���h���> ̟��n��OΘI�Ȱ� ���jF.��M��p�[�����DG}��+��|G<��k�����!���G3�FO>n)=n6�S�)�d��{I�@��l狚c��Ί�-���A�� ���AF/R�š�4���V���|;��G�p�d�XŃ�'ﬂ��c
�5�5s��l�*��y�$��؅����+r��.��E�QkD���+I���F����jwc�r�[ƥ��Q6�����g�Ogno��fh�w�<;�n���b����� ���t����W�=�N�9e�>�Gz��.�a��V1���)��³� ��9 �Z�(����<	��2��Շ�@�U�=���L\�g�~��ʦ����}mJW;���_�l�g���:vG��.~�
��ӴdC��$&�#���	��Z���D��`*h��%�>sGA	���U\&��V%u�h/1� }��& FL����_�((X���W�Xs$�%�>4�DD"`X9ll_%SS<[6�����)@�]n�u��?YHS��SX�_��Ky�]�p��o$����X�a���
<X�A����B���82C��;����гU�p��Q�*�?��v�Y����[���}�YE�|��?G�ͦ��tk��9M�	o�<�� FL��,�{��`K���������sF�[�M趾I$]BB�[��y�-}u7�F+�PiP(�}9�M!�1D*>��8�n��sEQ�H�2ժ'u����{B�E��@��1��{t!B��F��a�5ɄZ�r�>�c�P��7�`��SkMu���N��������a���l�֖��T2�Ԉnȿq�����Wa�/"2�kp�5���Q���L�Y��9�o�t������{+���Jc�H���ݙ|v�Ͻ�d�3��E��l��7�����ܮ��"T��ޑ
�,X��FB��F�Ô *��ς�F�3Y�Q�p>����t�o�.��V2��qh����[�E(�@p�&C&v�d�Z4��;\���{[��;�n���6��~�,�匹��1��v>�n�(�%g:��@Z�"�T[I�X���d�TM��)�ry�3�uf2?�t�>M��q��,5�G�JJ��?�	-�	
E�)/�8�l�30txh<BU����.�Pj*�M��%�]i=�%/� �
�Y�\�8�͎T�B������m{*М��&�` ����+o��������N\�]X��]3ӣZ7��nۆf%s�a �X+����#�V34��?^П�ˀ\�M�Ɓp:��Wr
��`���V/�D�֧@�#���>2��H�W7�ϬR�����N/c�� t�����x�.��=p�{&窄�2��2{���ߤ���~�����ό��J(�=�m�8�a� Y�#���O��0@�@�/��	�3�4eQ7_o��1I�]q�f:����zt��:�Zk���{�k�ɾ̵��}N���$e ���HEj*���^�q�b�}tS�+�S��y'�C��� `�f�0��~A5��c�SoDЙan9AۤÎve�*E���4�
9�6m�It�A����8˙�$����:�������Q����2{nf���hw�I;� (5��y,����%�	��B����B4A��[���*Lo�����B+�R�;�� #kRE�d7Ȁ���&��91y�h�Ċ�u{��s2��~!������qO�c���fh���<���2�)�ᅅ�N6�k'{!�㎆�c�f�T�!�����>�+=v��]�\�8F��n]�|R�yo:�h]�7o���V���0���.6��;�v^��c�}"��Ҩ ��Хb�2�9�&�#�1eb���Lㅘv5��b�r(�B� uB
w���L{ܨme�{5�nPڣ��0�t��R����ux'�S�vP����k�DEw�Qu�>|����H�3����c�.E��2^Ό�yŘn����.�Ȕ�M���o`�]��.j�����mp�(�g�I���e ��>�W�@#��1������^��4M`�l�ĥ
��+�"��ޭ%!�p���q_Cd9� »_6a�d��؜y�f�����H��C��Ϋ'Z���gd��6l��,��rb����qm�q~�\�,�� k�Bw����yi� m��&��ARE���Q�X
#N
	G�¶<q�:f{��ڜ��V�W���o-o��$H8 ٛ�_������ ���������t�1B�5pj��Pl��rw�a_�<�H�T���ϰ8eX��[4喁��A�#_l�85
VԽ��b��㊣0�5��JXF�l6�zђ�@jB��i�y8��{�R�b)����.�[%�a͏���mo5��3�����	����] �v�j������(ơܞ�[j��z�_d�2g�����^g���v��t61������A��ݼP@��B5�r�z썄Hi}t2쿍ã0Hb��W�Va����	Bw�������G�<ó���~�X�)'�����FW.#D"rz�p΂�5����3}5�����h�OS��j��x7��%]g�>A�ղ+!渖$��&� �ⷘnr����ǒ��P5�v���9���~ ��:
�J�ˍ]Ts4+M�S�в6�i�� ������V\)ӛo@�1�#��7��,z����� {:��2�@��G��2BB��g���f; ����/�G��X,g�5Yv7{ayK�*����ݑ䉮���2�;X2)����s:�������o�Z�+Qi����}��8�B1�Lshs*��8)B����,��50&"��ym�	��@���\�c^���.�+cf�|~ȳ���?�(g�͹�������U&}�����q_,m�}��y�s�0 �y.��Z�o�u�
E���Y���0��s�M˯n�t@��L�4�=6��iK4~�{�
�-:zݰ�4����Zl� F8fm�:�,v?��#�I=�l�3*�˫ goΡk+�à5����L�G��P�\�'�(���/��m@��J

�8��c{�W �_8�Nc��}ʒ�^R��!�g��o�h��jB3B�FT��g�.F_w��������m�)�5j��ha�]�s��d�s+�@y^�ٲ�yD���-� |�s \UP7^��&�oҪ�?nlv�;����C�Ǫ�d�5��W4���6�3�Wx@H�Ģ+�0�*��nJ\jd` �\��`-��9���� eq����ք��l|#�)��y3���	� �s� GYa�>�ua�e�Y�A�T��|�6�~,s��"���I9����-�'S�-V_���LC��C�~	w�nm�����i����MW��Nv%�斗=�R�=�3���r=��N�kE�p�q�U{��=�l����#6y��{���+Q�z����n�/1�RO�ܢ�D�H`�K!I<T�6l�O�vu�^//W��>���E�ȶ5��3.�+��0��ֽ��_�`ya�?@��H��b��4Mƕ	�Yy/H�bq�!�Q��,t<��ٌO�t8��`�F}k�㡟�C��7��-�Ѷ��:iV�0K��؏y�4�$j<����N��Y�Q�ye�7��%C(��7�ߨ���{j����.4��]�X��NF��{ɘ���2^��(Yst{�~�v+y!�B?�|��!��%o$[Gd��.�+o�rĒ�� ��BIp�-r�5G�䛲Z��!S����}Kqz��Tn'g�Q�T���vx�a˅Dy���4`
C'?Ft�0Zz2��5�H�<`q����ù��8�}�����!#�@���u�R7ۓ�ԦR���g�H���=�����ZLb�yJ��sQ[�MQ�b�����Y��V�~]��>r���ɵ�Q�����O3�0"h��j�y��,������c��rG����sֶ �ĵ����q` �׌�Gߟ�h��R�}��b|�x釥�&li��o�z(��f�ˌ����e�����쇡�8�ҷ?f;�:����-q!Y/9�2�ڍ1$�5������t U�Գ�q.p��J
Z2�QMi�[����"��sm�0����cAĪ�D�J�D~�1��)l����z�u��Wi+����t�sn�V�fj������M�U����"me�����Yul1��<�!Y��I��l�?}y7�dB���H�� �B=�M�y5���Q�Q8o��-���&i���*�S�-ۑc�t>� �U���<�s����0B����a�vo��߶!�"�2 r+�X�y�Nݤ�iow��.�aY //��Ȫ^3 �Bj���T1OsIܳ��o�|����&u�-\�Q�j�i�
 pj��@��/��w��b����D��8��X�PX��z+���5���ʜ����b+�1ɸ�kc�$�NB����!#�wq�$���؍��WXL�%X��V�� n�@�	�yͬ&v����� ��-+��W%9Q{�k�> �V����*��mi{� &���>���D� "��9IY�TW��c���t���L��$��=4��k���¨��+N����L��,]�ĩC��yɌ;yǍ���x/|�����aKw�����yd��Ӗ�[0�&?�����s��U%�n]'�*էZ0��x�D0��o+���S�?ҭ�
i�]=��m}:B�Gc}�ꭲ,8<�f��'�GQ+M��X�2�n&�o�u[�I�1Sv(�'�	�n�� :���&]�u\\K�=�8���c}2��nX7zH���)�=:�i*�Lβ�֋�6c�1lkq�}�l(/k-�-���t�NTޯX���:u�2~��٘b���i�ǟFt�ԀZ�����lEoK���/��=\��&�>��ݤ]'&Ƙ{�.��2R_����O{~uk�"���Q�z�SgJȃv��Y��~����9�kW���`���h��M���fS���خ_����=�Т㯽��!7���ԍ�ձ|�T{]Q̟l��i�g����A��:1�\|%	P,�1����#MPT2-Dۡ��5����jJ�ee_ΒA�M��@#v��a�fd�ɵ#�aN�˴=�I�hw��|O}�Nn��1���񜣆�m�i\*+e�L7H���(�s�4o�x�B�`$^�_G2�C,�Ȁ�oN�8�ܾ U'�;tL�{kX���%A�
�L&����%��4��%���|0�:A��G߈e��ĩ5$&��� S�*p��2X��5~��� MŚ_�P}��}B�^�0��_g��3���##E��g�``����q���d�8I�,�T�����
1�4դ3�#a���C��bİo�Љ�!F�@���E��B�e��A/x��r|1ؚ��0���0C�BP��]���p��H�q�h���j���R���Ԍ3���ka�ׄ����rj�Y�^6!�c���C���z���r-+��R���/{���_����k�hж۸f�=)��y��Яɚ��A�2ww`�m�g�TdW�^8���f�S��t�۫�b�nM�1�o�0.���>�l������y�}<���`���U��^&j�ݔ�5=;�,��x�i�N��#$��G�L$5�Ĺ�0�@�c,��Y$E�#�&�5�v��	��]-���N�؅#r�������0�4�4�Ky�R��	��|>��"P~8p<�]����9��p})����5����8nI>F��tD�iv�2��_���~*���`�9�R�#7��J���@c�I�\w��5ڰ=,J�&�j�ի�l��2�KwTJ_l�3�[��ʂ�UK}��lP-m#��zk��PT�����ث0�J�ʷ�X�C����@T�T����|�J�l�	�tO�p�4�!U�����5+��� r S��?M�L� �H�	�H_��/�JN��IFmz�8�Vf@�z�1���/m��B�sʙC�-�����Z�@;k�k�\t�s�s-�%����)����3���8hmKn�Tح|K�1��O�#�[4K��l���wj�t����n�(��8�סa,^WÃ��3$4/�ϙBν��$;u3�֊�t�?ݧ�/R,)[��D��P����"u�7T��F{+_^�����?�X-�)	�c�:O�=�1���ɔa�|�rz4�)��p�����V�<��t�K�R/p�A<N�;gw|��9l`3��CG�j�QjI��{��SH�]����,��u	�)Ј����U�7���X�:��#���`>[�q��y�B������Qzs$
��![K2��c���Z�G��;$�hjט[#D��h��k�.=x����9�>l]���jʫ�>�:I)�d�D��9^��g�శ����i{;��k���p�d�x2�.Բ˯z�����>������W�T�Uv/�Ʀ N�W�M ^W���A0cRFՉd/+�.2����#���Y䆢>�L�[�ld��p�U�Y�J��x�_���6(�rO���[��'Q��D�ʌ���~���]�
��������1�$ε�q�"q���L{8�mnA_�H��^cg)��>KE»��Y��	��`����?a�� �5�p��WsE�YHq ^��a?c�O�?Jn��_�:6�]� 5^�t�E�S
�h�WA��	�U@�� K�^g*��!<K�L[{�� p��b�]�H�q���;U�;���-/�P­8Ju�l�ja;<H#��S�����)�Z)�}d��� ��/]��1���@yME��@L�p�b�`�P�F�
$'�K�S��FNXy��m4	{�� ���:�7/,�du)G�����`�{=���`Oeē�.�BB�-�!����@i��k��	�TEW��)����D�}��V��1Q9*������|ü�a����g� >Q�I ���dK!���1F���a{�%�Z�XO��e����E�I����l'�Jď���D|�3^�֩:��g�q�@��H��oV���$�4Ay�elE S�E��D��h���yV�Wk*�[��h�0��%ٲ�qЮ�2�$*�הbZ犏�Rg�d��~iU<����C!���FC�-�D���,����Jr)��tT@�V�x�vv[�z4�oV�̸\��|���H�0�e��:��0I3Z�uo+C��b}�9��~��#�F5^*/s��E�p|��$9'!���砡�ˤھӬ�9����]�$��5M
���c��i\��>���'kG�E@�Y/
Sә����_l��r��t�`�L=׼,%t�8�^�������ƀBY��S^D"�W/y�cc��s`�u��"�	L:�E~�������)~�"�Z���1�!�����"�D+z�O�m6l�cFt����7�֎!���\q3�$+�V��ZIUkw��}�T����@4��1VQ*c��c�<�=a����M�*&� ���5�B5S�:�X�u��2��{�ˍZ��ҡ�s~��s�p�v���"�Z�����m5W9fu>�o��"�|&|�Ѧ�Y;t�ܱ�`���	g`��� Q �[�!E�8����ހ|����2� ���v��Rjj�T������z�g�ض�����N�F��O�!�~�=�:���Ê�a�0�˾�6���bL�k�+�)<c�� }I������~�rN�����k����7.CW��u�g�uJ�/����&��֑t;��Z+:f��Tn)�Ls6�d&
'��L �i� ���/Cw�3���o23�%�h�"%@�E�z�P4|�'���Q�+F瞂Ĵ(��!(��a�)+Q{���6!/�]�Bl'��ĸw��ϫ٦$�	����@w�&7����*m�{~�j���x�Uά���.�	�Y��Hے�l�M�!Nno����wo+��}U�W�m�a�NasH�$��4�~7��~���Ǹ�7o�Ls.��e	0ћ�)互�$S�&�4��n��` o�#�s!.v���`]��]D"$G{{!��]G�g/����X2����x�|���,����D�8tӽN�0<B���0OD|�Є���o� �f��?�zC��/�	cּ��}�H�NB�Ih��l�sq+ �G0l����)q�~�_���hZb�ri��m_(�u��5+YI����8�h���<��eه;Ŝf*
��~ z�3�6�cm���_?�,j86;H��C �*�>uR���{�*h��ڙ�*�X~m%��P�0u:�=?�S�+�ob	��{� (s�� g�5c�(	!H�o�;BGe�Z�5���y \y�{�v��PH�9�7=���e`�eE�nd�i��%W�����6�j���y��u-"�%/�Q�����0m��]�ݡ%����e{~>|�|:�FY�&��M��ҥc%����IM��5Y@�H��ɣ�c����XI��~f�C�ϵ����Q'���W�u#�Z��_4z��VܼwhrW��5��^D�����u�u'��<�{z@�l�$>�o@��}�71o(��嗒%�[;��>�x+N]b!ܴ�Q�9ҜDU}�n0>��O>�V��V��
Ўٺ���[���;��fl�LT�ce^�����CgvD�T��������h�����͡ZH??����"����W�� ��9� 7�	�?S�.T���`W��_�	/c\�2��C�}7����j�N�%&g�\ZNҝ�5�
1�b?�fn��O�5Υ|�q
���Δ{�"��x�揬7�B~NDC����,�yo����
�@���w ��8�����A�7@K�*�!�o���T�7�wn�����ם��6��[�Ϭ��[9�O,���%$ս�b��#�2�C�[���iE7�(���\b�"����dd���e�.�����C*���J�7��U�ش���3^AwNsu�xc�H�YS�yጉGyda�
�y���~���3p��nh/�+�W_�����AW�
N�� ��F�!�?�yT�� ��Lҍ� ��A�Qjd��;�rq�ak%�N6i̔�-Iv��Èq�0WE6������3L�6D����3�@������_yڏr}�#)�|�^z ŶR�|U���W�`Ѓ苈2ٰ15��A��=P�bc)]:����!��(��|+�̧D5ݨ��Mp�y�Sos�L�v�I����tu�2�8���E���0��*�Ҷ�#�Z�����ٵAΙa�Wt���͉��t�v�Zqp�.�~($fW������׈ڝ�-e>i��`���%����HU��!,�9�Lig�HF�&?���势7�?=�JS;l�����6l����যBv��ރ��8�;2,����.�b���t�z:���Qq�-N�@-&�=m뿾A�yg=C�e�?�1��h	�ov@6ΐ�t	��ȺWȻ>��G���#�&Pd����3�`A\��y#�� )δ�@�5��[!��t/*��S�������p.$ZA|�T�Ȋ�i[p���8��A��`�T�x_�$���P�`����
�l����;z�j@yKX�.50� ��>�wy4��j�[�������p(�#��u�om2/)?\y����T����g҅L���`��S���V�����(9����+H�L9�F���b�^-̌��=�иJ�'W��yjU�S�y�(Af8v���%[Q�a<�)u߶7�K�ù6��kꎭ��+qR��ͤca�g���\���y��A�Nj
�I-�A��@��_R�,������Rm��!$L�ߺDϨ:%����A�^�>��|�
#ra�c�䲠��f��,E{u]�
�xͣQ�:��o�����V�P�u}��?�yc4�g�0&��}i�b�W�"C��:o�\�ۧ4��L�X�J�B�p�;�.��6�}n��zu���/R\W�zt���Ji�?:�ϱe����S�\��~@c�0�^�]9)���1A\w�	�Ъ�=�᰸<���F  �+}z�ӜdƔ�f٢�l������6������eygМBs����^K(����ZēF���3���y��G�]W�躂�BlISD���[�c�Y�uV��0bX�abP���*1��tW��߅J*�4���}�K;��d ���E����!M�����-�*�v2��_�׹@ׇH�ޯ ��Y(�S#��T�&�V$��ڷ�ը]�����2 b��W�c7���c�G��bVKjl+t���éf9F}чGi`�SzH�񉏰[�<_s򎢐�(��Z�syD��T��,�;�Y����5?CL�={�4a*���O}��c���H�"|
������'�z�����ʕ&�|.�����O�}>>����n�of�7sN����J����wL��Asť]c"g�)���(}��0˱0/��3а��L=�Hs?'Q��pRI{�qB3̒^1�xXzb'�ۧ�k��%_v�$��.Q֛~8�B�hp��TV,�qm��/:D�U|S�7d�%f����t���r;m�4�a��mf�1V^�P�j_��Nߨٔ�F���l��{��Y��u�,_���9���ATIS%���;ae�R���8^�/ �:+׶d�V����$B�Y��Y�����P�!zr%��"������S���QvB}r߲���U�"�g��6	g�}ك(]����O�JD������+[e@�eOz{Bt�2jP׬�����������0��rf�uO_:���_��ww)y�l�)a������г3��bp��������$�<�����OLH[�jZ��&X�f����5�B�'�h;�Yh�1�=�U��R]�N$��O���!w��ߛ�0���/��A_hE���U�����뷍тC�q�f|�,�/	�oqn��C��-\n�^'��4��oXwSo4㓖Ǆ�EhѬ�>���n�� ��_~��]M^���^R,���a�]����l�e��m\;����\��9(
����m~ҍG_e�$a$��z/[�c-��e�_m��"��(l� Y��M�z����k^І�B�s�*@�� �x��_?N�a"<����z폷MT'�Y,�ƽ4�*��w�@¼�zD4����̬�:��.4���g������u��Ց�hl��Q2��8jC���X���e�FB���B���/�����ޫm�0xɾP<2��zD�5�?��i�]}]?����6��<_AYȍ��,)=�-�s�����$�" �!��?D��<��܀|�N]M�ӥR~R-$��e�sԇ�0�R�
~�TW���P��
�jW2�v�E�CE�D�}�!%�� 7���������'D_ح�����#;�EZJ^��KYKb9�
v˰�Ұ���e�G���}u�
��ν�[�|��� �uyQ�c"*���t}�?��ð�7"����5�g��$bڨC�^���n|z�!�z�Ͽ�`u��Z<��L��S8��B��0��yu'�Ƹ���b�g���"�R� ��7������udm���)i��n�o�F�dO	�V0�n���1���s�⬣bp1��g=7�~o��V�RR>�S^�vIʝ���g%���/�J��3���v�mX�kC��|��E�-�S�%��XA�J�0�鰚��2�]Ʌ|ݺ1�[�;�#���xCJ­r�3�/c=åQe���*�d�w������:V1���u�w��bp��B�?���"-
I� p.އ3c�$����:�Ğ�`X�����x���k��}�{kyƝ���sk�|�	���a)@ԋ�{��mQ�ןD�=���᪯9�-����F3}$�Ɇ:ݩ�tb6��"��ҍ��z����owPj�\�����;������T֓Vp��}y�6ۨ黨���H�3����+��c�x�Ƀ� ����De�0$i�(�G�4��h�aO֨ ��Y�{qˊ@o���Z�~�b�U�{�����R��7��������9F�_%m���s���wp�?(d7�8�w����g��I��w���mz�2-������-�4�����r���<2UP�ES����J�~�m
��X\Qs:!���e}���Y�(-��Y�*��,h<j�҄pZ'�6q�PLҠ��ɫS�d��Paٚ���AnH� �g���T��U�S1��[ZE��'62�����j,L�ް<�`C�Y�16��� �(��HJ��m����z�����d���b+$��B+�}�a���U'����X+�ű��&�T->���B�QQ��U�ͭ��E�
���Z޺�j<�"�ީ�{5���!�6rަ�S��*��ۥ\(��\�SG��y���4I��v�ޅO2���\�ëvBk��G(wu�.���86�*���+ү������"M��b�Â;r1��R)5-m�ԍ��b���&&����-���{,E��v����6q�4��e�<e�y��F~#�rW����OH���]�h�P1@w�S�l7[n�=��|*�Fю�ٲ�}�s�I�@��x����yZI�����X �]���i̱�ഗ|ؐٗ�!\���_���=��t
�){O��_#n.F��ɕ�!x!eib�t#1��:Jg����f�LA �=�Lc);��;�S-Ix}{d�-��x��P�J������_�V���}K1aPg��z��{���9����O�HU��|����]<�vI^�a]8�g�wB�%\<aIĻrV`��f��;��g+�rQv���G�>3\bR\u.>B��<A�yã�0Ԁ�Z6()	�
�)�A鄜�:���~��R�̅��]}r�M#GL���aV�)Л��$�M�f9������ª�ŏ�3 ݅A���2�7�
t��f�*��|:6�������ۣc�'=����:����� �/�C��3�ڥ+A<��/�՜܆S�!�[�(�L���U5�>���-�P�C���I|-㘆�B�Ng���*iF5$��<��Xh�'B
��yni�[�)�b��w�TB]��$�Z ��T� �ߍ��=5� �}~}�8�J��ThO�؅k	ݠ�bV�V���Rg��.u�'n�#��i��^z��4�JϟY����U��j]Y`E%U�;��(�����Y)$:���@�_H�q30]l[���]d���U�%�M1pݻ �C���	@I�?��tcUw��kJ����V%���+�������6��ʏ�`ȡ�p��M>0�C����xS�p�/����
߱�W?��k���u3�B$<�v��;���(-��T�<��'%����%��؆��ɿ�ji0�o��í����Z%��)��a���M�){o5��Y:e�?��2��l/5� �Q�k)�x��].������=O�m�ɲ�t39����$t��N�5�RnTf(��P���,b��#�&������V����x,�0mWs�y���$7v��d�Z	U���w��D��m�/����GRt�]þ��	�~���jÍ�V0W���I؋
tQ�J��G��WsJ�� ���ſ���
�ac:�:�x�>`]CYˍ:7�n,8|8�?�b�m�|)�G8&GAx����ծj��4���Sr�� �vǌ���§�� � �V����?
�l�Lo�}h<"yۏuĒ�27���$�k��}�u�(FFj�/�)0������s�|Ʌ�*����ߤ�)�x]R��'N��I`"�5�G<�cv�ס�#��|(�X��m"�Q�q��B����B�i�V>���$1
��T�aj�����0���W9G�wsYԚ���%}k���:��r�C3 �ڠ] ��^¼�}la<2��D����1t?۠̊Y�� 
�|LR��I�"��fvFg]J�ĉ��>��[y��S�C�>���O�`�s�aX[Sn)�9)2��YE�rL,<ԩ]Q��i�ȞT���8q���9�Α��Vi� � i��{���c 6�����S6L"��`��$�q���.*�Kl⬳(5�6Ieon�K�O��T9�e�����J� ��mwP���, H�E��R�����BN�����\�2��zS��X#�}Hy#�h�>������fGdn����A?���4=�y�o(��2k�q"9��Z���/�m֬�@�ڔd�e=���g��m�P7Yw.�!R�d���n��0f����������9�b����� )/�)k�X��E�-�Ăsm��U�8�Z��{��7O���f�� Qդ�X*D1��y�Uk���H\�Jj�=�m_��x�L!������
;��C.s���|��)��W��g*���9���G�W�ˌ���X�i��D�})5/� H5+LHDM��_V͐���@��X�JB�b���'��M�
h����ݺ��Q�������?����	��so�D9�xY���+�U���g+z�����ȋW��ܧ���W/tp���hzaN�^1���B������s8o����{��%ߌk	�O��+m���D��3P&)�v��9>mk߅�N}��Ʒ��pJ1�Os���8M�ԍ�d&Ylcn�>5.m�Y����잷�Q�����q�3��j���F�Q�`���;��TH;�.X̧Fu�us�F�)��N����2�P��>��k�RQ5ޣ���<���MW�I���
�H�qRŠ(��Ur��FI���'�3c�Sk���	0-��Cr�E���G<߸���yH��gL�ma�U���v|ԯjYrˠvd�J�X.I��#t��z�(*�6QCg3m��1~��|����P+>'�^ؑ�ි��GX=�z
g~��ny��8��%�՘��rSP��</>�^�S��%,��ҧ?q��;L6��QwK'�N�-
�����^o��M<�}Q��VP�SH��$O���I�斃�%��rMm�/�S�\�\?f4�Wm�[(K4����[LLQ}�A+���E3
�y���̼TRb�Ѱ��o�`à*��=��X��-��;������1g�tܒ(�x�a����S;�����A]}����S�`�t#�&5�Y��O�jF yqb��}��u�����y��I��|�t[G��.�S���\�l)[G����үۜ"ES`�fm�ak�m�+���~��Z�Dq�E�Sgז����ˁW���:��,?�f?T��8c����ܝ_.���L�{dC��Z\�bȗ,X ~6���f�Y^�����;���2@d,��$~�������s��ُLY��W��+r�C�Hzv\�J� �rI}�)?\R��֙��4��s��l����Y��-f e� �����
j�lt���]<����S��T+���9��_��ķ@�GyR�#lre�������i����lـG���X{��{����
:Cn1=z�A��?'ӷ��y�7��X1�oE;���U�j����8>���y=���"�u�N]4��T���d��e�<Yl~�A����W��Of��⊿�m��H�Ki9�/ h��6>ۘ]���R�5|jb._�,b~����U�f����l�<4� :^�}����2:N����mQ��L��qI�m��~�k4&c�!��a�Ͳ7cgR>X����G�2�լO�ʝA�(����ym0�d�:�e�r�b���B��!��
�o�L�at��z&NB���̥9Y��*Ң[Ix�7x�Uj>J��0AY�.q
lWضH���ȷ����5I�^x����%�<Є���<@}TA�L�Gn4Έ��S�S� �qG�K��Sm���|4�GԌ����u�O��XЏ2SB D�5���������	���8��\B��%Dr�dP6�e�����r��W��,+��{i�Zo�,a���N+������W����B.&�ާc�6�
|������\)�]�Qǧ���-i����z~
_ɱo?4C|BEW�մR�#����+����D�/d'i���ּ��" #15Yͯ��-%��qw>��ר��d�i7�~�tP0 ���M��&�&���}�e�cx"K%�f�@	�.E��";�{��8�
^F5�e�����>T�%��]��\��W�ZE�t���N]3�r_������OY��F���D,�E&��2,�B�&-k݁8r��ޙ�h4]u�[�w�����H�bh��<=;|3�g�5(����m# ��������N�3sQ� {\���\�����
|�j�Ϗ����TU�����؊��-V�WLaw���{Z��)�#N?_bk�K�=;�zw��
tm��6:Kj䦉�ӂ[d��.�Gd�8>�:�bq�G@�I���ȪL��~��s� 2.�d�W�90��<���g)�u2�ͦ�"=�C�塧��0�E5��M��9W�u�-o#93�i#�Lǒ��}��.���v�=s3���M�E�������0�K��������Xj~'��hN��c,�(}�c�����?F�~�a����N�&�.��\��ؤ*��(C����fN,O�9��G�y�&q_�y���"������G�~��OYj��ƜN{��})
�R�Uj�Ks=�xS�O�+g�4	ٕ������)��LX�Mw�}�k�׸���q޳	�%�Q�=�)�y'<>|�و�*V�	1Xr����m�Ӿ�L��������m�ʈ�Ws��.)�@'��O̥�h�:�ܬǪ��%��j�Y�[ft�(f:v��C�^��A���-HC�>��G�ԟ"��LHE4�J�!e��õԱ�0��]�~��4;��<����]��n��rJv�L
�Q�0M��]�߭�`�9��N� �zSx���̙5G�ۉ=:S��sQ@�Vs�"Y0k�%qA��Φ����^Zl��}g��b�np�Zd�f���;���Xᗂp�*ǽ�$����b5��*�2�	)b�8���B:D�+Qz�����"�rc=[�vU4�V�v��L�o/��A��h����Q�c���fw E���# ق_寰����L�e)I]�
����� �y^َ#�HtC��^b�<;d�#�'v�5���!�$w8ra�I����LېicT[;��9F�8�&~���%��EqX�CHⅱR4g���&̍5����O���b"����W��;I��,5m<�{����_G�����e���谎B�-U�o�|bZ���.��icۈ~�0��fu7B���0`���3�|ȥ;�!-� (�I2dUS�W�:Vh>z��_��.[������Δ'��by���8h(/c�A�̗��*Lch9k��zй�kn��?�Ʋ-�xA��(��T���<Ek�7�������<2��me�CW
�Ƀ�V�މ�Ǚ�gY����<;%g�l�P�7�g����ֹ��3ր{bz|]R�����=ԓ���L����j�`&� 
�����dі�� �f�=s�F�:��&qZ�:�Ң��wi�T*�Rnd55	\L��4�a�11 ��uG��>	�kED�K#���XR.��>�iý�/7j��zꚗ�/�:���C���ݝ� 
� G}�:AO_Xe�ZKv��O�}�y����� �/9m�Yݜ%>(�H�\U�p��|��Һ������Xh�0����E�Rt��pcRf�w�rv7e�5ѿ+U/��B��T(�t_g��v`l&3���
�9�՘7�=�p��D[~*���)d�ilC�N���N^�
m�݅M� {�o��� ��d��\S^ �X
w��lDq|�-��T�+e�n��w9$�{�+Zܜ&�|TÛ6�%�+�l��NQ�q�u�ó[�J��^-�����:�k�H���B��Zyqh�����\��!�����J=S7�&3��n0�!�P�+���� mJ���ysd=�*�Y�F�i�E2��gMG��3v��'�2A�$�a_� ���Z��V:M9
��!5PJ��/���QEi=� ���($zQN�r�'�x�#ڜ�D���9!+θ񪱙�SP�#���j�+1�>��T8�lk!>4 a��9-E�Y'c6Zל��Y��8L�ܭ��J��~�4�G�`{�S�D���Ηc_b��i!��᳻�t�i���$f�C�E$e@��=#ߐ&ԅR�K�S���:Jq�&nf������ヽz,�-{� 1�q2���V�ɞڰ	?���0�*�c��p|cٕ�w�`o'�HL���|;R�?�娴�YW��mIӌ�y�q�A2������}�l��ޣ[o���3�E����h>�{��e �ƒ��n�F��ِ2>H�x�B�*cIov}g��sڪ]���C�>Ɩ�8���-0�h5� f�W�����PGg�I�M�(�$y��sHf��7�~K��X˘�p�x����i7s%x�۶ͦ��t��$u���xa�MU�x!�̈́k���Sf�,r�,z�2�t9�J�.Ʋ���
2?B�����*i���EDG�t��NJ����)ä��������M���xA�?q�ݍm�|1��K�&`��ka_y����m��Ϩ\�N¯pT&��$����Z��	�pj�nvr����_�'�.� -�Q̲�����累i2��J�SN�n�\�R�,��A/��Î��?��U�r�s[��T+��5���O%��t�3��A�h�P �Q��sP����5����x���5�|޻�A>�VG
�Eh���_�
��%OO�3��Ni)��m}C���Ԁ���4&��)��Ng�E����D�56Z1=�a����������ؠ�@����Qed5J���IW�qvNY�\�2�!�V�̌x%��x���/Y)c��m���<38q�����0ޣ�!	��x�'�X�2p�8u#j��XU���rR0�����H{�Y6�%d�@��g���2V����grZ�e�N�١�A�vYO �Gk��jz�Șs�Q%��˛���}LI��u�<��&Xr����Hn"��G��Sj�����<�l�/(2a��j@1�	��w�=��)��ޙ��o�2)|�H)�^(��p��nY�痪���:�z�Aw��*`��IGS��n%���If+a�Tk��%��6V�[\m)��h*�1��IAB���p���Pޅ�i�E�C�k�?o�ե�	MZKMб)�'E��&��h1�Ԭ��!x���n!��'�([3& �}��Ϡ:W���3sӟ5g��^a��G
C����~�1}|��n�� ,����\7��$9��'|P� s�}����P~F�o��%��P-��=/rJ�&jh���/�͢��7��xlHn�9r�O�ʸ��������K�},���x�Pi4Q�k5	p��^�h��7�ɘ�7�B-㌵��g���̆;�� �pbK����؜gX����
��F�ɘ���XӠ�Xm'+�v݀WG��Vl�
j�ө�h��5	���/����A�bR�
C�ux{�'g�w�B�1i�d�Nd	�Ү�\Kj�S�j�cT�a�ԲԂ�A�>�T�m�W��p����]��b	�s�>�:�8�߭iZکS[��y)P�����.�j�d��6���⿥6�ߋ�5DE��L�0��d�O���"n.nv�_m�+����Ɗ{L	q�α���.l4G[����'%"�\1m���Ґ���ך��+�H���Ǡ[���dF�X�N�I���z���~Ȟ|\j2Mք�n�	����	WP랸�@ ¦�Cğn>C��Fo���B�c%�Z�h�;O�߽+� ��d��<<��Ρ7�	�L{��E��R���'c�b�C����=Ty���%�V����a<_��7D�pϢ���k+U�ƥ�eZs�o��eUl��k�:��� d���s8T<UP�>RD�5����4�Y�p���j�ZxA�''��"8A3�ߘa�Vn�j�m?7�&��3fz��D}�k]�t�D�E�n�f��V��?�}u¥�!����\�z*��"T�1_]mO���H��/�O~H��Q�I��sk����I&@(���b/&�?v���J>��FG�d�~���_��`7C��x�/�+
���A�,Q��S~:��p�������i�ζ06��O���+)��b�䅅HĽH�D���J�)�
.�\~�wm�e�#f�P��2@sk��	�х`���b�0��ə���V�=y+�o$��K:l��mI\Nmr]����&`f�� �(���Ev\�]�b�W��%��F��(�fY�� � f����7��hP�.3��F�F��b����2́��^��^��sHU�-YÆl>���>�S�����GN�֓�N���Q ��&�d�fY�G�6]B�i��������y��z�uS�YJ��rz!�&��Q>}�y@�fBp;o�����=
yV���VG����L�HK�����E-z*3 k���5��y0h���_"-��Y�y���V`�Y˓3ة����C�X��L_*)23��Hʶ��޺Н����[J]�����?a�y�sE�ҫ�G��x�ڗ����y��>��D�Z��-av�VK,։p��ŶQ�ģ�)|s}d�233�)L)��Clq�Ɖ�}��J�d��m�̣WE���Qp�S�	p��l��ݟ�w���e�O�N��vd��7g���M8�Ó�Ma�Y���xcɶ��'�=�)(�
�:љ&�).�!U�q�LY�U)Dq3f6��k0��\��LJ�R�nښ4Q�o4\�Ȑ��#�l�a�w!�һ�]rzm�d
�s�R��������J�Z�?޽�Z^F&�T����-� �Lu���
�9tȒ<�;ڝ %x.*��˵8l��K���|D����dE���N�A28S'c`֨�#[�=�(	�T �
@��(BO�ɺx���I�
W����.����7���ZR���U��@� &f�f�ڦ~�M^3I�K�X�=�����.&�f�8�X%���>n]�SP���~w��H߃q�Ψd���!j���W���m׾��^fW�!�(�i�K�)R�`��2]���ݷ�y{~]�����X-�|\���++�I��vVі���!����0����E*=4�C����l�z�����+h�q��	W��FO�.7���E3��]��3�bbKFٜ=�?SA"j���(?����]��:��)y#��]�M������S��1!ҁim�����5����"����n�������plW'ݷ�;���v�xl}����^��,�������б���s�.q�uc�.��{�ǅp2Z�����¦E�ɪPWL*�<�:{z��W4��������z�C�<��[�����^�K;Z:(�%�+Ս���Aa�3�R͓5�()�M�'*���)?�
��ֱ�C�]�Z�i��i���u��Hc��j-<e��� ����Jȸ�""=L�[� r�8�ٶ�![���2����_�;%\��_�HI�	1Ot���[b����N�D�e,OG�{v�B�nF��#p�mi��S%6��RժL�Z�������vfі��s\��	8ZI,��l ��ˤz����\8K�C��ݤt�$N�|bBd��?��'�3�H���4��"��QNx��jcg�H �ye栎o����{�Rgx4W���"q���Vg�W�_w}
ኬ�/U��:`���&��wְZ�H9�=:I�*����Y���3Å��r�P�Y���.�%#as��Ѻb꿟Zcϊ��<�j`��Q]`��L��7X�i $��'���6�w���k\��	����[�D����-�ׂ0)d2ycu`(����IVn���|��\|:ӘS����'�c�T�C�����;7y� S��&�x[��',TT�x����[+6�PuҔ��`��U!X#.�<���?��Aˡ��}�?�N�/�������������;lm�B�~�EA���,�wj?��Ũ�r9m�7�]�$j�x��֊Ti�ߜ�?q��%����OƾYNK��͊z"���'r��&����r���r4��#wW�l�͂��V����Ko�]��-���V���$�x���}�Н�����;�ȃ�������J�?u�i��<�+h�	�_�J��Ђ���O��8#�;��ÍDkf2�KR����em�^���GXm�&mh�$Z'o}_f���H��<�r}�6)۝����a��І:��r�v!���=��^�\��c��fe�x5��V���x�wtU��ZD����&2����<�P&��25m$Aѱa�x�� 噸:��7��
,W�It`��8���7��0�
8�Kz�}�co�鎟4�HK	��.�b��-��s
3�GE��=>R��z����ˁ�(l��?m�D�7,�(�x1�_"���C*j���������(/T��$n0Uп�{����d����º�v������Eu�8ɝ��(��z28<�2K/7l��Uc($7&���%����3W�� ����꯰��fSj�L`�Q��'�xC����t�͙��a�Ϻ`F��	,_��ߪ5��ހ���"�</H�og��՞���M�����zY��"i�D�hoyb=����� 6�4���_E�U �9����2����t�jx�2�Lӟ���-N���OOx	6�L�����]�NV��y?9:�w�P�b��{@�smm��<�.�f:IG�vj�=��������pk�K����O�+�?qxi���?�n��>�ٹ�2.�!�P25����H�Ej�
.�)2�.��\��rKP!���9?e�,�n$��|�7�.qAf;tl��c��+��K�'jÌ�n�Gi��K��Q���f8G�O��z�_�ku!��J�zǟ�+v%����1�(���"ȹ��{����M�q�8�ώ��UB�-��1�����E\�%Wb�6;�gp��XS� �N�\%����\����b�+�?�^�oF�	�������sF�C+O���q.\�|k��^�2)䵇�����=������~���8�%E~M�|ˏ�ꅎ��% ��M/�?G�BmT�=*���H�?" �)��? ��_]�T���H���l�h�&���h�k~*?��>IȺ�X���D��)3�`y:So��k�;�T�֝�<�Q;`��d.���`hP���׻��A*3<g6�i�6��b�e�g�ק&����C"����u�V�Ap���L��x=f	qZ��w��bw$���! }���0��'HG!T��:ڣ�ĸ��P����h/�k���x�����r��z5���D�JT�4@pԌi�{c2"�=��,k�g'��+�4+���Z̟��n��Ì��PG�g2��3�AƲ5�oq'�;��?����~$D�,����it����-u.��UH��+�]{Z}�y��İ���h,�#x�,Ob����>�~�QZw��@�ez�9�^��5h�wM7��72f�2r�I���=��)�}	A�	Κ�7W���~F/��r+'T%��pJ3��VͻϞd()�����^�����T�h�:��N)�����!���%i(8���~��ц:������h�ȏ��c��	�K���n����ň��a�#�e;���2m_z���H���Q�]�K������-:��m�hr\&^	c0Q��ё����g��$�:����(H����|fb7��=���E��
H�qM�)AY��y��M��c�pL���.� S���nG���
���J{����LYI-$�L���&3,�����Nh�P�6��6�������F��+���7sWS�=Rvu؞��<2�`Y�96p�=�e��<{έ>v��#UP&Z�^D������=q����He������I�*���y�1ǉl8/t�D�(4E];�O涃�4�r����/��L��P����}0Y����)TdT�P��ˋHQ��L�i��{����x:e߂]��`� V�$3�ʺ�R�O%moܼ��}�](���[�k� �0�r#���r��90>��G���ӡE�<ё	~�;P�V�*Cذs�e�Q!�O�Lk��	R��]�xƸ�U��Q?!0������Z�&;8�����v��j�K�N���E�z1`l��u%�d6$���a�t�����f.��ۭz��bw�@R��-(htD�����vUt79���������W}ÏN�x��h���T�*Ю�xv.g2(���K�*s���mK�wDT�/�̓|J^�3���%V�?9ٶj������[�)g�I���t����Is�	��h��FŦS����T rɚ�#�f#��
I������$�e��.h"iL�*�t��4�q������	=�l�H��t��ǋ�X�d�،�`�BfR�A3��LZ���ذ;�"� � �t��(<��O6!���p)adKܻX�l�qDխ����0�+"��Z�A	��X��v[�J`����[����B �F��`��@԰��x��鄉��yr8ݚt���Vݞ����qIf��\�A5���+���I&�=���:�:ɩ)4+q�|�S<w`����G�&��W�t�il{�ΈJ�|{�c�0\�
ϔ��us�����y�"�v�~^Q��7E�̼��a�R�I@1��]5Bs^'������ו{��}�������ij�Ưd�F�� C7�oDB��\5�)S�Y\OS`K�V�.�Z2軮�Dia��5Ĩz֩��oV&�3��#.�  ��o�?�u ���X��� �c.�N��9[��UW@ҭ��p������o����8"=�����B����=L�x9���>�*U������g���ʢxA����u��2P���<\����vH�9D)��UD}�zT��3�~�~K<,3�)��S��t_�*��́M�a�w6���\��VϢ�ƅ�S\^��bL}��� ��Gd�1�"6�)�]���|�2ٯ�u����_��vB���A��2}*Yۄ�I��7�YR�\H���S��?�d�CyEiDNZ�%M������|�D��S&!�.�j`Z��~�ѥ}�,W�-*Ve Y�	]tl|��R��I�ȟVb�?�$�}w\,n�!�6�Ya���`����#fY1�9�
��Vкs5V6�ೋ^Ɵ�5��'���yCך�܆�A8%*L��3��X�/�@��m˩��;�a��G@8�_�{��B��kR��X�+7�%�ac�82;^xY"�<�|���Cu���X�6w��)��&�h׮�ٲT���ͯ�y��P�u7�Ђr-��<�K�C��KS �
�*��lb�;C�Zs��Ra�^�� �jω_��-�;`Yvd(<����5���<gy��Ě�� e���gJ��S�^� |��� ���}��q��=���z��Z�����B�sސ�<�_hv���<i_��˂�o�2�>a9�4��[��e��HHU�cA�/z,\bB6����� �bAW4@�pS�')މ'9���zg0?W�؞���P<�2�±��i��gj�b;M)֛�G
Þ�c4�B=��H�V ���r��{�+����q6B���SP�L�N�T����s�eyj��BP�����kH��G���0�j`v77mș{:�E!�U�i�$"2�� �)|$�z�>%�ROƍ��}���� ���db�2���kAg���n'��)7E��c�E�"�j�6�دbdYS�c	\����{`�F��똅J<	TЋ�
� ۷BV�������o�4��J�u�@��3X����,0\��k�ƒt<�6����_�,1f��P�P����b�����;Bv�_7�n��ðh���I���7*���'c�FE�xbXK��)�kȋ���}%b0�Lh���E�81m�4x<�s�3N�ǆ�㉪�����rm���2�h�dd�;xa�L:���C78�Z_�u�=�FmA!���J�?��B��*��DxlhE�-&���s�b~�oO�z����/�sw3�\�j�tz8$=rpE��j�n�e0����H���;D�>�K{)�J������5���SeL{��Y��Έ
_F��y��0p�� m%�T���0�>Hʯ]&�T/b24�L��[����Zic�D.
��;y�2�	r���i?��ꛜ�R���͂UU82����*bx��h;E;�jq��V�������	��\�"���7�|"��v�l�Μo^�]8=p\[j0�ӭ2�:�>�p�Lʨ��d��C�/�	�
x�f���F5��vM-_~<%b��BA�ա�`�i���.����Gl�Být��]ez��~��IT��8IV��L�|#�uZH,wbDA�Ҧ5{N���ߒ2��T�T��f�g�""��3<qɸ"A^7%��O�q1�� ��'��Ljz(V���eE�<����&C�Q���_��t���`�] _5�/��� �W���Mf�y��\N����E
O�P���!���k�ѣ�6�� 3�;�xyB��K�=��;U��F��w׵���gV��q���-ّ��xa��!�{¸��#������|������>�	gZ�/x"'���
�Z()��-q���R��n	3m�IZ��p�=
��A)�&��+� ��lN��qi�cbyAsDW"���K�'TkvX� �)I�M;�#����
h��H����r:��D��~L�Q�k[�Vk�$�Y��֓���-�AD=W��O]Pj�opș�7������Ok-Uo�e�`{�=��͞S\�Q8�]�!����<�^���j��-�O���l�+m��E�s�=y�p��M� G�#��AVDm�A������|��z�T-���4D��97�L �s�:\Q��/t��HaR�X�%�$�.-�������X_/��r{9o��I�)�}�+aA��+Eh��>���D�x�ۖ�ZO�}�,/�1-�dY�dU¨�(�o�?q�qo �N����7�i��8��g�z[LHu�ڧ�+b�;�
lM�G�>O�v���e.���Pبaeib���a��V�����	q�C��_����ꆱ�]ڊh�d7Zd2�j`���#��N��*V��/l�͢/a�Lv�F9-��I5��>X�8���f�v��fc��ìE�s����!Z�-K�UT��u����H	~��u�ݺ|/Z��{>�"\c��]m��>��Е��EK�GߋEe��'�"�6��z·X���i��t���g����dBw���S	��T �,i��^�Y���f{5Z(39����s"�Q�D%b��Z�m@�ũMr�j��x����>k�϶e(��������MB�A��(g�c���H1�,L�$����E'{���(��T&U��]^pOՄd�WU�\�u���ז�*�xK��9,��3���=鿩��s��9M��<I�X���'�ɤ�W� �fbi�TRΏ�A4�EhX�˅��>�4��~`7Wŝ�!OQ)N�U}3�H����L�zޣ�u��*/E=�T�T#of�qz0z��Z��Nmg�jk��?�m����$s�p��QT��]���4��P� �/���ⱀ��*8uL�_��N��^-G���+�ų���9��"��`^�%�D��~l�f �������Ԩ7�z�"��'�X��ں��-�~��>�>�|)��v�9��*Nɋ���b�i'
;:n�Ʀ=.�Y6�;�@Փ��3<�ᒻD}�v��=sF8��Dz|���TlE"�j���#|���wH�NiO)���5�1jPK�]�{����|��4y�ԗ�4B��vVU�pq��zPp?�����̅~�v�5�1*�Ϳ�;JP#9<�s��9Du�K��ŕ�?|�0 ���Yɯu����4̾�D�]�l=��;.q����� .�\vo(�y�7�^�y�����7F{̈��N����\O����	��7��	��ZJBuB��փWM%J�͛M<�y̢A(���72	��d��iچ8�k�|rm�?�w�i��j���Qj�t����u�6Ǌ�R�]I25���z,Z��X&�}��a`��3�~nS�)��^�zGے<�-ū�t�}u'V��X��4$N8{D��q�*Y��m���ryUi{�E�H*���R'L��-���I�o�;}�fX�j�m��`�e��y�k_*{�����ѫ�+�c�n&��Ɠ�$J9�$Sx�8�����OKIF./? �C�x.O!S��p��ժ�ˉiy%#�9M&@���/ˍi��&o�m��,��<
��&Z���\L0'��5@���3T��%�z�%f�ȯHB>Wo@@���?kD(���s�|:Tuђ��e����;�x�"��P���0�ِƍPHW߂�/P�Ĉ�����3D�T���\�:_gsH;ǻÀlTn6�yu�R�R2݌@�������E_���0]����)�Q˝�j*)RW�'�(�x�ja5�Չ�����]%P;�r��4oU�즧"���f�G*��={�e�)#�����H�M��ՙ	ݻR��m���|�/J�~,���K�F:T����a�C����@���Pk�D3�@ЇL��M����=�0��,.v��tXRǣ(z�7���n��6<u�)��Z5.� ����\Pe$ 0��DޘmD����u,��g$�r7�-��έC���ɍR�IE���߇��u��^O��.��?5��#b�N>�G�93`�*���:\�<5 R/��.q�3�ӟ9h{���҈�TS�K��Ɲ`R *�5�+7�la@�"	d84u~zQ��jv�q0�;/S!2`}=�yF�"�w��r�)=k�ŧ�㈫�JKh�E��O~���AE�����9�]�J8��l�۫�0�����V�>�w`�ϧ��G.
�%�Z\��cHN|��)䉈0��2�����
��D5E�Qb�P;Bw�~V�9Sm�k����\w��G�Fv�N�ӤEHK�3��,G�h����4��x������EhI� m@�
���_��Jsh�,��I��Lomk[?��*�����kw.����)vL��mk�`�6d�!2��^�:7i���?�2��/�4���-c��d�h�N�oMEy�,�p(���[����1I�����6,��XnY�N�K��n[)�|�n>;�,>��g\FeL�ޒ'�#2X�T�㢐FI����I��� u�ddjyS��e\� �t鉳g�/�;�8�^5��6x��ad�a��Ե�L�<���Y���̶ݜ��h�L��ŵ���0 �m߼�[ ��C�6x*ƅcW�����3mD���?h߻!5��\�!~� �C�jVWXͧ?���!%s��h�=��҂q˺��{n�S�3.T�5X������-����-�X�s�됩`f��_ΙM"��q��dM�ܒ�9�__pY�؎���0�YZi�D� ����a�91�4٬$��l��)�&�&&�<�o���g���1�e���X�
�$�1�vg��	!uR�u6��B�%�g_�'RƗ����*���F�׮�Y�V'>�ѹ	b� LA�����f��Qx��g�:������X0٤�]�)��B=��&�{�P���n��<�&Z)@f @4|C��s&�|]����'o�%�;5���y���o�:c���� l�����s��h���qx�s���R���.,~S����;3I�?��r0>خx��%�W!�rq� "p��	&p����7�b�q�n
� h7:E����8�f�~q��c�Y`K�!�w�� rҿ��j �4F��.Ms�i=�ٞ#���/%bB���(E����"f�T�����7��_0�RvĒ|oj��}$�[�M�:�5��^��A��0ˆ���w�6���TS_��S"�k&��.<�b��7.�
���3��q��3�zr��{�.�vJ/�u����1s��g�m�#6�N�C���`ؙM��=a�yp�.]9`�<u�r&1\ۂ���R��_ee�@��G��1^��V~�mg�k�'\�k+ 
����J��K�_8��8��;���w��x�B6N���A)<o��c��%2�/�fIhlМ:]
����xV�,��~�D�j��W���9�g����dnE\x�/l�y/��e��b>���@x��9�zFI�S�;�]�J�e�=O�ƨ��W��ߛ��2H��S�}=#`9�Jc�x�oíԴ�AFTol�p��x-!�- �B���h�Ԧ�;�la>p�aׇh��oLnaR`�S���v=�x�b��R;�Cw�V����DkZ��N�d��+5F��GZm�bġ"����E�Ia�1}��{P���v���|]�W��	��z�k��q*���3�C�Ux�#�ª�@ �	��V�����5H�����`}w��,NT·����	�]O
LbR���&Õ�@k\9���<�&��k@*>��>Z��rH�WK�w8~$������?�C�f�ɗ�+:�+	�	�.�2]!����"���O�����n5��j�S��{NSq5��&/%���{(o9Q[�9)сRSD-�{��o�����LAec�Ow�D|��q�'႟���˗>�)J۽�0O�?�TA!�?���J!��G
ߌ�Yw�@��s����mN"�z�nj�&��2��~�t��5"f����ƌS��J�C4O�ke$��R�f�>�����5�]�q[�Mm�\ċ`K�x����r1fi��DGf{M�pk���y��K�����.Qj
N���fV���P!��k		�ț�_����{p�������W1|�-4�,������c,'� �(R�'r��A[};�N#�|��$��)��d��kuxB)}Od� P�=8š�m;fã��7��ꑊ�-���Ϥ7_*F䉄�u*��G����#���p# ���a���k���nˀ�GTΪ���Ø6��G�[g�ÒL/m�ꗊ���oނ_���+ �"j���Z��
�V���W�L�bT���,q��8��έ ����a{af�\�fg���� T|@J�4����6��mJCru��ns��0Z��K� �F��F���lu.-"��A���!`�@*N�y�d�NC��% K���>�5%��y*��&�Q&��9�2Ͻ��=2�-�o|5��⌉�ch�&e�]��j/� 
.4�6�V�$/�� �
������Fr�Ј��ژx>�%y�k�j>ߨ�;�9-���,Ǻ����7Å�]v�X�56ύql����F�+o��-�v�K/�꼯��4·��������P�B�v�-6�Y֣��D�(��
2;nE�2�A|zb��-g�L���a�)"t��$o�`�Z��nmqh�|�5�HLj(Jx�do2�u�G�gRu �����lG��_z���{���F?
?���)��sq��<)�_-��V=�uJ��v��l����ߛ3!2���\�$�ʯ�sOq�#��9z���g%r�/pıL���ki�:D�+�Z�,�[�FS%�4��^A�%�>!zk_��SƊ��9a���c��l�q�<��f+-@��������YM5�27x��C�N��=�k�:3�1�؆q�6�������&��LR�ߎ Q�bP�3���@���t��/G��*H����s F����R����H�19���+E�����Uf��r��k`��l	'(��ԽY���GB���$�Kd��<*��B	��M�h�;'���1r@���7�����C�oo��d"�4��ezz���
�>x��'v�@>L�� ���U�-�eWF���-�-�znD����c�ӧQ�qD����;�4�֥{<�@
��X̬!��f�F�EW�A�n5�n�EĈ�y�����J�v_DԒV1t	�l����	�h����>�ɳ6G庀���Q3҈��'1PWpǨ@	>a����t�g���r����]5-\��[q��Eơ�.E��I�\έ�K����_DZA5ֆ%���uL�.m����;a�=�B��q��"�����'WDX`	�C�k���9�&��[6����@Ʃ�;P��Qf�Ǐ�R[kbg��';.d.*����ɇ�RA���/~;�79�"�I���,brYs���E����*o���BD�Ε!ZLp�vY���oNTw��w{~~چxW&���HoX� *.�����X�W5�#�k�RUIȖ�ha[�_u��}����Hq/t�]�ϞJY���L�y2�1�-@�|�GM�;��R5�m������˦��|{S�BB%���\��ea$�f�?B7+j�1ЊK���UW	̆��L�\]�Eݤ7���\�|:L�9\6)
��n��c��\{����*NXo�ω4�Vg@�`]?�= 3^��T���K�����Lܝ�<�7����OW��ަJ��օ4����l��g����Jxx+|�p��0��	7��YI�O=�NW�;b<�yB��l�~��d����m��3��9��̦	qd]�y���g��d7�<�w��IM:�y�*y�~Y_#�&������() ���nT�}XO�m��#龁��B'��>����RF��.i��c�|�Ӈ��q����i�~Z���]e�$;<��F�D��x��ӄ�O�J�	Eo&B�]�:�ez/�='����6L�83)��ň�0/�B��&|��k�ZD sU�v�c�9B�	9�]�>�8�����:�:�-BuEW�{a*?��*�yH{�&��M�]��s^�Zk��� �R) �x�-�h�^"��l�U�nG�#*"<ؑ���m�j��>p��Xi8����MXCɮID
h�y����#����&����j]�-�a�tv��"����/�z�Xr
����y�1;�+}ץ[� [5L �ϲb���>��8���o�f�3��0�8�7YV�a���"g	�f���� z�T]� A��yAU�E�Q.�����
�+��_�
3�L�0�B�2v�Q���Rȝ�$m�<a��2�u�a �v���S�q� .t�p(��){�C�``����Q�V�Ṕ7�\7�2�sEE�J�F4p�m�˖`��OM�����C���U��K���ܠ�Ç��np��������tG��=f�瀮$@��57��	�H�U��S�f0�	-�.9�_o��	�Ҙ�ם.gх�k��oM�8!o< ���^g���;~�����"9Ϲ�#�|^�s�<�w�-t&ks��$1gͳ�S���Zk�Ўn �2�;������>z}��$��y1�Կ��ٓ}oж�"^����
�	dȥ����~��(|�`�p�Fa[���ǁ��paP��R��S�ؒr ���������\^bd�S��x��YDTEۇ$��[�t�cn��X���ڤ�@��9	X����	�i����;�!�g)�(l���'��w�"���%�)JV˼��J8�R�	s��i�!狎6����	'�V7:��Ϯ=�'g���!�+`���.f�����0!K�/#C�ME֒��z�ZZк���,�_͙�vĄ=���2sՔ�J:��ݣ�/���T)~�k�V�I�09{������}\�Y����_��I�G0.��斝ל�Uq�a���8���`"i1K龞x�g'G����6�V& �Hhj"i�,�◚ɰ�C�90,.#zcċ��T�U6�����6�B�a&"�k�=ç����2��͋%Mߴ��9]�3�s�����hW�LizP=ɨ�a�A۬uR��-�7�������`ݚ;�qH�
 S�S�+��6dW�'���jq-o�fV*��6 f��z�񋟭2�;���t-�6�K�)~ʳ�"��_��L�Kږ�
_����p�@սq���t�m�&�	5�v�rh?�Dd�L�d�h�����'O�n�\�6g�+	�QD��:A�'k���1s<���9��ړ�
^Ѳ��pA.�������1 ���C���3M��0)��d�d��X�X�~�� ��t�]Bw�v���JG)��`˾	3DD�#�wOi��\���%��������"��'�.oM�>'޲�%r(`��B��TvB$�8&�k�h$�^<k/{�^�G�M_�
� A��6jE�rͧ�:Y�S���g�_h���9��c��\�~ִ�W���ۍ��EL~>Uab�[\��v�D��r�1)���&6�Y��qk�p�3�+�x�	ω�W�e��pߘ)�et�>N�����[lhR��%"��Ԃ+�wLcx,f<�g�£���*Ϝ_�8��P{��l���YU�n*� ��T��Qh�r0��^�����վ�1�<�U���d���B���z�w�_-�,5Y�O�l�VE��l�����Q0 ����ު�z��A�L��R�V[_uvKх\JNS�)V��ƶю�ކ���d���=&jqcP9�N�l�=���y���jb͟V~?%p`�\+�7��Ḃ�Z!�t���6؁!�{�W��0��^? �+���ߟ�<]I�����r(�_�'#���^�O��ч�L1��8Մ]�k�g}[�x��	��8&v��%�R�\L��!b�~��jg�&X�d��1�N���,n�P���B�6����A�[�5�r{��|�<��KѺ�:��Ů�0�R{&	��,���u1�ޜF��M�.�q�R�R7�X�F���gl%���R�ѣ���M�f�z��9*yo�k�aw=0��$T�<°�NaX���n?�Pe���Z���DҤ�:JE���]����-0�M��A���J�����A����eN�[쥂����M�d��,eS�`��z�ָ�V�O���**1y�HC��!h	l�v)Ano�>�g��*tkH �"TO�Gv�ߢ�[���������Z���ܚ����e�,�q^d���+TwH��{V[�RE*��#�x��5�! |k��2�V�x;V�����3�c
�F�e���ΆR�z>�3��0�`Y�`�]Y��ҒY���s[���/�r�5��\�~Y�{:]��P3�MgA)K��<����������`�&0��2a!PӅS��F��I�<=;\01��G��{�7'�E���"��C�E��ɒ�����sb�v3���	���Z�"_2�XQ��F�v��86/�3�ss�(4\�>���Ma�{G°������%�>C;�2|-��!
\�,1�X�\y��*�g�h�T���f�=���a#�I,)�y}}e��^iXҝN��z�Ukt��aHxn���ȧ���� ��v�S�mkNL�����D���L�-����4�Ɋ���z�F`V=��t��{2{^Ŷ����\����m��U��~�/Cp�,?��1���OӪ!����K0��&O�';����iXJ�������_��3/P]h�#�5����o��ðIa�j��$��D#`���='�T����2vL�zQ(Z�k��ȓ;���n����eF^K��Fi����/3F��"q���S:#�	��W�N������G�X�hp7��7�Z��pS�Й�|ʙo�y�V��6\�[<���_��Й�E.g�6pF��R$��HF��)�r���0�	tCҴ�$�cͪ{7nwaqq_����:pg��1E���u�ĸ\�-���묑�NΏ������du)�����f�]l�v)g/~���G�U��4@e|u��k�K���眲�t������O4!2�*�R5h��zjH���̦�oh��B�Ȫ[dI��ފ�y~�و5�1�OȶP�(���ܖ�Ŧ{Α�>һB��
��p�d[X�?���H8BP!ַ=L��'r:Tj����	
���":'�Cpn*�U���`�2��>7p���e�Af�`d4�LL�6�k�3"�Ja�� �I�~��5xN�� �>{b���������)�~���S�Q]�%��xn}�~!���A�)t2G���=�ʙ2`�͆�����˅w�h&�묞��A���c������7�$#���� oP:��І��P۟���	"���ٵ�V�Ӵ7� 9�ZZ�lDީoQR���/H��~�{l��u_cE��5�1�x��>XYlҍ" �+jvx��լ�b]H�Ȓ��v3����3�adxWܧJrD�|���].�qaоJj� d�]~u��~�*�yQ
�-"����ֻ8|u�N���GAԼ��g�G���Be��ʟx��b�ẳE�:#�w`������y���3������"�����R6���!f��Z���<%H|z-Y-�o�D�Nr��=�N�M��)�T�Ǽs�;���1��=Î�U@��o���}���P�%���}�ϯ�s$F-�'��ugACTx���a�O�j�&)!�&�_c�̾V~/�`�Ƀ�4�	�j����O�G��� �E������A�E��5��t�gT�P�U�E����C52Ԫ7Y�x�v�T�ʔ�x�ѩ.m3�hc���U�*���0� ��D��-Wh"��`=c�k�°����9�P�@P4��Eo~w�XK����%Wy���;T���+	z�c����Gߟ�׃ܦ�+�oA�g[5�\�4��s9l��٧B���$(��?B��W��/x �[ˉ a��;˘j�\t3����3�k�E<)R	���M�_�ݙb����O#��s�3�.��4�"tL(��_�K�[?�Õ-E����~�Gh�9c�bwjVF��F�sa*7�O�ZG�|	�!j`����Y�����O��ʎ�����)���N��|E���y�\q<"���n-vt����:N�J�.�����<��\{��͸l�o����Ee��x:{?��\j� ��(�J�j��BH�j�X�`��~Kd�H�&�؛52�:�'W����F�4�?��JGe��W<EFM}�<�[�^i�t�$�ոf�������᜵�egb�!c�ߎ���LP�D�b:+SR�Z٥�<�ĔP�柞"��pne���ڝ$�:� X��3_I�>sOC�n��Ȳ�I�<	/�Pwä�^:��D.�����?Z��\y��ua��r����y�2���IZ���G?<��B�!x*��V�@y߿#ir�Y��K����.x�FEWl=���x$���[������z�4s\�)(��T
������*Ӭbf`an�7�Օl�p` �u�zU���͋�%�`S2 ��c[�ᔛkL�3j�W����hm�pS�M��_U�$ ���6��|��N?����01cޖ�Ɗ�[�S��<r�CU�qA{���:����w&\_�����YE�����]�G�pW%zWW�G�[s"p�UŰqC��y-�%h��v_��'Lz�����C鰼�,c��S��n ���M\��q^,t^nَ���t�K2 ���9�@#�/)&����f�>
r��`�1[�o��r-��֝D���E�A�ru ���j~�`���w�\G�z���f��9�:�"�q��1��5��ɈZ9��>#�	��_�V���r���� ��׮?�c}���*����z�"0/v��b�U+�K�/^��Zھ�S��O�Ġ�vt�π��^�A�|^Z�Lp?�{�4 ^l�Sܤ�������w���'Z2�I��F!l[_�L�%@q���Ŵ^�}�`�G~��Ja�8%��{�е�Q��i`��G$����kh(hEF&�O�oɌ�E�V�Eɡ�#�IK�`gO�Ll��k��,�����jf:h*���ŗ��4���N �^6uiȳ����O�$kD��+�T�2Œbf�vJ����8��R;�4)�Tmƀ��::�,l��ID n:_�.��5�MЯ�/5���%;�[k{���8x�B2�zmfD�>�!����"X����b�a#�P��ҹd"8q��Am��T"ҫN?�	�"�N�b��|=����v�{Z�N&��S�?�'�j`\OXtU�7q�����Q*�RN�`0��x"����i�~�L�^�73��m����W���UAh�7#N(�yj���n>������ٚ JP���4�(������"�c�����~���	{ٶuH��:��G�Qu�p�N��X�#�l8&���<���̃�{	��&�B�b����'�9�n��e���ҰI0�w�A��.*)$�>
�qXW/���]+��T6v�ٵW/ �� ô�ӸC����.����^������1$,�0V��O��T�BZP���gW���`;�cn�73o!���������/���0+{�D��՚cM������Q�va����'f�+��K���:҂MZx|��|��蝐�Nsڍ(`3,����"���z�%:��dN��D�"_����[��P�^!�F}�b�s��]AL%�1Ə���ke�ۤ7>�S{�;@EW9��{��ᤋ9A���ǋ�
�5��,�6�Ƿ?i�c�
�����!���������T���'_|ea��r�� ro��y�����P]32�X���rm
}�ARUƇ"�P{qw)IȻ�"�Κ�'��7�W�1��w�W�IЌ�*�`�������&���j�iua���IF�,,Q>�zz��-4o��R��Ӟ۽W�5���u���S�ɩ�76�kk�z��:��i[���N|�z��8��p#;Q���R��j�Y<2��F�{�'wJ���3�M�Lw�iOj�_���=Yd��w�O�8W��7q���gM�<H);2�	{R�l�iS�2�
��q�f����I9�i�lP�a,�vAK1�%̜>��IS�R�����	�MA�G��ٲ1yp)Zx@u�*]��_�+-�<-�o7�/-�aMۏ��Io��������� +��Ā��{�˟oSS:�`�N[��Ң��ւ[��:M��N����e!nM����Gfi��o�*|]�;�zi�'�zH�қ������Ԝ�v�S�Q
��o<���˕�P�����URH����^���7��xSB�ti�U��'鏫�b��n���*w��ZA����N�����UlL�U,p��=��$39*��u�{��2��Q[��d�
�Jt�s�b��F-�BA]�]+�����u.[Nc��"��~��
�rA�h#����$a.�A�)k�����\�z�ߺl�y� ������1.B�F�>�v@�����u�ټ�jG�\��� �AD��rd� ?7Q+h
&.f��E�@�X�>����f��Oڔ�v(*)qV���Kظ�J+V�M�[�������{���L���jO-�R���o��}�U�I�(*�:e=̼�1�����_4"��ŧ>����!�(�F��[�AEH�eL�<V�iD��T7}rs�(Rc�첹�٪� ��'��eӫ��-g�ܿ[l]|���6
������NOz��nL|�����l˓8 }���c���+���������j����T=��t�v��R�*��f��eMw�)e�0��\�O�j�����d,]=�!&�ڙ�7�qp	7I�d#�/��B��7�W����+�Sƕ'{��CR�3��<|��!�N�N�oK�|���ގ(�4_�C[C粝ъ�ɪ� u�ܔ	u�r���PhD����Gi�4�����bd{u�2�m�#i�q	��F\�Kv�H-`�;JgH*vL�{7r�u\(��E��������(C�uLe��{�k�Y�v?��J
�q{H�M�A%��d��#;?�H0�ǈ�\�Y�
���W�,vQoف
M��<�{{i����
�?gW�e�[y9$���A�.5�M�'���-Ưtzv���*��VR:�,��۴T��6S�f\!6Ha����E#�C�YaL��넑-�i��	�]q�����|�,��<��2���)&ʍ�+�K;���Xy1�C��H��X��$y�=�X|�eئ2g�]Q�p�1�����W��'������ 쫑o�:�ek��s�&eE8[p}��f5k/��2�g�iI�Z1�M4p\�E�|t�%н�#���g�TZ/�SN/�7�O��(��Ć��H	dޅ��G�)D}�e�N'�W%}uőɛ
��YKύ����=L��^58��kD��*�Q����+׈N��M�4�8�ú�%���"H��P>���Q�^Z��=�ۆ����	b:��彪|�Ј*ڲW,�;	�����*���7@-��c.h�����y�1�<C���휑�a��Ƨ�B��H�f>Lů�0�	6��Oq��L	����Nad��>�o�n-�]�*b	�h?�R��j�:8~�������A>�:5�A��U)(�I��+��{� � Yv>ߦ����1}����R���i�����qt�M/*~�NEl�:���P|�8�k�aNK�H��)I����xZ�(yf������+�D<�0Wk`�@ٸ~T@�T�Ǘ��;]̜���{��2;2��.�ռ�q9D�À"�XU�3�$�`[�#�u�c�t6���m��DU�]'��f�1���k�[�LI���#Q��Ι�J�F)%� �G^�n|gccw�j��0qV���E�,�{+�IߪPR4 ;��_�Ic@�V;Y��L������r͉A��$Q�	M��+a�����mk�"�Ld�fb��5��|iy�{�@h�<4
�J5��bȡz z!�?)9VMv����c�+��9ԯ��b��gd����Z"�n`�;9f�x8 )o �����7"�tP����E�R_Ϡ�R�q#��J�8��A3ӛ�${�zo�DƣOtU>$�����PmOz��l72y����@�_I}��\�VA��Z��	�s����+�G:��Gg�v�dv
x��V�ޒ2�漦���e� j])��3]���Me�!�]�@�ӧQAb�����M����^�Ȅ���&b��� �Lbpk.�R(���9�"T�,�%�d��k���G���R��]ǽ�;��;�/ ��\A����+iv��	Q�\�2��^��7�T�AS�f~z�0���Sҽb�z�C�佼.%��M`�b���4,��K��
�����C�L��3c�3v�9J�A٘��d9ȡ���=y7�=��&-��R����s^�󕳘Xڻ��$P¤S݌~�Ý #�pQ�[?�Fk@y�<��F8����?�vɄ�����?�βh;��v�:�{xl�����m�j�]���\컑��O�������j����A����
��ƀff�@U�7��D��z��H�(9|�V��-%ϭx�K[���g�|��.stDY��p�Y�RN���Bx���:c&W�/��;K��s�Zw`����@�^�=�ٙ��)�~hX ��m|%4���*x�d�~}�q�X	ߦ���7��+��7�Qxu�s�Ci���EY�sֵ�AA�E��=~B��������^����YP��y�Ǧ.{��A�qvfs�I]! ���"�ߟ�'���M��m�v�g��V�yx :�~|_G�5Ř�Y%h��mZ���h8t0Vv@�ib��/$ދ;XM#�)eQ_;���"R�%t�����Z4Ó���66Tp��x��X ;�u�q_�����#�7�0ml��.&
�� $�?��Ų��B�	Y���^�Eq�{*E����K���ȇ p�����W�i�#��G��ʇ]T�E|��F5�z?�>��<3���c��m8큫~������L�������[���4YG�k�X��E�qz�G�C���z~�I+�v��Ţe���w�t���[��ʹ9��iU�V?L*ۭ��&�}`�QeB�8H	�yO-Z��B��ҩ)�:�V��L��`Gk�@�wJeo�~c_��M�3�i)g�c C~���y��Ұ�JBuk����w�u]�ӓ�F����r�4�ft�|�#ۢ����T6W��R֨ ($ N�7�k*]WC���	�	f�I��uelB�Z�1�Jڅ�'��נp�R8��N��v�� E�����>��z!�u��i5��N��L.�Gr���������ڷ�
�t*?wB8�t�H-�h�a��&��yڨ��H������%�)�Pf�3 <�Ս��^Iԕ���?ݘ���9��s�V���P;Wc�A�lpb�H����������*ϰ{ڃIy>���[z;����u[p3��k�u�"Ʊ�H���&���n�ˇ���\Um-)��;V��.m�+��k��\���[G�ں�/�K��6�=Ρ�� �e)U���1PJ��>;Ex�7�Ժ�M[cʫP�5.�L�k\���3a�Z����c6p.�{	��]�ԏ\q��tfG�Wdww�T�Z2�AE���P��������hE��^m��1]�S���X���(0|_�o;�6?YVn!vRҤ߱��{�TɏF_?�����^?���Evp����u��:�XjK�����%]�T2W-�c���r�ڟ��ܘE[l2��� E��KM�w�Mwf�{��%���%�K���d�F��G����K�ByR��*ɪUs����+jP�Ó��8���,�-w��X��$G�j���B'�����"��w��#�yg;���R��B�Bt���a3V 	�@%�`9:�#��bkri��{۹YE鏰whm�k�ʒ��6I?���^��AQ��~*D�F���M��R�bI� 6I���P���rn�f��1���c���zM)K쪺���F>\�D�Rj}*��A��n5�@�C
L|� ��c̋��U�v�A����5*���v��f\��*=�'��d�6�B �a�u�`4Q���Un~A�{;���؂���n{J��V*n���
�r�<O�|qM�&�H��c��mo��v��zz.c�k�"MW���Z�%��PY�,�`゠JF�>q>v]pӾ^�s����Z��o2�:	�^[^�M]�V��������J�s����T��)���A|:B�%�^��z�N犀�p[����N��U�m��.挞��J34.)�W�5e�;�%��sb��Wp�k\�Gj��\8���Q<����T�?+�q5�� �Hm=eQ7d�d�:>�Υ�o�ͣ@��\2ۥv��َ�x����XLK�5C�ΫE�H��	���r���p~�3�,6�Ȫ^vb�g��[r~X�n�}W��\+^��5�%:XUS��~8�qq	)=Z�j���^��W\	���
Vw�7;r�л��#�#��	��j�s�/����Z������>ِz�b��Lp������"����������|�71"��NG"�@�AG!�\CkI|�P�/^�Q-��qF�zȄ!�*&.N�2��>�x1�mc�&��@L��#u�UrE��޶�ӑC!�|P
�%z�۲��u<ё���}��JMnHC���"+(����$R�;U_��;ʨ�
�ѽ�\��N� ���
�grYy�z��/���}�	���k@�8(�y��S�[\�a%1�3�����GL�Q���L_K/�QJ*Q��b�a�n���m�c�X*���h�t��Ǯ�o����^Hd�El���:��X�S�uaހ�`Mڊ�0h&yD��S-�7��j����ߜh�E�a�q7@��\��|��}��ü{������ ƪ����jeI`9��<ѿ5	�}�|��k�e�� �5��lF�s��3�w�YK/�����<$.�d�ݤ�@�u�ygU���l,��\.�]�㕺_�pH?h^J�����B���E�RsƻϽ��\eQ�a����{-\g�̡����D��hɣ�qR�\櫞��C�,d]��ũ-l�^>��)J�GwZ7�'@ƻ�?��i���s6A���E_5�S���>�oD������$�g�&zDta�b`ϑf1m�^+�k�c�����%~^��37H���<��Z������6Ү�ǜ�S��;�]	��R�D*�B����H��ُr��I6Q#<�8H��HJs�w�Whv�����ĝ��\���1� ]a��d|�e���rT�/=�0�	٠9>��[;譒�b��ranpB�zM [�Y.�?�	�qI8�+�'lɆ�f����ˡ+�k�m/ك�@��69�v����^e��A8$VJ�����5�q#�?>���6�-6J�A\?F��邻G�t��ؐ0�o��d�C�̵u�#mlt��A��vq�F=���W��G'o9Pi���C ��~2+q�]��A �����-�]��i��]zN�4��^͑�7�0��L3`�C��JKQ��4�t ������ �(�-8��U���H����|G� Iܡx�jdDK#���梂9D�Ƴ���V�D5��^����c��(��W�>���
f�ߦq<$<�ۣxI8	C�z��T���,��]ud~A���a^3ER��H�m^r��[��!�c�\�h�r��2�4�
�Qi�}:���U�u.i��� ���.KN��i�����H�>�n�2��l:.랡�_N,�[��,�-Au�M�\@��`�7.'��s�[�d�Lx�+��ʰ�K�9B~�E��Wu��¸%@x�?�����9_+��&���پ�+���ct�(x�à��+�adIJ߲�ڂ4��hX�F.��'�����+Q٢���7���Fz>�o�cn��z��{v��m'��w^�Z�Ģ<T�(�[����
��ۭP�W��B-����`��J��!��;���]�K�(�\���L�ZJ���� �j�a��1�7�߈iM�4�-��O&�"^i���1`.D�V�k���D�-U�.�+^��X��;�OO��a�?HEт�ʝ���T��a�j����J�ߟ:��g��%�31�
� �����D#����k Y��"nl.Ɇ]������)m�<;V���3��-�W{1] �_�Loh����ӑ�p��r+�U��7�:�g���Jo�����5�%8��ή�/��rڰ�j�GC��r������DD� �Ŷ�xTF����C���@̕V��E�X[]RO�t�Q�;����<S�CD(�w�d>�H�x꼾x"0k��/�e�m�-w�g��uu�r����|��s�5����@��}�"\��C�� �C�?�a��c����v"�ؿ]�fX.�ލ�#�{�� 6 ����ӐC�j�褢(K1�B����Z]z����ӣ��ܻA����|��}�J��k1H���W�����o='�6#����v�V^g����"G���{����S��@F^9�1լ����'�~5]�c�;B����薛�<��>�z�x�c�{\Gc�;i�z�F_���w�L��f;L��8:^����	]A�V���e��Q����t���hِ2�F���]"Ѯ�j�<N�_����ٜ�n4:;S��9��Yd���������[���������܋/�\8K$m�}U����~*z��E��ɲ o�Z�1����s+ Jz��}�StL��hu���y���#y�:H9�JP5?�����x���sng�X��sOșkw�e�gXĝ�Xߜ ��̷�h'>��!i5a���74��m|�}����\Y+o���
�-�9C̄�y��I='��T�E~E�
	%��SB��<Y�~�e�!�w�C�2%vhm�����!�0 I}���dt�?�獫��� ����������O�"�����M�����%E�Jìf����ѷO���PҨ7�&�����[�&�rθz�Z\^6�����ᴹX^O�G�4���^kJS�	"���4!G�b�sՁ��p�Ӟ$�\Le��P�����+b8!��.rN������3��Үڀ�eL�������ۗ'�n�Q���ȩ?8)���ߴ�A�o�v~�D��L�;����Ƹ���L#�&�,�.�\�Y3���F�x+O��!X^������Z�E̚�|���y��W��9y	I ��H����.�m�f�����S�嫪�ɉ�2�f?j�>�|�0{5 r�
AaJ||� ���Jm�X��L�o�ɸLΤ����@r�ox�n���Z��#��-OF�ӆ��m�/��ʉ���X�ǔ�u����C��K�L����7�l#�TB��o��x/�VU�3U��������<����02���m*�7�'e5�R�sA�cw^�����"�~m
�)����|4hS�-����;�.8Ca�T#��oF$�W3���q��e�Acd:+�� ���ٶ����A����f�ks%Jgh��o?�g��ȆЭ�#7�����4R`"Z��TG_� ֍��|��z#�9���9�Z�B�Yh@��6�'ZAܺV�=�_��X��E!iP�o�$Q�\"��1�:����`B���u������,��֑�ZϺp�s�Bn��f(�D>U;Ҁ���/�5�[l��&`���?�����8�������aw.�͉�S�TJ|3�qg^��E�wZ�Eͱ��,�Q¡+a3	fsK��/Ւ��8��C�=�i=��S"�,任������=<��Y�R�:����c9m��l�4A��?*߂��ذ��7�kSBkkH�L�:�����ن5�CEb��ө��χ�i;�{���T����'�s�%���adǦ�e�ťEX�Z*Y�6��5G�;)��c��S�Q�=.�"%?c��XF����������q��������4E�#<�����fQw2̕��|�ˑ#�yy���&����MG�K֮�����k7���$Ò�g������xqVy�*������6�I�mU�P�u�$F{�%�Ī��O���q�[��y<z�r�!�#�Kљ�������4
�.�qX��bڼ�	�F�ywĶv�_��Y���5���Kh���'q�v�G5g=hU�lG�@s�����c--��ĆP	F͏D�#k:Nͱ���}*dk���_�9�KȐ�d��B!�o��$����`*sp�Z�U4���e�s�e��j���4Lz^����!�v������徬xP].�s���<�s���kII�OU<ّ�r�M���e�� @Δ��zz��z��7��u+娔~� ��x[`$�'j���t{'3f�hr�n��M���S�K�朁���.�.�^���Q�9σ�hN�훔��U�+�!%��ٵ�>~0Ts�r��� L��v�P@\ut����FN=P3֬�}�����@��'�M���$Ў��XUݿ͛��V�ӻ�u��t�����z�m/���\#��҈�8@����"��<<��V�R��ǖ�*��N:�>n8�ʼ�ÍF����<�mB-ܒ��Л�4b����o.qϺP�%3�.?l&�~\����=��W�wv�艹�zy�:7ݪػԯ�f��I}�/l:Q7{�T��w���s.]YZ���ww^��EW���Kg6~�Km��BR'�<��'$*�k�!&`:�&D���xC`H}��ȭWT��욮T������䔑d(�;R�nBz���6] �;x�+;hI����V�
�[d��/-{b�й�߿y���M`�S'`�O�i���h@0G�e�H�̔;^g�p�KT�Qk۞?+�V������Q�Zv��U�j��/ZV����Gv�XxoH�8�_�^���j'���L��\�E:j�Gx~ϒ��ޗ��9�蘵��U[$oW����G��Ν���rNvelKMW?�l6_-4�?�\���?ߝ��x;�;)����z'�Lvھ��QKo@��;H�}��@������'��Z��Z<���F��X��,�%��{Ը�p��r{Ơ����"#@���K�~�U�όI2I��_���J=��*X%��~e/��,�W W���Ҥ��]{$��	.�/K0E�ӗT�{S4��n��@��*����m�� �k.K��c����'$4�u.{Ȟ'LO�X��;^b��g�ěDu����у��B/\�v%����Iբs�q�
)�Py���~�827��[��������/���<ݳ(������h��͹30��S�K9b�����Shm����ʚ�3�W�@���k��f�0F���zA��mjؽ�A&u*@�����N��ݓ�"������P�-��M���������0��1���h@��QvCZ��
���k��7��W��T��5%L"�(�Y�p*R��p��E�q�z�͸����3�����J3,��kF؝�@�����[}'y��=4��E7�
o��g�q7���A9z��/�wDD�{\�?��R��!%�օ]Uf�_ņ�gηO<�p�'ʪ�?rߥM /�yX�~n�۽�A��lM{��@����d+@q��}>�ht>�!��=��脂(�LT��}v�/����w�:,X跿��Á��j�aCB���n s]i��R,�#b��v!�uc�B�Q�wf�1��ep����r���p��9\�Wr��̵��	�M��L�]X�
޲�誘�\�#�z��*2��~E�����mm�
Z�@��z`��T'��}@��P1Y��i�����JQkw\i�7*�_\�����je�T��G %6w���ʣK���LRK�B�\�n�>z���@��"��(�n��v[��R����A�>�:�K����cD����L���8GF,��5�^SSHF���6���r�B���}��A"]�2JSW�8e����?��_�����+skn@���i�����������kI�?��|t�S'���T�;9�JŃ�<dI~vhd!���!�%q���T{�;S�Bk��y��G_���ܴ��6�v��
�����TL�bu�/~>���3�>Ll��[�g��^�`�(�֑����hL�޲�O�ݒ�G�0rmY�?|O��	S�'�[��s�k����uVd����E90��M���b�-)w�R�uB�NZfQdj݈[@��բ���$/-�P��ؠƕAbXe)�4�R�4	{��7���nE�"���8 �a������*i��
0˿�[R}�AEc�#�dˤ��.�R{BA���s�����ɟ�x���y�ExO1F��7��f����l�u��k�l�wU���b�Zno_I��m��M�۾����)�O�#�8�ۼ1Ώ�E�ׂ���1˞�޵�!бn \����i�D[1jB�н�+M�wL �@�S��e��,kL�������U�,��p(�:�3�����F���ܯé���cm
�-�?�����44؃��V�F�(U9Э�:.8��y�'�Ѻ.�v75j���}{?"�H<��퍨dw� T��h6m�����=�>@�J~O��5�vC�(M*�d��o-:>͌���e~Hx��$�к'�� .k�s��E�%�#�n1Heۺ��}|��=�\{	���"2_b���%Q��Iar��G�]NI�olm��&�|��|��?���U�j����="��^�v|R�v	p��Ku�~mBe���FXA���O!7�� $/c��i��޴�D����*��<�7Xx��lC��=���y�b/�c�i�_��H��X�C^'�v��L�5!DZ��Ł�B�^��<h�"���o}��ŗz�ל���K9N��S]6�z�W�櫌��P�$�bz�"�Yxf?�f���+��e�uXl��A�R�%��"�mΘ��= �;��	7z�_ᡡ��#��H��˟m��+T��i����ࡗ���əT����M����or�A��?�Z���/�D����`�H�a�x���",�\��^09l�>!Tp�p��`��#֬����fT�����^16�\+A(cYA�gɿ�｝�';�mVJ`��=X��D��^}���?����( ��$�|�޳�	0=�EY�y�$�g�{4������6`JB'R�7dŲ,�������։w�|���OKO�c�7�H����T���3Kr݉�cwl4��my�?
� 3=��+��$�x�X�)�}N�X��|�5j�k��?���X�2~�hK�ꄥۄA���y�NhY�.�K�	�A���������w���ea��7d�D&���׳c`Ǩ���BS	�)�*`I�2�]`5�� 9{�{kۆ�ܡm#��]A�Ai���tz.=2H|��f$xx WrKS��s��+q�)���lp�.A�}��Aس��e���F>�3������ `y^p�l�PP	��υ��$7������u/��<���2걚����tpÍ�;�S����[h<�e�Cl���Ց�#����CC�㠞��.�'���A�P����Y�O
�t��{sG�^y�C�����,Z�&쵾���'�u�����πRYeX�%H�Be���΄�K��9	��=�*� Y��%l�ejx�e�����G�RI�$��]hv�u�/o�4hB��Yzk�.�u�n`'��T\�i?
8 K�X���Y(�먦�?o]o��CK��*��sP9T�­:���E�hH�P��{F�歔���6��R�������f���ba������%���dŌB��\�zC;��&�r��0SY��'v0S�/()����ʌ*���*i��ꦆ��O�ϊ嬟��\�J^�!0����U*z]�.Pߣy�BRf�+����Z�?�n]����X�z>��S����M~w9s�=�5;�J���G���J�瓵����Z4A�H{���ē��]��H�6��Û���#����v���ԇ�#,�*Iw<KPf(�3�X6~W��r@����"s���^#н������4c8����o#�����4�
���o��Q�SZ��pI���=-WO�J��8����k[�j��' /)�����R�ٞ�p;vx8��!�gmld�E���tYO"��+�����_��a?������͟{ے���Z�t^����%�C���hNه��6��{��'ˢ��Y�M�	�ʮ�`O��;��"r�o�ڌ�a���ruՕL䂉İ]��=�~9;0"̜=�e��{;o���s����<5qn{�'S��s{*������fj�>�w�/�gq��*N�M�i�zORV�J]��3�C�����kߣ8�)��ɓQ�%]ݫ���|G6_�K��S(�	ٝ�u5���x��g�;އc��e^O���2��_jHn��,4����Ӏ*��Դ��Wg�+
��`J��,:���;���v��i�"F�#�B��ܞĜ�tC� �*Lߪ�ݗ+��F��M*b���4J�����9J8�E��n�C�'KF)�
0�7t�"c�>�'�,�AZ��
�T���]ݖc���'~�m}Sܾ^6���Q.a��$'�F��.�^�g�ZH�E��F�[~�Q_���U�.��vr�]3I���Ȗ�d?���ӝ���?��C4�0��KL�����e(��1�eG���R��r躷s��'���\㲙M�H����CN*�A��C��@����v�bd춐�9#t)
R>?f%$�WMU����� ���ͪvQƉ��EV��3�x�sG�(�r��a�ѳF+=��(#��Y��`��r��\_#����3J��	v$�z5^1r9�m�*�h�q����s�_��f9�VϿw|�!��\#�H�	�:�4ׄ-JJv��ޕs)��~�}by�Uc��+���6��:�֩4�ϣ,��e<��EA���)~�,�\F:��2���ʠ"0Ȥ��=L��yO��b�c�F^�;�O�ޑɿ�@b�����~���WDl���� T��/mP�cGl��	 ���>&�@q!)G#��ֹÜ�݆O�&Bƺ�{�sv �[�t�b/���Pe��!��F�է�=�{ʜ��*d�%���صu�Y'E��T<�s�_���G��UQ�o�3��lV˚^�:��i���5$qS��D��;p���9F�k�Fc_|h��Qk�K�O�|��L���n-n��4��������5jq���[��~ƺz1��<�ʩ�zG���Z��l���NB~Ɓ���9C���i�ܱQ�G�6���̈́r�bUR>���=���g��};)�Tn6Y�Ⱦ~ki5�Gy�5�����"=��qU|���'�8��R`G�X@Y�[����\w#��8��R�Z�f�!�ϥ�m^��,!��a1�rc�90љ{������SΣWa���?��f=PT��2&���3�Ӗ{��}�$&��tL�*z����RZ=�a�������*)=��\�+�'�9ܫ�\Pjc�g1�ក�St�Yw�L�P���ο)��m��ى��Y@X�Ǫӽ>�<�S7�Zs^�#ʬ�b�Cy�4�%��ك�1`r�����oL��"d�=�('����sщ�����d�V4[��;�<%�7���	R�������7����%�k�l	"�*���49w�c.2�7�)ATZ�"U�ķ��6��|ߺUT��$笀@��#��&���Z�[7�E�#�,Qdv��]�ϸ�j�e��R�,���HY6y�7cg�j��onR�D��PA �c/N_&�^U�iY$M�A"��W��mgR���_7��'�v�ꢐJ+/zo41���v���;{t�����8֪&�J�5��g/�2��M�F;���3�Fڻ��Wr#~W�0�q�-g�M�/�	�ɯt�0��Å�Ûl�ٮo��ʸ@P�(�9��y�%K10A�'�Y�Ip�]����)�d?�e����C���QK ��?�H[Λ�����5�����Or����w�F�l�||h>d�J��ٌ��˿!?q
�Z9W7�F�9m�5~2i	��᦭��R���O�n���M���O��H���-}�Z����|�[��^>R���
V`���|��~<uK���$m �f��D58,l��$J�X��GlSow`g��sM��"�_�q&��R�|}ƻ�{��ij)�ۖ�+#�Н��O�"J�k~e," w4�*c�L��J[�9d�:���M�z��G'��r���͘є֜%iU�>�h�&���:!���t�|CF��:L,���C�&#S�����=K��<	O��#���a"�a�h��5�`%�����|2�?��4�����4�����5�=9o�H���}k�f^]9�;�z�X-5�-���7(U �dc�x+��0��in�p:��(o{��2~��Z�˂�ޘ���;�ʘd�d�3^�V 4FM߼��T���r�\j��^5o���y{%JX��V�=�vj
P�w9\��6��_�m2±��@��e�%�����K夼�:�)}.�8�"��9���N�"0�2�n���/�N֦��lEN���f=�3$�#R�A�=�����j�p�ÂL����]�݈%�Jcʾ���g~�M�~i�t�|�쐎ESh>�q�v����Вg�������	�Y�yX�%;����{�=ڵ�.��#�JP���-_-Ckew8�5-�,]����G�j�M�.r�>T��*�B���!m�d��c�x
̰w�!=�8�M���Mx��Q��Ȳ7��D<�I��ӛ%���\xR�ֈ�!���pu]��jH��a��C��ߎK��ٸ��%M�+D�K�����Lc��`H��:B�0����s�� ��a��(;*���!Dtp���8�xK�-D�: ��� R���I��
����\�����9UV
O6 ��+��3t����|��Q6<v "��9Mn�Ɯl˝OR�&� J�����w�.����i�T3~�{n*^�;�6��gϪ��_�<��a����,���`�ߐ���G<FP<ֵ�d�J�v����G5�yk�� �\i�՜rf'��
x�l*,��5�ң�چ8ucz��W�W Ÿ=��J��\>�����*m����k*��h�m,X��?��#�!Edi�K��K�J�L{yJ��ރ��&1m����`�öɵQ,E'�R Gq��:<V�d|��!7�J�΂�-%$��(�^����\2rzPr4<��ͳ��{�����>g�S��}(����@ak�7���%�4Ћ����썐+��?G>��0�\&�fn}#3��M��Y��,��N�������X.�;��㽐.�<b=S�<Ɠ���"�:�ob=��y����	�%f����|g'y�����O�ݪ�M�]���Q�pB��U\s��c��x����$���ƺ��y�n	{�rT9�jc X#�5�g,�|��A`I��'L;�J��~DyZU\���
|�@`?��Un^ɝ�Qp5��^���x	H,��U�9:�
�<�
��'��E4;�&`븊�1d�;e|W�<�|��].�9-�_��I��B�����<�u��h擸V����6(�����u��HT�Z>�z�K������(�R�˛Z-��w�	 �v�9� �Rr��i&�>�6�*�/$��{�׼2�MB����p�����-���b8k�-�AK�B�WX|f���>曧�������5e���c�����Z������L*��T=�M�LruzP�������ĕ<I��CQ,q��0�ҏ��&Z���v�

~1;�B�->���{\d���@'���j��6� *�q
z�����R8�brm�B��{Le/���A����u=*���d!�,�/`Y_ �[�ۧH&9���)	��oY��fy�gZ�ѝ=��u)L��)��gu�
���A�alZ��ԏ�{c���s*@�3q�r���5����?�j0����r�����_��[���yR���o���s2^��@)�:���
?��X�|�����������
{lϸ�,�νEe?�|�axk�٩b���@y��÷�� �$�#Ee�04C��g����N�M�|E���H����J�T�[.�\�����u�S`�>�f=��t<��q������F��Ő͵�Ƈ��L�]��B�j��{����#���j>�+&�$�o�(�]Q��(ɸ�H�vX>�-]��D�}]��G�2S��V�G��>h�ǩ������*<�bN�? �����W!����Y'�0�H�D���Rn�cS�J�Ka��A�.J��E'�p2���濑m2�s+����
�#�� �37�{?�Gg�=m2����r�֧�����sVc�Y�Vա��"B%�����Ӥ���5?��J,��x�����R�P�1@�(H��d�D��3�y�|P�|���S�.+�y�����:ڝf2E��5G�� �1�X��'�L�f�-��<���S�F����7��W;}o����u��C��>q��Y1#��y��� jX!f��0e�Dwu��,�+<Vӝ����նC@��:&l+����WJk+��t�W�c�'�Z���fo��f.L��$$�P\��,���`�;���b�>भ%]-cy�v�VqTc�?�s#���S�2G�B\^��<�nމ��xZo jB�@�w�$q�`�v{@e�+�b(z��Pw��ߦA���-p\�&'�?@Ǟ��mgf��}�ҡ�����r�5C����b!����ؤ�V;��T�?����6��[�.QW=V���7��c�H�*�������@On�E/�|�\�9p3��u�v��=�1>���������M�
���-V;�;/��GEt#�[�"`��@�M���s������b�~m��uXpIOҵ�Ѓ���(�t.\	��_	N$��7h���fh����=lc|=�f��K��^�<1�d��N�-���K��ntT(� �tf�����B�_p�6��y�o�|�6�`*�;D��DOo���4��-s��w������>`�}*��l�)�����c�2N	�H����q�.��Z�-93�Z����b*��;��h
��|�S���;ω�_���MS�+&=�5Q0���e����
c?	�\`�%��$PS+oA���ҏ,L1���D�3�#\�^�D�	��T�E>M��x����%��f�k�0°�6X�bW�)t���6�=�K�d˖ޙ��\��,��� =4���Yyh�?� 2���AƊ�x�OL]N����1�j���P�h�J��7DX�S�ߣ��&��y� D�#:��k���6�0)��DOF�X�`����*G�#)$��	`��Q��'������r
>��ұ�?�^&X��K�(\.o��e<�f?���x�\�m����!���������!R�sC�~.af5GV"L�����I����T1(���q��=��ud��G�����
��f̍U��p (U�We!M	��D��f5�?��ź�ʡ1 cĸ�ڏ#�e�`g��
�C%qY�s'�^i*�0CG�#\].���Բ~}�kX�a_����L���-!�f�D��9���7B�P�sR��I�Qx���H�A(m���3f(�;��lI���+��|LΏ���hϲ#'��AZO����o(��9!�0���S��b���?�D�	�xC�@i3�OY���,�Qdh���k:<��u��t�bQ��c���hX��yF~��ja#UI_##��D�v -�L���$�Y�5|�P>,�f=q�3z�����w����L�.�T1�(຃�V����ca�<�CE���8=Q�;}� ��*�`N|~��	G���:@os����D@]��stF��ӻ�%[lj6�ǖ�'��2�Ёb�t���*��]�t�L���c݄�@���G� �=y��������)o������:2��i�渔��K���0����X���5��(����=�Z�'�>���=R9G0��i�o�����Ѯ}��<�k�%Gۡgv�n�\�W_K5P�`;�1P�����9r[Y��\Vz�:��Yn��)E��(��@�!N��;��L ���h��;_�`bM���~�>rn����RQ���rVh�P�`��<�Q.�ad��n!Lo�5����!T�
���K.&>��B޼s�ټf�V�h
E��k��¸��4p��ŵ��d>M,|��@����B���9ܯoTqDT^m<W��AY`�.���i�8>sz�Y�9�M�@�	��)I7���4��[d�#FNF����w$�+D���8KS���`��v��h�]��9�s�v����`��X?l�Te3`���3{&�m(X�ia<�"qkq����Ʈ&�)9���O6�O�΍���v���ٰT�~���y^���k7�(0�qn�ڲ��Wl��=#U��>�����J�n�N��d%�x�����Rd��;"3U�$���S�ն��o559v�.���E}�S�{�0Vn����N�D����e:��&e/e9��M~���;��Yv66�*��Dx�Fp)���J����՗
�����|q˙ɞ�p����F-�y�(��{6��
,�dKg5(r�0Y��;��;����8�$Y�kŖ��8l@"���9��݇��6M����i���)�"|�Mh�ҭv%����Wd�	+�ӺhOR��%*�84߅N����P��Z�ԙ�N]�/YH���5���16����������7D�D�ϙ�H���)�W��^��W��)�*� ��!�c?JȈ��*�]���{[���*�p;O�T^���{�&��e���R�Wy2��@�����-e����\L�@+4J��
߾xBAӒE�n</��ˠu��v5��!r�YL:ӧ���Qș�7� ,z�}}�*r�%P3��� �! kz��� 7����ӆ�9Ä
Q����u
�t�p�43�t�A&B��m�O�L��x�ϥ"����t�1�"��\+:�aR�f���E�S�&Et?���a^����P46/&!r�8`��<$�%�O��7~�,��̩DN���<!��Ɓ+�m�A���?�1:�as(�^B'z�c��݅:c?����E�ab���P��m�JI�(H՜���=Sޭ��3��i��[��t2�������W
���o�WS��Q��v:Ԡ��)��*.-�����:��vec���ܖ����A��юʆ>ϵ&6�>�;�y�����H��P�6��� �d�j�u^���Tb��I=�� 6�L6���$
�5b&�Z�{m��vΠD�P\�o@
���ݺ��%dֵ_4z�	n��J�
O��G�Ht��p�J=lЭ8Z{H[�-Q�F���k���%���E����MV�=*r���� �ȳ�>�����~c7`�Yx�<�����j�i#��G�)�������0&QaK)�$����@�V���Ȟ�Ii]ӑ&*\N�i�(��C�ɤH�4?�-<�yNI+\X��*lA��Ky&�V�]�E}�b�Ώ�OGQ�M�}���ǖR3KH��v6
)U9����pޖW�Tp{����ٛ�5z}���̆wF��� �~asct�"�oÊ��-Sڡ�3�as�H��a����ℚ�V����|�h��!���h���
O�^�:�|ȩz�j�2�Y��_�|�Y^��2�CV=i��O�$̏�Y 񯾧�L8Fg-�:w��>���2�uG�V dXvL�W͟\�����	kZ|��qA��h��8��?.1~�4i�:_B�J��n4�����a����v�x�I,✊��O�ϟ#@!s��NbI~����8���J�����GJA�	���J���h�MX���Hلe��!�|vp;��9)>hS�2����Ž��6��Btaú�Ax�| >��J^<���Ԝ�l�[�uL:�7�C� �="�>�O�Z:����$���9�aVʇ��3[�{��Hg�ư���`�g�%=V�@��I)�~��ǼHJ��f��*U,�_-0��>�4���O�FV��*��gA�v;�әD�T�Y�8 6���ݣ,72L/xN�o6�[�w?9۲.e/�X�'�llg�����g��6�S�����xc�Y$F,�f�=�`��t�	�kB��iw���9>��W�۟��29eғ�E�c��+�J�m����Pt���9�{M����'�a~�{����d��$�����U⾹v�#�N��MB�!�H7@{���{�Jr<�Ч�c�s'-5dPIMKPV���V���m�&3�;8�J��ǒ9���go�4t3s��]��X���b��z��-rGN��Kyfԛ�I����Æ���R��mS���s��ǆޕ?8R|���U��2��L7 �ؼײ|t*�J���|*2��
�q-�AaIu�<��IBj#N�K1�(����}:s�|:XWm������:*����������[9X��P��>̀��r`�Q#�mab;�6c�C<�	2օ�,mzA�EՊy�|���5b����'&K�AQ\i;e�٭mt<E1isw�0����щ3��g2��[򨶳_Ҡ0�V��Mi�.�p۴��#V;��UE��c��}�4�4kq��Fu��7�`-E�⎲��Pa��o\Z�F�g��釠r�#�>�5�T.+�u����C���9@J�$��>�D$�%G���)�׍Vt_m�W���?���\m�{1X���g޲��4�b�\�b��}�WvRSu#�o�]�IyB�RY0q�]Y��6��:���g:�� ��8��Cl��7cI|�jߺ����H ��3�Rޜ���ָʗN3)@Y"��Ú�Xu�7�(t�]sʠ�(�8���XU
�x���Wq��a(:R�i�Q�J/��ğ��rÂP��h%���@2e�F{v�J^*������q[����z��j(��i��Qv�C|�4�
ē�qgE4_U�0�'6dRS�SF�i��<+���.���v�Q]�״C��83\˝7~2 �.�R�6�˄Y؜��UK-_��g<����O�q8ځ^�7�&lDZ�n�.cd����c�͒}�"�������&���U��w|k,I�o"
��x�!�G�6l�[X5m$��������`ւQ��ר�Ym|aʅn�|TN��濇P��?g�k-�w��y� �MM��3��]�\�XO˳l�:	���.�WV[�$Ak�B���"c�����_��ZP.���:�E��0�E}����Ydfm�W�(wy�O�m�����qa�G�v�ML��֫L�o^���lU�u�0R�d<�y�F�I+��tt�Hإ�V�g�ZҐ�?�K)�C�L� u��ȱ�"޹�SF��0^IqYQ_<R r%��B�Se.q��Ġ�mԎ�Y�l9	!�N�p	5����[Q!�%K[��e`_��E��#��+U)=�XY撩"�CW�Jx���qPYF֘��	��Sۃe}���A���=��*��n.�����c��2-����Ȭ��e蓭�"==<�.�]<��KHe<3��2���^7&���~鸛9�f���A��S�h��w�?�Vk���!�&l4^�y�ۼxH[X���'����zw�M:�j�|���O,B�k�lb,���.}����Ģ�08���l"�\�����,��J�JM�Cx5�ܐ�p��?܉��#^u���⮮<|��)�;9�b6���g��Cpc9w>�#޹��gg��Ww%��@��2�po���o���n���U��!4w�!_x8�ϟ��n�:���@%N���O-%���:�j� ¹���o�6�OޕqG��s�6(:������=/4����Ix���4�w�,�L��L��~w{�$	<qb	�(�����#t+�x�u��d{J���ޚ{@��� B�U��$EPf����֖�q�:����;�E7u9Y� �A~� ��ΞH���ȟ�JW)?���	���~��ĝuz�/�O���)��*VqV����jSDS����������㼳����·|J���S':~�iZ��\��=��)�S����B�����+���Ro������̍Q���vٹ�`�cS�y`u}x���a��}`V��Ėl�5�:#t��IAI5�;~���X�_H�nxA�vҔ��ѯ'W)�R�@4�h��)��C�= ��jp]
�Wz��r2�*�e��hrEi�!/�v?�\�S�j,���9�Hf<��
�����ێ���(�5>�=���ef/���`��0�< &�@��������k�?��W���\��n����*���Bi�S���Y?��ﵬVB�4 �*���kyȦ�˂Gh@aT>�7�Z�sQw�"�Cu�m�=�&`0e!�~Oq�x:�x�|��D�ϯ�
S�ﲩ�_ Cc��zL%_S2���q|���0���A�.H�I�#g�8G,7�DѼ<0ZXY�R��,;��(�����&��,�V�,���t��'BA�}�6<�jӁ�(�C�=���8�e��M
u+y趟������]�B��?�`i�Z��:kXr5��~�c�؛��$��1��i�G6��uy��C��n9K��Ǜ����ei́16S�9-�un�:4";,�5C�߰5T�SD3=��u����_�����	�\��b�_t���ʛ�lT��-�ڰ+�1�=�Bp�i-�,?)˶� ��	�2Q�����_��j�dZ���4l#?����S*�l��e |pS��
�w����]*�v"�ී�o��:�{�Q�
�[�yi/y��E:b��m��B����&�@����{�cD�@rMed�fP�d����������q��02����[]
����F��Z+e��D"b�8l�!V����??��$D?q�Qk�|�!y��O4�3'_��l�i�H�X�Kj�)ke6P�N�`�Տ+[T�`���2�}Q��A+�[߿*S���-U�F(7�0�5m�@��|t�2پC`Q.��s�aתᇦGɚ"(�ԁ�3�^�O�y����>�� �`�C��Xd	1[�r���ɀ6������T�F`p�t����@C�E!�ۜ����M��a������{Wr� mZ�G����u_<a�i�}zݹ��y���O��C1,��_\��¢�p8xw�.�CWz�Ql�|'P��(8��CnՔaaݲ;�Īa����t�o%�M��'/�N������H����>��H/�3?���ac@���P����M���|�v�X�������>�B�1��<�wo�>B��jFKa:��!D^@S�˲9b�;������\�H�ӻڿ�h09 ?-����t`]g�R�~�n�nK�&�)G#R����'���~+��/�����=,A$v�2�epI��p���ìl�I��6+���{��}U�:b�5[ƸؙOqW!p:bc�r��J�\���2kIs��J�6�� 1PWq(��<�_l�������� ��& ���������E���q(#
�G\jm}�џ��f�6G[K.r��E�hl����6�C�0�B�\	�3�N�j���^^-�2.��,�l���)��Y��qX}ʍ5����du<�%Jn�EA�L$�EE���A�ߕK{N�W\���$���T&�� s�]K΢�Jy�7�n�M���ԇ�o\�~Q�!-���30�\�F%�Y\{Ø�f�0�9�C}_c�8����:��p�,ҎW�� �	 ذ3�O��Fe'��f��J]Y�?�^�G��9/E^ReO�^�.�.�;�*ˁg\+��Z�搓����Jo|�%�~���~�)�qP2T_}P����D�{L��c��""8�� ��2_�l
ľU��r(�e�O��Y�Sn�?�2sxa�Bޛ�����&G#�5�ϵY�)��j�Y���SQ��L#4�S E���U�S>g?� �+�&���q�#DB��ON+W*�뮞1�C)r5�-j��a��,�%5s��'v�9Lұ��H$�5C3O�k���er��w�Z�4�\��*�K�=�Z<JMJ�@�4�T�=��zSpc��_���:�t�l�1\�دf�"W��q.G<��Z��R> AGؽdv�J��|T��Ir����(�x~�-d������0�Y
��΃��ٔ���2CҾru����V�Q��̆�����N�`zL9�= �Ul�g�R�X�(T��w�p�}77����M�2��2�_Ľ��K�n����\��	�a%#��D[��IS����R��s{(��qq�Hbvl홷�����z'Iɉ�I��է�$I�v�v�a�ZQ�y�Z䭣J�����-�L
����$�E�jvIF8�Β���,�o����U�ӄd�}]_<�E ;�s�����!#����^1L�J�)<�.���{$S�tU��f����K�͢�X���WK��f�~,�; ��M��!=��~1�{��������c��+�Fa�fIQ}|ξ57q�6������k���R�ϧ%^2��\�V�+�3���bm�[�������5��ߢ��t#*�܈ދ��+��\�gu! EԾT�F�2��V�H�5-`�(%�R�^��Mܒ��e�]��P��p� қ=Qe��(��Q�/WM0�ְ'���`0�U���nj�撍X�S�q4��hc\��e�G�2P=�X6����(|�7��V�y~�5؉Cf}�����_j�;"x��m>�^E��j��ۖ�ʛ�!�-���ev��iWs��<���7#�������{0���My��zG2P�Vr8]��Y���:R+�������u>'���N��;6B�²�Ϡf9%�,a.|[e� z�]�"�>��7ԫ��6����g�V�z*3/�두�� ��NDڵ]��]7����N�Ln�v�ru�F8R��PJ͟��Q�F`�̦���d�E6xGr��H����ga�)�G�o��7�%h�!�o�L�G�uA"�h��ȵ����$����F��I����G��+�6���4��1f��杝k��[s�9�M�wM�c�c�U�ΝY0�!kcz���A�{��_Q`!����>5	���
O.��.��7�Q����>��{b���3A.��h%�e��!ݰ�+XqCۄ6��$�^�*z�(}���\�u��@b	�3OA���5F�ض���1{�$�̬֢�!	�� "E0[�(zѝ���;��#�G�=��t�0�3ٛ�ֳ�s�xi)��l�T�(���P�6���5�_���7�?������X��n0Y���ҕ�Uj���栅�MZ��Y������~��'3�M�@� �\����
�,9r�Ǧ�\��Wv��?�LPź�B�ॷ9�A�(�bQS�����P]5�E�5؀G �ӡ!LKu�{��#*��:3�-��	����Я(M�[4_X�VA�#��R�7rBm1���?���A.GR
H���t���<��r���N$�y�"�dT>��z�v:Q�	 Bh��w���h��� ̋�+���зÉy��n�,�oM|^�p�OpfM�ǉj�<�L�}�����=GI�S�D��I�K������g̀E��L��p@9�)~pb�"�bz����>t���T!�a��<|6�Y+�Y��Ku*��ɖ�w���r����A6^�Ah}��~t�R�W8y�%�Xx�
��E�����ƊRR��j����>s���I�h��ܦ-��+�`t&��O�g�����Ѽ��ZӇI�G�̅��~D��j�S}��_*�.����v��n�}�}�hU�}���B������p�zL����\�s{Q��� Zʩ�g�6ɏh�}�/S�Oٓǋ��7��e,(̫�U�#��f��p��mȌ�o:c�s��6�����7.%ڡ�[	N�q��@��Y��Ċ%/![��em�9l�2��q�9]lhK��I�.1�@��ڏ�ɑ��|ď��p[��<W!芾Y<-�Ts	�.��Yu�(�Hڼ���Lw����B�������A��Y��7�<q�k�)�I���� �D Ij�i�衢��T���}͐yv6JF�"��3z0C[�z�B@��{B)���o}H��/?���O��gLk�<�-��`��2�����\K/@�+6.L,�	��L� ��e�"*D�0�կ-}pe�"T`*N��',��h�S�o�뙵���D��zLA0\����#�SV˲fɨ,v�5���&4�m�ҋ�Z��������2	�d�od��',�݁�.#�GE�0��,:l�ʉ1��٤3q2�y�������j�{!�U�S^��1̌�v�w�����|��:ǉ~/g�x-$�`KS�ˎ�&��\��E�J�N�_��YSP���T C⢧�|#���0dp�Dْ�v�@�O�F�Ţl ��]�0��?�^������B�cYm½Q�tu 
y����� ���$�Ra�0u+R�s>`�<9�]��P����,.�y��㉃H�FlNw���Z�yPì���>ڰ�xZ���'L��}E���b:�G��=�S���V�2��7
J�SU�Fv���5۴C,����=o�O��ʁ�`.w�!����7��E��K�W��#K܏ޣ��ְJ�7�Ȁ�C#���v��ď��~ί�F��$� �8����<6QܘgH�Y��F�mqp1�ӌU��F|�'��>�����L����N��xGP�'��:ħy�D�ȧe/�%�EQ܅�E8Tu��6�����E7v�.�O�;k�VF%s�])�!������(v�#2�]�����F �t}l/�c�k�L�e�"����Ԕ|N�*���UxDe���r����ꛃ�0-�3�i��C!�W<ߌ��BGd��&xQD�oT���8���O0�",����eO�f��Vʺ@0��`&J�HN���<ϼ(��ؐA�s����8���$〠܆��9��w��rC�z)�xO}v��� ,W��7#Oݕd�f�v��`�!q��'��/�Gvj2�4_A�@ gႫ?�qXa�d���:�|�NVwh�T!���{`!+�j��՞��e���YyG��L�8�}�w�bDV�+���K�$ �m���
1%�խ�ʀl�I��R�^.ܽ��9J��-T�����h�Fq�nK�jc6y��i�\cHVP��Ղ�m��S�߆� u� ߅D�qY��`rmf]*J7tI���R[]�Z�ebY�*����x7�G�(���$ 9�Q��]��NT�&�	�P�b6��C�e��^q�a���EC����Y˷��v(����;���AK֎T���]�Z�FUVU_vM͎�u[��8������p�v|������Ŏ�-��p�%'ymS�{�S���1(3D�L�N���b][��%*e����XR|��]p'2��|1���+r&.�޴����[=��5�n���n������.C��`�	�d���R�IK�}���ؘc��ĵ�oҾ��$Ý��##��Z1�8�p>ϛ�+�֖�'�iGL�䜒��8[;і�7]
By�N��E6�"��E=el��Z7=�i���0�A�!����_E�#�����򃽃J��� ͻ`9Lw�{�9�q�5�sZS3���3�\�@!;c
�A��$Z��h���q=��7��mAK/�a���� a��5�s�S�2����q<
|��o/�+���`����-,��͗��;]э䗴�x5G��2��|�,�����25���x�
B6���nv�u�d�O}W��&��g�#^�HMvl�����qgU�L�|�G�+� e�!)�p��VVj�������P�q���jM#����q��ߩA��lzZ�(jx�� ��n�E����]0��������eX2Ga`!L%(�wDL���ޚ��̓p癛�"�
!y�Zi<G�����.&Ԓ���%_�.y�e+�� �] �<�����x���Bv�`.Z	b_W�Y�M1��5*�u�pH!�)�&�}������֍Vr���A�Td4(E$�*�[*k�Mp�2T��ú`n�_� 
���'TYp��p���g� s{�G��ւr����d� T�"����<�P����m�v��0С��3�����D'D*�����4��j��*�ҹ�ȵ^����5��~��RsBJzHc��[
,\��R��K��dƱhG�+ ��:�-�:����mS�c�����ZH�A){�z�܆���Ν=�j���Bcʺ��dV�z{4����Ex�ҫr���V,��Cz�h=�ޞ��1� ��`P)S����F�m�Jf'\ -!;ǓYd!T�]jo�L����r_�bFp\�.���P�zc,!hKS��Ė��k�\��C��T�DD��U�Y��k���C+R8�	�쇇}ԇ��q^�"Ul1=�`e˸8r�XӨު�afq�Y�;(��Y��:9u*0����xc ���iQ�%���)�bi�qB��j���@>�X&dw堣�ٸ�����UBf�NR:4j�V�����wSrȔWz���Yx��H�0C���3_)9�J�y�A+'�|�����f8nF�&%�@ƙ_Vm'���?{�_�g�@���ސ�x����$��\���O5�����l�\��_&�Q�y��,�WHm�������\��ϡ�a*ɔ�G�R|�	 4�w�1�5��R�	� �z9��~�b�t�"P�&��r«���ɽ�6�X�$��M�Q��so��C�zJ<3����fU{�=��W����p�d�rLnZ��l/-X��	�bD;���<��%�����F��E\VI���"������8���Ĉ�D����fbd�7P�A� �"0'H]$�&���w~�5(?n	���F�C,��ȏ� .��#tC,�6U�.�iV�l�D���Dv�	��������,r6�cl�|�
`��\��]�
���&80�^i�MWaȘ2�����G+�5�n�)3N;�B�`$<�GBSG�I+�.�/�v��\�͋f�E����YϜk�=�Xauо|`����u��ZZ�nߏ�ɧ#���J����(jSM~a�7]]jp%0�M2=��P�h^��Q�-3~��r�&{��o�U���l���>�W���$;sZ��|�,�#P�M�b:%��y$�L%�7����+�}�P�t�I;���\�
io���2��0�:��s{���A��	�u�1B���&2X2�І�,3�X�����&��8]��S(sF����P��_��?�(�q�C�h-�욢�˶c���b6�Y�	��1� �l�
I�2g�⦙UǠ��"z��Wy�\j+MB"mTn�'�9J�Z��������l���"E���fysw�"�<����E�fWh���@.���(��ܔq`�J�	}�iV_b�W�3�?:�R�6�7_�x���*����J!NH��k8��XU�p�|�e������]xO���z�OB�����v{}54��\���Pן\,��{yv=PC��y�?����PBNH=b�f�`�L'_,����.�?�T�o<���g�~J���i�g��@���2Bn|GO�ON.52�t��T]����ђD���ӽ�<��B��A3��iՈ a<��l0Icj�.Ƴ�#��S��O���d%�ߛ�[Э4�ìdjI.��I@�~���Q��a�������~b���{\;�Ik���A�?:��d�r,}�(�o,�	�j�Y|�%q,5	F;�,� ��,��5�ȹ��e%��4�Ϝ�E���4.���ٛ2��3c�9#P�
�l��O��P_۝��Rz�eA�f���-r�'W'�\�ާU�������ܰ�N/��b�c*��� ?�,��ğ=5w��@����hRK�_�R=��_m�N��	��,�2�S�X�a���*����f�gJ��1S9s{&�.r�
؂�hك�6G�T4"����3}�����aaPp�Ym�Gox�;t��n�ɴ����+�&e�����,�q�I\_"��P��X:�C�1��ʐR_�D=��\�p!0���Q7N`����V��
��߼򇈶�k,b�I���Ġ���9��|�r{0���z�N�#$�!c��و�QS����"�0�A{�z�Y���&=4gF3ZbD&%(B��ϴWL��7�`�`r���m�r�&gnf���8m>=P[WF\�[�&��P(��a%K*���J
���4�S�$��!v��G���X<������El�\>��Bv� ;��%_�b�~f;3}��D�
h����b�G|U����Ğ���hq[��졧n�/ڛ��#fu��XW\D��"	?�G۫� )�qv.E�W��@��P�7��Ca��3�͏��y�"T����(��D4$Z������\}�t����۫���C�"v\�d/�A4��t��+��w�&�����W�?i�0�`C�}�GG9z�@�X�єG��b�iJ�F�c"_k�>�b2H��K�e꽉걚�d�F��r��I�uM��8���(�^L2�(�U�l� e��ЂkZ�{�ꏅ"̶,�$Wn�F�j��:8X��� ��%��R��)pt��_5�aPz?upv� K�+'��V�Z�bf���ȢwpA��W7A��+H��{U�f��L��Rq-2wUz��ӼK7�F̀�D�w��]���T��2�f��4@�C���T �����d֋�As�1�վ��P!b7�ˠ��̹�7d'{����͡�)���r3���e��6���u!hX1�)�u��^��D�5����3-�)�+�B�2w��h��k�e��}�n��r�=���Gpc�܃�,)�l������e1�`��y�X_�7@������@D��%ߎ��k�&u��H����p�+�4��y^볯e1� ��Gf"�D)�۷ɠ�}��ҬRN�r���4�ܛ���f+�~��|�߱$'Q
ƶ$�����ԭ�΋u�
�W"�S�\
��yk����j���-C��rFa�1�j�7�-7�d0�ؙъn\��E�r��k��ߵ�_��"r�����Tl·[��Mx�3�̺C��8
�05�b�>�(^˞OɖTūd\�1|U<#/��8^e =3��#~�j���
�0����T:�~_��3�L�M�?�˱g�
�~��8�~�m��eۄ �"���!��{~�&O8��L�9w%W�V�Y�xo���$��j��]����+&$��\�D<���黴�0�����D�<}�2���Grwl�� ]U��� (c�VY��|��|�����ld1ͅd���{��{�E�z�m;�#�+x@T�EǷ�vgVWh�%�Z�� �yn�
8�~�]z?i����"'u��GV�W�Oe�`��>����=� ��H�=��T�eQ�i'����cӺL߂��� nA$�g�1�I��"ΉqP}�j�c�H�,�"����A�$�R�%�8g�)g8��U��Q�gM�(�|��}0K�k\�+�L�[�hNTÞ�TĀ��q�tn�B-�=6}e-�d�]���E��"�#��m�#A_㰯d��X����4�^[:�[���!��m`�WU:Y"w������2�l�_t2^��z�+��i���>I��R��e�l���6��1�0t���a�uqy����	h��d���*0�g?.�la�?�&�����<Ęi X��/����a��滜��f��і�r[�t������i�j[�~Zr�	C�J���s��GG�ci�K�3E"���M��'pq9��� ������n�a�?e�s�Y5Z|���A��Rޣ
:Ox�H\s�*�T'��g�xVE\6��	�f��b�h`:f�qĞ��^t�}��$�Y^�!eJ7���,!��Y��ř�ĸ��"ܯQ|�:gc�v�`�� %N�+T;L�ͅ2�eyT����8ޢ{�Igf-F�"\=��w'yq�0�2	�LX�X��D���=Z?̼��s�^����l>*�A��H��7w!F<�Q5_Q����t ��d����!RSٷl���ķ9=�fn���v����okRБQ����4�E&��n��-�)�K���Lw��f��jД c�O�4��.:�.Ac�����*�9\i��kΙK\���n	��b�I��0<�R���̒c?*Y���	p����6��t�}x����rsO�t�޹�i<��S�u�"	(&�RtQ����r�g��i2M�ȵ̝�Y��q5Q�د�R0*�-&�t���
'Oi��RNJ�3[(s�nw�Fﱔ�U��(�t=Tf�9���{��ΌNT�*�`�e�(D}���*H���\Pf��Yo��@�l6k��S�
X.M���Px�8t�<.-O�Yxu�	�z��,�:�ԭ�%��aP;+�\N�F�*�iP��a��8�R��>���@ͪe��< �P'����cQ��ӽ	|fS=�Hʓ�Qc�I��i��aR��X��#�S�4�^b�Ui��b��b�������{U��/�4�Bǽ ���G�����Ӽ�#�����`�l��*�,;tV|!������>�X��)�P�˂3�AP��x	�o1���S��K���Hh�X�r?fmKȮ.�݉�a�Ԋ�x�	o�;�������L*�<��6�o��í-�_ì�5'˯����=ˀ:Y�&��o���������mS�/�p�:M��@VqC����qTvPF��Iwf>�1����Q����]2����ʼ� Z�ծE�&o6�Z޾�c,e�i�5��5��S�I��Θ��_�.�"v�	�)G���H��Ľ�Qb�B?L��l [{��׹F���ZnH��De��`�x����ήS��{��;�>?����*�e2�ZL�RhV�l�h���ٰ!��x�{��N�=j���>�{�Я#�.o��^2�ǌ����I�\�S?-���
���H���'~��J�M�����s!�^z�WS�W�G�%��8��r�/�X!��c�k~�P��H4�K�ӫ;����l��+���*@5�f�r��N>'��l H�(�Ջ��f����:���B������{�@��C9?�%OE�m;
��d�\%%��� ��:�~2��l��n�(�Zj a,ۥ_(��TIy�?ȗu����+���S�,S�^F��;�s���2�ֱ���còiT2����G��BN�@t�[d\��4Lu)H���#�N6���:�W�X�Q�Џe ��A)����͔��O"7��'��F��hּ�FgL�%O;�,�L���=�޸��(SI_Mt3(硊�X�T���b�[�TPp6�~�%��ڇ�	2qt�����aU,�.��V������æ+����^Y4!I����P(���:�E���~s�����#R����m
ĝs&U4yWd�Ĝj���x�(��e�{T[�_�u�(��;ϕiD�S-����cY��\Q�G����Fy ��o�׬� �^��D������7��H��j���2|@����'�o���q�j��������_�'~;8&�W,]"���i5G���a<Q�v{5E8먺}1|�3'!h].�)��1N�$�(u��o�s{� �(����-�X2m�E�M|�M�Ô��{������%'V�|x�>A=X����Bf�QR������M9�}p��Qȷ5�✚��շja�D�������,S��9P,���ة����>|��Ӣ6$�XG�]��g){�K��V�곯��!V�|�c�)�Q;��?�B�X�b����f_S�h$�L�?*h�D" ͞�@�X�E`[I����}E�=�4a���pn�{>361�_C+Y��o�B㢵�9����'��7�9�P���[������xd]�9۱�����U�����4��O���xk�	�տ��!_�ԡk���m��}0��2iRL����p���̖���cI�������C�h�ԾiK��جC3j�]�M{�ؾ��V
��L�; ⁻���	�zR/Q�1T�hJ�[l3�J��ߣ~�9�f��Bm�z����2�m���_=��B4|���:�bShmW �->z��A��o��&2@E�Q U*.*o�d���ݖn�� {z���<�q�C�0:^�n��fw}sr��e��j�i�B���=�d��9��p#?$�j���[V�4���W0��e�1����z)������ Z�as�S�j%�K�d��VL�s��VT	�=!Coأ����D�j���A`���|X�n������=@:�Aq��)����F�$]�8��A�y�6OdZ�F�>i�v��ғĘ�f�$�9�Nj��v-Vm�*��F�Ru��k�H�i^v^%TL�w�̼'@����?LMQ4�BG��,�}vHM�ϥ���61U٫��eRz_h�5�z7���(Ś[2
��yS�p��o�X��.>G[�U�:��*#!z�+�B� �q��G5͔��ۃa
c�4������=E�}q�0��2u�~��MR}��G��
�J{�G���k�_[��f�׾'=�����w6�-Ξ��u�`�a����S  z=�#�R"6�U�>�,�|X�xN_���k��6ߴ��9/���$yX���e�s�*�#bI�Y0�
��z�$��z��Ò���m��uB���� B�YԴ�p��xht?ե qu,��'"i�3�#�����eĬ*�$�$,�9Z��	5��?����� �����uV��v�,���u�5]��=�ra�uZ�
Jm���9w�p��8���Q��Xkg.�Ꮂ�+ba^����5p7�b%� $���u���p�9���Tw�&D>�$��,��@T�k����3�ˈ�+T֗�u�#`SVHA���5m��/o�~#��":�v�[�Ѡ׼��1n��o3)������u�!��g����G���(�8�M$�۟'��2�c��)p�)�7N|'_v���g��:��
�Lu����f%�ڠ�4A����ш��w�O-�(J�w�rB7`����!%DU�M5��8��v"jF���r͡�2mK�O]�Ɇ(d���Y+��)�����c��zYF�(�@F�QnBn��P ��/!"���$T�6���N�������NA���O�I�"ѸPUF�<n�B����ºg96�^��(�c�c�DƝ�#��6Em��S��F������B�E�S;��; �����(�ҝ�Vo�Z.�Q#T�R21)�V�g�OOO�?bR>R@���S�ңOd��&�����$��(*��H.��f��6�i�m����ڱn�Gu�hw���[ ��F�;����x� ]x�#�S�!�;�!/����$��� `����-Y#�mȠJe��+�L/�	�����M���-Q�4�P�\��àc�Z�j[^�Hi&�Zff��ސ[�y�re�P��Y�3�;^��)E�x��:�K�)2Ӹ��K�.��ǋ�������T ���4�9�^Ҿ,L�u�
���[N�`�������s�hTwL�+�2Ih�@7�'C���703��ʚ'��7�BU<�l:f߿r�x�ʒ�FV'�z+��O�4،S��:H�en[��g�-Ѓ���=��P�!����?oR���&�[�ԡ���d����pS���LH@9�*��v_�<?8�Gȉ9�pZ9hH��k��<���UT����;�yy,]X�j�'�W�&ܰҋ7Q9����r������Ø���A�y�D޺���QIbP@�>��t�LIo#m��I]��`S�<ăR�p`g��C:u\E�Y*Jw�Q�z�煺�3�p�������A�Q=඀FA/v��;�\����
��W�c�!Pt=�#�Ag/��Ru�#*DV_)^�v&���EA���}o :I�KAU�>o�2Q���ct�*Y����<�/��0�"RN���L���L�n$W��@/z�� p;l��h����
��}�Vn=��~����XiY��> ��ѷ^���۬�p<��Z�ގJ��C�� �9�_���y�xA�e�&�Ȅ8d$��{���BJ ����������N�N޲>�͒HV�]�m@�쳛v��ˮ��Ȋ��K9��d�&1�(ኟ��B��2.�yv�������P��#'�A1y
��v,A�ɥݮ)C	��% �{֟)_ߓ����A5? �����lf.�?Ц��B�D;pӾ��s�ϑ�J*���Zs7�t�<� t$Џ�9g$�΂xN�9;��ٳ
Eal��	����9�<�(%��XGb�ns79b �v��oR���<.6���Ո+3�̶`�-��R 
��5n�����/r�d�f��-A��Т�g P�6B��*���K'�<�%e��֔�L�(`5�G�BG�r�%ъ�x�ͽSDrPv���f&m�J����B��l�!N/����9l�)�%Qp�X;�]c�%�f>GA|H���؍��.I���o�X{Y�h�hTё9��3�u���D��}���5B�%䕘:�8���.5B�5��>�C�� ��|�+��:�?O���u�1�Ot��~�'�J2k��CYA��TC�m��E5��X�l*Nn|�D�Nښ
K,e�d�\l��/KZ�'�^^���,�d6����D%p����0���I��l]�	��3��9rl�r�	�����se�O�g]]<����-@�n�Ǣ�c��z<I#^�qz�쥪� 鱈¾*{�^H�EW���lboPN'޳��O��}p�_�3X�5 �5����]���>�9G�ë=l?����Q�%kf�1QgG���?V�D^O��X���R��Vhf�찀�a���?O��v{�b8���c�i���=��F������3e����T�s�3>��D�OZq���$j@zC�C�@�:E�{�ڏ�o�E�rh1,D\y��s���D�u˼�����ذT�;��|<d{s�¥�Jω� �V���c�o�Ac#�������!�8�J���PO2�˶�v���lk��"�c�����h8zd>'��G�����n���rPHp:XL��̐jm5{�U"�[ �;m���"�M��7JP�](}覃��&b	O;Di�ﮨ�u�q;5Tݹ�z�{
\�؉$�?"7��YyG
S�/�]��F���E�Is��� �MT#M/��0�++��8��9k��*݃�E��^JO�HrA�+���6�z�V�du"���	%�5�5������
��Α
!UZR�sV�f�On��Q����,���N1$��j��L�R�h�A:np�`�6@�ִ�`:��ŀ�J9̧��wN{�*/����kD!��t*����#�J��F���F`S���CG5���?�^�OC�vj�a���w�f�B����m�Qzzr������s��
J��)���T8B�/��/�����C�T.�� e�a�I��g�ɤ���<�^r��P��fe(�����g>�dxܠa�1�<a�(F�����x(����K8�2ˡ��T}*�Ϥ�@R�/Ȧ��v,�	t�H���Y���2�y+M^ NF{I^
���,r�����h�4��ԭM�칱&yq_ZD`�U2'���i�܈�b� X�U�*�g�����+ n�p�[E)�џO�r/��n���%�c^S�\P�Z%26��CϤ�>�Q˳S<�O��z�\� 5�Z�*����*Z�=�xn���$8�%��<���B�NC�	���0�Dt^;�\S����S�u��g��@����B<{�My��;�/KV3�W~��U��/z��R 	������O��q��F�ZD{hE�*�������Ӈ̼�{�rm	��%niU�x����w�unLl*9p�j�8�&��J��r$���0ׁ����UN&x7?*�
�a�]����-A����.�K6-A�ı���XH/��
�O��R-�hT�9cVE�ӫd��]���c^ o��L��
o��C}u/��d�"&�)'!��qZJ}�ɶ����gC�e�5�ܷ�0S	sP�3���NzYʓ��am�`ԓ��N�ۮ�u���M!Θ�p#JA*,V�U����s������'Э����^+G֡���h�o%�V�F�!1���ꂠZ�w�9���yK}B_I�h�\L;\i�*�>}��FU	����z���j)��T��=�F�Y�Y�l�&p��vi-_�Lo���������ֻN�����4�d;��Ě�o�p�%�ƿ��0���0G�9�	Y17�su�z��T[?����6!v����:�pP&����y�M�W�dq'.��#DD0Gn̖���^��$t�؞�m���4��9I�qɞ>�t�5�Mj��T��IX�P�w�MCS}ǋ%M6]���ʡov%ǀ��ԥ�h� �>��L�h���=H(�y6�u+�-v%3��nx�H]��$T��E�*FP�|y�jKx!��h�\*��ރL�Ⱥ��ͥ6���K[.�9�S���9����HѯNf�+]%�L(��`��=�V�7�����gO�����qk��dC>l�S*t�IA�0��{�"1g�:P�7{a|��P�2�e-�����X?�G/ò��^������B:,	��B��ʗ���QwØ4��� �~'���m��NbV��W�̀�����~�lV;��P��4m���I�gA���z�z��%�q�ؚ����-�)�ځT꛲�#��B����I�O(j$?�bn�q����0�ھH���&��a�V�u��Р�֏�h I��&�oW
�z��.�ݳ%���k�7�
F㵥�%j���v�}�~y�S�%�
/��u-nU���.�|���FTV[ڻM�NK��j��N��	<�o_�<W���d�#�ܚ"�� ���a�9�"��f�q�F��N�TN����q�=��.����Q�]<pʺ��PӋ�k��h%���z�v	��(*�#��o��cέ�ݭ����o�-6�����wJ9Z �����ll�Ǌ���$��z�+ɿGE$Y��pg��i�N�1����7�p���~�C������	�������c�ƙwEֳ�7�/"
�A�����?$�s8R$P�9��9TH@�p�y_�(����NS��_�Q8K��5��՗U9f�S-K$*�.��=���b~Ո��H�C�N@�n��S׻5�*'�x}���$�{�rh_|K6��}&}��x�z9��m.�o�}��� ��{=��l�bΤP�D{~�̳n*��
�J��ǻ�uuN��@aZ1�~@���'�v����}`F�������ԟi�s�3<�~�_�� �4��4�Y��]{�������5�����	*7mfa�.aX�\;H�4O�(?{1�E��"!M��������@~H'�>N6��]s�G�^�h��-�T!�v��+��0�>܆��'�e�p�'�&��c���b����*mA�a_�v��d��6�	��� M�`W�(�c#Ԕ�v3�:��y'ɡ}mTů��0�Rm>>��^<������'�-�KƮj�����]��De�O����|n�Y
�&Yϕfx0a�+��<���¬�od*_z}06�Y��÷g��dE)0�!��f��8p�(��V��ξ���ۇ&�2U�M�7 �U�D�ȧsi%P0���f�U^�����BPe`Q`��1��W���x�C毈M�Om���6�S �|t)���"���Q�!B8.Ͱ=B�����o:���j���[#�G(e�vرC����VE�\�q�p����u��d>�?�'�i�&|�ξ����-cK��RN��9�]�w�
���Jw��&�Ýg�z6̘&u��u-8.�����>��Ge1�������H�(������_Z��`ct�E�|���$W�߯��O;���H��o`1씟�JN�q���A�~�>,��U0B.SQM�tO���i����*�>J{�����G�:Rc�F�|�%n텄��DW��"���J�Bv����ُM�z!��S�����m��g}��B2�K��E]7��+�n����4�p�7�a��o�v�"Z�Ҁ8�E�1��t.����шh1
���J"Ö��E�b�E�X~��w;gs��m��<Y~|�5<m/���bX��ixvPl�c���q�k��z��o56�jeLHG�U5�/����UIQz{�s>R���:F�}��\�������>��s���T��)�3v�-�f(��3Z4a;m��=���r�OD7�w�yo���g�5h��0{AlŎj��8�o�5R����^�ʿ�)s�-.,�G�΂Q�:��,�������z��L�12�Wi�h (|P�i�ny�� Sض��꟎�z ����,�s�g4%	�'s����p�7LF �=��ku��]��+��WK������)���93���|�Q"1��%���Zɔ"B�f�_;��l�7a�ُkB�^E�7�N�#|��wK��ά����V�hd��"���%��s�h)��Ē�ghp���B*�+Bd�ñ��獸�9T�"�h�,E@D�ͨv<�����N�Ep�^��2��J��)qh� 3��+I^p@OXJ'{�U[�� w��2y�.��M�F�0��`%x�ĩS�>�:&���_$�hF�D��:N��ڊno*2�W����L�dS�dL}��Zb�Z�-��1n �M[V�Z�7�k/2ʬ%:(�d���Y%j��G�k~�n$���w�IG=lE.1�2��m�� �w�
�L8������Q�ǀ}lΛ��\б��须��?�usN" *�q�n�OH��=M��W.~z�:ּ��M7��-����T	��s$��E��g^$�s���l���@+R�禍V��i���SD�fHm����l��l������/����~cM��GLj2�o���kġv6[�^���}:񇞽�V�K�f^ L1��A;���R⣕�ʜ8b��)$�]ştL�$�H�b��f���y t�<@�/Cl��0����JA��*�m �3�Z� lS��#�	$"9�'1cSP��-�Z� ���h� ���f���<�,+�y�]��!�G<�u�"o��T|��F�y�Z0]w	:*^N��!��{A�݂��_���gh�+�Y��yD�>c����{�`��2�WYd�l*iљ���z�'[��Ӿ�nᨥ@a�^����z��%-�@@̙*�	�Cq���Z�Y������~��vou�-�B�.\���:C�Ԭ��eƬt�W#!�gU��$����˪|Cuo:g�e����-���] 1J����^XXC
x��UW?Z_f4.�Z�uc�Lc*����	��\M�B(���̞�T��h#O���빴_���C��qώ�z�pF�:}S��ў�X�l�sW6���w�팑���l��:�F%ό�/�����ƹP���v�'d)��5�Tj�/�3�&6XN^N�/<&*�Y���n������3����n⡓\�R��wWT,BWYr�8��wm}���� F�ޅ�Kv��{�5�|\��V"kD�������8sl���H�	�e�|�PB��=����z��ݪ8�Y�X���3ېE�b���l�h����Q�0+eSG��,YP���h<�2� 
1?�~����g������[�L�,�{-\�ʺN�@����.=��;v��(;��x1����R�Е�DRI%l�
��&��@��Î7h��$ϝָT��ʻL�架=�]<��u͡�>��->\_�eYɥ�x}�
7���X�@�W����7�)"=j�b��?|�ڒ����$t�g��|��5�ӬjuF��2ƚtE\�n�ۘ�E�R��m��܍S:�s;� }FEE�����4����E�,���X���h[�t����'A5YԲ�ڎԚD98�$���灜�nS^�L�R�`+eb��G�@qm��
+E��W�`�3��_ٓ�ɐV�Ώ�ڥ��׳��w��{�gۺ�
B�O��_.I�u��7w>ba��Y��&l� �-��-d���ȶ� o�����(���M�������;�V�s�R�Z������j�����A{��L+�k�Y�mS�16���������͝�9�4�\�鲁���R%pm=X����r�Lw	��h"�g��'�;��n�[�xM P���z�*��O���D��+Ig�]u�S�53s�sCT��E�%~���^���[��)%E<I��ݵ|�шwe�J��!�_���Q��*+
2(%=uP1�v��m�
�4���E��7!�m�ul��1�P�'��V�B�(��r�b�Fh�)�}�?o� h�
��� �3P��a�T^�$c�_�Kr�:�&+{a�`@E���dr'������&[!�U���8��~��[��!Ugy0��KEY�F�~�֡P5�S17=��4sV��`Y*0�e�l�ޒN���-���݂���Ō ���sVS��CPe�#�hS��y��+�Jĭ�z��Y�m\=@cB ����ڏ�C��(ŧ�Y��ؘSݣH��Q�ݤeu�=�C�u�U|/Lsd� �!�8!Ñ�j�7������� hT����.�8�F�N�n/��>��̰j�	~���Rr�p�M�������k��0` @��d 8��Z3"��]���(�#�C��f��S1�����=U�l�=�/K#��h��0K1���p�c���u�{ �yPƻ�X̓b�à��4�h�����[_��f���q2��K�]��1�c���~�H5���uz3����$ۏ�pX 9���\���)J���k�t:���0V���so#s�#5_���41��@��x�o��!%�z���j���X~1�@��k~\���p��]�s�Z�>@�3���t7/�}��&5��.�(�+{�IyE�q=�/������3�T���-�v�Q6�z�u�l� �7L�.���(#�O�E���f�?& ^�	�坆ጱ��ӂKus��VV03%���ȫ7���T7��4�RD�"
�FSȳ��*���1�$9���>��(.
��b���XЭ��w:�v��-�峑@�p�r�"�8�R�v���EH��`�{c�X,�Qz�v����iZ��r�<��^FQ`�S�z?'���M� �E8�k���CڭD�l�eY����%��} ��p	������k42L:���Ә�E��1�nk{��F�sH,�*�w�o��ۺ0�F�0��A�m�O�,w7\�=������!�3{��m0x�˒b����s�� =�-K�k&��3^��q؉�yni�VP>rH��;��6p��l��]1����g�]`鏁��G����U�1��&��K&��Q��,�������|]��yԤ7�Mz�XHB	�b��a��|�F��%�� ��4ߝ�d�T1ۆN��r���3���!�p�&i�*c�2��V���Rl�b"2�=)2"�mp�3bш�h��f�	�k(�F��R�3��i�p���,U���V-E$�O*9<�� ��l� �og�k�Q��x���9�����l�[�M�U���ɩ�4�2	ڹ�p�maY[�~J��(*���:�Rm_�Mt3DQJ�\��ղ�5��<<�%i������ �=;��٧X�ޅ(x����%`��X�ģJY��2i��r����f����z��dT`y�У2�ɾ{�˕��矔��#�w�|���E�k�<��9%�X�"����F���;������#�i��A�"�QIY�Sj)��v�n��!_����X�]9y�g�g�I�/,b��W���)�s����.�!���I�晋9�R�~�f3{����D�m1$I{��z6-汊���v�K0_[��¡~'XmQ�PN��`a.��X���VL���f�&����rI2Gi�Xy0]���%\]�!<���=�q�P5�=�z5>	�<�[��S�T��l��B�R|m�)|{�����M,+�VbP�z?�k��c��O��[[��Kp���H��1	C:H*@Ȼ�ۄ|̷ߕ'R�Z�i���?� �ƚ��}�jvs [7U��ql�@40�V�j9ܙ�g�7zS`�.	3���aP���s�|��}ض6]���c
�}�O��rpx\K@7��d`��6�#��0�P�HhO7s�ρ�nT?Vn�;��c�����A�" �jP��s�C���PAk���J�	7O\�1��C>4�eCM��cN�X����	����awY�J��7+�?��8e��P��H0B��x$"���H��ń��c橜�5�HR�=�̕�4JF�=}#��@Z�a���т�&�Y�K�O0�ו@��D
8VW۪f�*�x���1�Mx5�Ý�`��Rw<Bkep�~[��m�x��B-��Tutk[F��v�o���)I{ә��p�Jf;yu-dO����֗�kxf�dC�j��q�� �)i3W�ےD\ %1�E��:���Xx�r�bؖ۴�Ć!��<��6�_���5d�v�r�^*���$��|=���~8��p�4�|�4��:����/O�*acm�}I,�k��)#G.Fn<!���6�ZM��>�9`M�o��ޟo!�Jֵ�G�s�[��5a%f��;�ާjA��A�ۨ��`���/\�߼���$��q�唩��x��Q_�Iw(��z�՘�,�K{��sC������dR���-r��O�F6#~��ze�>ҿ�)t���/�ֹR:�b�ܵ�>�*V��X�q�p�U�s�}��H�,i��,#~Z�u.%Ub���B/�)���"�� ��LR֓��Oy$��C�Y#�������?Ӷ�8̲���
��5"��#�˜�3kQ�0�ڙk.�ʀ>Ոf��{<O��^6g�F���M�� S�E���)��d��d����^�,{sxJ	�ow��Eγ/6��Zx��k���M�A�o������(�_����S�5����S2��!��Q�}������#׿#���/����0<[���%/�=���:pW�+h�bb�0�����d��)��ٹ҆+���7t!l\����xM��c���)E�]Z�D���^'дl��^�*>q��n!����םM�nm?*I�.<H���N�>B���k;n�*�:Y��������i�40���K
sE�#��8�M�)t?Z�/��zш��)�N�+�^�D5�\`\Έ~'��F� �L[���� ��Y��H�r�-�j��P��Ӭ��<vS7�����o�o�~�'��	
F�ԛ�����!�/[*�߻fm�'��>�1x�+� p��A��!h9���pfm���� �]R�;��N���{�m���w>�L?5E/e���}ˬ��\��,����b�5��*�R��Fsi�� Q�t��p�t���Q}�NDHm|V2b���W�	.���B�[��>�8Rr�O��ɯ�yyҶ�0s��l�8�L:/#tEŜ��scP�JU�U�m��E���(!:��b�z�����\{�Uhw�O�`��~Ⱦ���#��"�!8<kT��l�M����΍��&0�v�d���d�fi�|�Mf�$BL�i�D!�,{P�qGB,i��.��}F�WA;�[��i�,e\"��T�A�П3'�(>�����)V��8e�Y�O�gq���0�:�W����p_��Hٕ���z�������˭<����.��ה�W���g���T���~k|�j9ui�0���}�J{�Jަ����:��>fzy:M+��s��a"61N-*�������OC�wӐ�_�1 ��v�A�9���Y�p{1z�:a�h��(G���5�4��&xM_)�:�ʍ,/K�F����!�O���36�P1��L@M~�Wh��ݦ�\��/��J`i�_��4�A���<�좵x�!�����Eх��v����U���������;�L�/&w��>,h���b����	Ά�|?-��T���+e�Y߫fT�Z�
N�|z�~#��Sce�e�a�<�7�S���)1'�iU2^�a�t'���')�F��ޱc����G���qFǪ���Ro*�cNf���4�:,2痍�n����sO�U��-����:Z9�(<?�ס}���,+�Cn�l&��i�f�XS���h���Q�j�G�,xB32��e���Љݹ��@����Hgnw��TJ�"r�������co�D���+�|� w6I�ű��P�@=U�^̙+TT0��bM���;ˎG!�_�X��� r�/,�"�3�t�C9��Je/1��r��$BT�CNN{��Č���Je�ˁ��IkJ�ue\4z4�3;n�������?bz�Ga�^��4���WU~��P�9�T):.�0�������|g�kld�$�FY��c��l�f򊄙�"I����e��N;���S�]%{Lx�s*�<�h*�	:��΋�%e�V�gR�k��@����Ѡ`l7�o"+,X�S�סך8BX�8�gV� ZF����A=�&%�;"��
�4��}h&@�d��UA�W�0����8o��#�k[\T�4�k=�U&����=������Y����x�%�LG`��ַC��x��l��|�ɐ�-�!&Q@�$�yV)����Y�ܠŕI��2���L���Iks*i�Ȃ*U:6�)4x��O��F���l�[dFLv����@�=�u���*P ���l�K��&_î7S�P&�⯞9qS���6���#�H��_���`b��CE.�-4NЈCf.���U_��i��!�F8��g�}����ý��C&��=Ck�)m�V�r��0��u����x��?���Q8����U�U3�9'e���c<ާ9�T0tº��G�3�S%�w�S��� ��ʪY�V�]�Z��tT�0ѕK١p]�X����٫:�Q���W$��澝��$�a�syӯ�qRPb�gd&��vVh��gc9�$4��B>[�g	��0�wPB��!ۃ�����0��w��v<ֱ�CD�8��~|lb�I��Ju�L�<�z��'������גws��?&�㑔L����j(g_hG�#+9\�ՠ/Z��ߔ�v3�z��ώ�������wy��v�i�������4�Y$ۘ^����?+�5��Y� ����9a��$��ßL�`�P�<��I�o�3�gt'4��y�ie�@/%�֩zɾ��?�{;GC��tp`n�M����+,)
PϹC$���n+�H�3��74^����0> l�m1i�A��c�&k���6�6���U�t�X�x�	��5C��J�M��^�)�#�����}�4uR�["�Λ���N�KkrJx�~@܋�����Ԕ@��0�R�"yHł��qߧ �UD�"�$�R�R�C��KkE7�ۯ_��Y�A��BVF��b�;h��0ϣ�z_}a�>�][J������4A�'��U+R�����M�j�4�S���@8%�H��Rr��,=��x��/��fy1��IwT|Ҋ�vG�31߰�k{�����hi�)�F%�L��;���c�ݾݳ���PS��=V�SD_���4d�E�^E"�J=��/ӷF�Q��ĕ��&J���b\�
m=Z�#��lk77���i��l�	���Q� N�¯m�����2�F/!�A���_���#n)��.*��]�ەU+E·�B-�jW�?�4��_�|B6^ �X^����3�9~s��d���G}�H�O�&���w���do����]G45�^�}�3�[|��`u=�����M��:��M���W�)����Q���a�}�<���4�I�y�V{�v��of\�Q��Y��OF i��{��u=~}���Nu^�->��,Z�F�Æ1��f�����&Cb>+R���%`�)LR�Y�3c���/pJe���$�'�>�j�fI�F�r<��~�}8*����q ����=�W���]���7@��n��k�8����z]š�J:0,N�����2"wui��n���_����jA�U�����i9K��譛�����S����z"��?Y^�,t�(�ie��36�p�Jo��Ӝ|U?��Xk	UT؟?�P�p�n������c��~/p��R�}]��o�K�mX�8��������w�%�  ���x#��yקF�r��{�{$�.��I��BM�ƯI_B��H��>Ü��M�(=�yi�%<�ry�p�gQ}Q���Zj��-�r��D���`�K�кɖ<��"�KB����v(!�	��K��S�h����D�-�A�H���)E@��#7������5i|:� tN��ƥQ���o�LB��h�)�N8z����Fye�9�Y�������2:��6@�Co����v#U8񘊀V�EP�����&���V@%*!��*>�88�B�.�Y���e��h�� ˇs�u+F��w�!���E�N�|i��GN0�<�Z�T�٠fI
���z�&7ah.8̎`1&E������.�k�)G�WI�o��ki���8QI�j��b� �|G8����/l��i�E���B%K;*��G8T�9�=r$�'M�Wc�в+g�� �`&����Կ��3%����4������N�l1��7B�([�J�ΑO��Ԧ\� q�zu�^ ܧ����G��bg'��Q�N��#h�M�����#�ΰ���2�qv��܁AB9��秋�sJN��\�ɉ�3���ܥ�r��V�K<��F�"���x����!��/�[bb�"/2�U���	�^S�#���,-Vjz�|'������q8���A ���U�
�@��i�S=�!OZ�ξ��^�!4�`m�͉��ec�~BhP�w�v����.�j�-b�zܲ��_L�ځc�b8͙�V}���d �}2aj���N�na`W@����w�zUJ���hw}�	���D����EN��m>I�>B��OR@�����S�qSb
���.�zdQeز$�61e���_1w�j�^��n�Q�c.�(����nS� �Hqkv�`��6��]1��u�g�"G�}\��Lw��-kDvچXw�!�N�']�$��9�i׷�TX��&{���9���9���Ol:���̉ȳ���Q��lV -1�T�'��QY4�x1ԑ��h��@sW��#�����44�u��QgHd�U���B��B�l�$��Ye�!�t3:L��b^Ha[��r,\�'�y&�w".ط���!���������D�fD@&Rw�Q/hσl��N�8�
d��J��3�c��
i����:*��z�ك�a�"b���u ^M�d��R������T�d�9 �
{Xv�{��g{},����lk�B��b9�����7Lj'�k&��}+1�9ip��c�N�[�2kS/��FK���
�Q>5\�� ���=,ڻ�I�s�0,g��[�>��8�g�69"��O�󾵋�/��h͍�'?���'�Mj���I���W���Sw�[1G��I3���$�}��x����.�s_�~�>P�A���T���s	�p��Ƈ^�pPU�,_�$�&�B�����gY�O��҅�%iAɩ�x� J���F����LT?k���8x���hX���Q�]1bcf���Z<,m"�4#B������)������1���u+4�1�9�m��E���a��g{m��KQ�O�g}�M�)��3�IU��<��A��Q,0���2�J���@��'���f����n+�U�x���k�&��6��Aa�b��㫇&j:�%90�_��`&�K\�n�H+����&�6�o�/ձ�I�@urp��G��MRx���g��"r�Y�]{�D���RF������?��0��A�o�8�8y!��bYM��� \Bn��ɍ�إ�
LnB?p�_�� ��Q�N?ka9+|��ꮅ�7[��擊�W14�ʽ�" m���J���DzGM9�=�3���d6D��W�z�����BU����0���c��Ȥ��!���~GJ��a���Nl�p-l#�j4ߴ��aA�e��A���o闠��kN��w��cJsBd�-�]n���ȆP��JS)�y\�9�=j/MwZ�.MF�����:�j��93*�_v��Y��wi^~֔k�y(��UmѬ����^���9�G�CD�0�[CY�u��a�����g��C����V�;��	�UmR!�T�M��]@�|Y�4�X =�/V�5��SS���JXυ�u��!,o � nd����$��f�.��N,(^x�8%˰"@���\�*�2������;�R|�u����R�")�jL�����+э���t�r.ڬ�b�s��9R��~����}�|�%�6�����I��qԺ�/��ye��;�g�RQ¿f2������p�9�3�ް2\��^X�V{n�;\�y���A����E�~ �3y�[.�`ݼ;L�99>�6`���9�C�\��l>��ZĶ~��Z�bp�V�&�ԉ6OjY���	*C���3!è��,���t|��^+ˏ��0��B0��`f7`9([�2�B����P�L*���t��>Ѵ#�i�0���Py���{>@v`n�v�s������Ϊ�?\�͔�}A��NGi'�UA�޷��mF��>�C|z���(c3����զ�o����2�L�!�[#�Y�-d�QP�ژmɈh� i �� �+L����)�S���#�D�2ËO ����RM�"p�%��=�#���_�\�-�Ok��,��Ⱥ��9\�K�n`��?pհɘH����=1��p���zP~2P�Eb!�)�O�H)H����jЮ�)�Rz�7�'������V;�0h0�y���u���9��r��'��m[a�x%h@_����z��;��a�B��2`ލ���.���h/zZ��^��*�?w�Y�H�P�h�C�����,��i�j�ՄO)�x~9I����#BM�#����ؑ7�8� ]ט;x�e<����!U:���:f���8�FK�I芑��3Y��-��S�T�MYc��`��SW�ݖ%����	��A�����[�fͪ��#Ug�V��5�'�Q�j�$��S���S׭����#G<>��:>��(s��z` �����f�I>�aѿ+����'�ac�چ�H��n��u�r����"��o�+�
��`-��ʧG�W��4tT������1|wE�ڏ���Q�whn}��m�G<��_@��z�?Ң�e��j��j��hx�u�s��D,�Rɨ\� x&>j�S9���k���gyn�R�7qL5�q*s�aiA�k�&o[����J�^E�&({��Og� J\�B�ǈ�����&�b�V�@�m�#0�a��Cb���6p?әY\!Qj�y���G��d���i9�����ȫ����ݺ��	�u��
��޺���� 3R,�|<0�$�X��xDfp�mr�ˑ� ��(C-������o~�KY*9>+-,�M���&��Sʬ��G]sI(�$}����+Ykxwg#�j��C�n��+�ߞ����5CeR_����pk�F��MGA[�8�{K�����n�74�~9W�z�E��e����u��;�~4㉓�Hx����^1{�LMZ����
w�;��$�;�C���!?�ʡ�|/3}��]�T��:����xo��*� i���H2�λ����2���!�pk�:-�m־?$S"��(��$���-MP�7l9������D�뮨����-|M�9��~�j��?��4W���Kd��3tF8�֮^-����n���&3�y���'B�]�ۈ����20L�y�M�q�� }��V���ȓ�Y7��4�]?&��٠ێ:!7�b6���t�%7�L�R�)V�|��u"˻ϼ2\?IB��*�#�<ơ?LcmB��u�#oAW�S�N�
�_�j8u�r�_���cz(�m��%� ��C�G�M1.M�����?*�I7a�S��ĠS�nķ��zu\w���r!z9��j؈�/�"S�ό8�Tj�_Z�`���tS��� ��a*»
2OS�X;��BQ�h�Hi����`Z��z���.X�W�c��G'��:&5��o^1�@
�j�a^VY$͘6-d.Q��\E>HV+N�����������bw����]�T� ��+��c���hEh��~�6	����f<���C��y��zuU��_!��5�1
��N�)��C#��a�-`Rյ��I�f8=��E��r�a�B���d�%��.;pB�"��i��w6֞���^b��&6���������9e�\6����,X^�-B4`�޼LЏ1�%j��:�A�R]� ��t8�ܐ������c�Nqһ"$�y�`C���{ǿ�:J4�яb)Gպ�����&m���dF0���y�=��f�a��`�5e>��#h�U)<�pp�_�[S��&�K���:w��/��Q|�<B?Z�g� ��,�}�8OR�A��O.o�[��jI��Ś� ����X���0]�B��\i�P��iDT��6 f�	��N�դ~��� ޵�[bķ竎a�)��Ԉ-���1c�G��Gګ�#�ʳ��k������Kb�>L��@}˥����)�ը:�ϗoqG����y���� [�-��l�R[�g��9��ۣ#T��`׈��̧����g^���C����q�v~�z&��mS�?�i�p8�V�=��\񎛔�H�����S4�gP��P>ǝQbǁR�_��ɢ�
.i��e���n��jmoE�֗����U�
D�$p����mLu��l��	�
��C�]SS�z��M���]A�0��1Y}2�eQYA���L�f$¨���$H���&�q�-J�G��D`�g1��n���+ʏ!�vBvTˏc��W������[���ZBP�pPD��VS��x��y�ۣ�S��{��fa�u ������ŀ߮_�vI�a��8H��u+^Dj��^�/a���80IW��`��q��M�t�~z�ѫC���ŵ�-EE.�2��t��C��Ǎ�lƑ �?��Dwp�#�9���Iנ(�YȀ�i�@��#���$����u�}`�cL9�<�s�b+V�	#	Si�	����-�g�X�@5t�7q��Mb�$ւ媎J����jԫ�PjjO *I*������0x�EX��&�D`w��}{Q$�L��'��̌D}��d")�s���Qi�������g�l}9�R#�!$\���VW���Z5n���?'�6;բЎ�>-�9<��f�mC�f�ٻ+},�&+QS�̡� ���Ω�R�����ϱ���]�oS	d4�5gtRK���hęj"H魣��l�%(D:���e8�8��3�]��:N�{��$�G��$�v<:Z���m'r*�豏m}�p�'���d�Л��g������Ύ�c����L~KO�'J?>���a�����vK�����g���!	
�8X�A�G�8V��u>��tLZ�D��E��J���:�JV����j?��{�Y�SC�2nΡb��}J�ޫl�8\�ȫ-��m�ɸ(���"���}阄�)���t'�]g��4��F��
vv�2%�s�GP�Hg���y��J�D:�9���\�$���|a�?x�v���b:{�k?�V��o%�|�"�O�L��Vn7�T�~������&'6������28��Ѽ`���6w�Yz��_�m�څ�Đ�g�����Ze	�R]�45�cwz�ꯊ���dsU<S��T
ڵ��~D�d���G��p�>�@D�.*�<�z��u�gHF�qh-�h��)��0D��mP2H�@��1N��e!h�E1�{#H��~K���K��w��NP�Jÿ�M�P�ڗ}@W����Y^���\���6�fC�*�S�7h�8�L꞊� �U94����`9l���,�gh0E}|/�)�V��T�sZ#���Veެ��P�6	T�"֡�|;qY�6i��Y��"��k�t2���Q��y�M˽�Bݏ̍i���_�1°�K��m�%R�Ѹ��s��ͮ{JEJ7�>�֚e�+�c&]� ƠZ�������^���a�/W̾� ���[,P���x$Y�eF<�x͖(g�W˝4#f���u�l������'4���X�m�Λ�����@������;�P�2a=����x�3�������U�Z��1ꭥ?aw�mz�#������O�L�z8ɿ����'mdp�@����� �=3eG���[�!���8.&:ϒ!35�v���R�^��U�H��y��hcI��u9�nl?�y߮�(����O�S2sW�/{=%��GN��{��0Ui�ŷ~cz��f���@�k�|E�߬Zȏ����v����i!d>���^�s���֥O[$�WLVs�CCPԋK�t�ԇ(�ot-�m�ԁ�[-ωe��Kѩ���Y��翚��)�;�����ƽ�L�M�L{�6r?�r�������qT��z��p��S$>եN��4�Tm�-U��?�̦��%X.
�f&�K�B4	��:*�q����ѫ*�.)h�E�#rJ���'��ţ��ׂ�V��A?���DL -��̾�]#N!�-���#�`��㗦Z|���{K0~ٱ�'dT����^��6��N�4���;bѪ��WF%qj]y�uh�y��n��٩',�#*��
 �����sU���>])}K�H��&�%�g荘l���2_vmxO1Sn��-ѥJ��' C�=�L�Ϗ�;1�����0�Q���5Hپ�ANX(�ɾ�*����U~�!pZ�=�/_�|7} �*��y�P����82�����%�q;���}��	1�&�JX)��bi{�G.Y�mu���R 
�b�h:�A)��ӡ����>
 F]*{@�jMC��z�S�|<b����v:�ZAĻ�K�Lo���v_�#�d���8")�h6���>]���ОR�w�]��u�n��%�����=*�z2��N`���[�pqڂ�G�*H����ژ�;����ͩ��qבXZ��2�-������ 1�ֿhʿ��$�*W�`����/_����nV������RS�(�i���4v�x��c^���@��/�:�Fn�N-����c[kAi�t�k���ڈMiM��E�$�dt?��2V�	Ec��L�6{;�fA�:v�pa���ca/i@�fq�GS=vsgp�DJ�H?�Z�G&��N:����4��Qau����'�	�G
�;%/�3�"?����A��
��Vk�Q��	�?�;<j��2>�Z�p�0[�
����G�n^�/���tR�_�D\Th��x�l�Ϸ���ǫ �I?��p�P8.���v���a<@��G���:� �ͧ�3B�S1]�=��Y���������`�A�7��D{x�^�c�|��"�~�Y�$v����X�Fޒ����|�+����bv���)��xM�?��H�<��6��L����M��{"-A�w���Mx#�w)ߗ��d�˄��!I�[6�n"��K���Y����=���� e�	e[���G��
�Ngl�:·�b�����7���h�HԮ����G)G8��x�]��u�B�r4�AT��#8��#���d?��r���p�\ی�Ee~´@�Nzn���<5��\��:DĢ�?����93��W��!<��t�����(i(��}�X�b\����V�S~��)B�#=��%C��y`�R/� }+�f�y(�
_����~��ЋD��h_�
���SNI.�t`��fhm��~R�f[���j|�Xd�w��f(4g*N兣d��t�R��OL�櫊~��D��ҳX�3LU�p���h�p(C�<`���Ҥ���o7a�)v�������Z;�P�� �|�{��NШ���W�W�r�;���w�㭤X�4��1�9v�\���q��w�ŏsT����4#�?F@r��1	�L�q�`Ӭ�6%M�0C%��W��S���
�g[S��H#��u��>6�3���`����1�[X��P��ݓSv���
\W��]��P���&͉��["���@�X�WF���֡o�6;��L���3pT#0Xq�9��^�<��Q*�J8gj	s�梽���Z��<9�E<�����
^y��L�Խ|tl�M����Pɿkq�a�Dg���YHnb�UP�#�d]C�����?�7]��fX��˟6���Ϧ�����l��2�Ɛ���q��$ѭZ�5��O�� �ؿv�x��+l�7�HJv����;ج���W�0+0K�b]e27F��-�Gn'�/����;�%��!9F�zr;s�������L��'�=o���* c�WGv5�*O.f�z$��nĕ' A׬�����͛�����;N��N:����		W%�� Y�$@�E;!�j��<X"�����c��������z��|*�,kK-U(�o�j���W*��~���?Ɍ���)�
z4^u�0�9 �k���M�V��x[����z�i���r/1���<UB�<�h�3i�h�%=��t�p�*�FR�Ŕ�$��,�Ѡ	� �63���svb[��0���ս�	���K�/n_��Mμp�f��b�d�B�5n�;q)������z^����	�O��T'����[�!B��a���-���7i=Z
�R��_�lLH���C���P��;���*s(ף���~��|��P��� ��K�G؃��H���(>WіȪ�3_�V`cgwd`��M�3F�`������`�X��� h�������I��wi�b{�%ۘ"���;j���:�䈵_��
>��Ӕ�"���3*�}]Z��I�g>�GD	hvM5�J��L�ؓ�C�"?�����A�qA�%�zT�/ �4�i�X�P�Y���Y�R=�� �,� E���8�S�3,����kGc?:i��h걁���x0X-]�b�41��|��e�R���:�i��,L&HMp�Էe@�����W:`���<�1'戫	C+'�r7���@�҅�lr�b�0��f�L��=�I�9�q7U��6�0�Z"T��Z|͹U��o�xY��4�o����h��)���I�ӷ���p�Hz&�]]�
$5�Og��W����WY�{�6c���Z���^#��)������9U����Φ�l?��	�
�����o@o�g�q��N�[���m����0p텮Eގ���T���h)J���n��@��ÿ�Ie�CE�Z��%����8�#���/� zM�@�G����<>Q�]�@��V>��4)h��)�I�7���Q�8���V��F&�2�����E��FH_�D7�\3u��@�vY��F��;]�m7����M�DI'?�k�����k�n$�j�0�w�����¯��ףд�I�وK��t
�q���+	'�������ZE�o����ݢqr�vf�n[D���Kk&zp�\�ac�SZ e���R]��Zt�c(�����Q��Ԩw��%샨d�+g�vdЛ�T�m�ĈK׋�6q�Y�����91�(G��_��5fM#"�u]՜��Z����T8p#�6�Iǆ����ա}m(�)�B��;��&���w7��}�t��c�fa���S
E��q�wRl<�84�b� W�t�-M�,Lm��}���I�%u��̚���!�z�����Wc,�x��۱���MQ>]+��b�U�N#�c�g�	U#��Q��D�'��w� |}�&�;(R�(n-�ɩ*�a�:�����we6��9C��"���!�+R2~:��e1[�=7A$��Rp	��r�j��A�I�E��r�6A���2MD�V@�'E��=�W7� ����1oU���x�3SO`�f��������deF
m���wtC�ۋ���<��w·͋�b����L(��	�s��xTO�=1ږn#ޘ>�-�q䆟bRѱ(4!�@ia"�Tb�rw���(�~�~'l����9U>^mM��M�K��� 8���EU�FrB�]K��!�tP8N�k������&�{5�CS�3a�qCq"�)ua��w�#���ϊ�U�ȼ�$����{�'h��j�qFx�!��R`\�2�/��/&���'�Q�G	�, �܌���+�_�񓊙����C�d9�֮�v�8�Ĕ�*1:�|�a�c������ A��PA(5N�ڴ�N��X[=��*0�ʣ�07a��#�e�M�:�c��8Oo�!~ ���g����ۖ�o
��s�i�$D}Q?B�,j.�_݃2p`>�~[�(��>vG��`�C����w?��R�5!}W���6�tr@���?�]�M=��v�y�Mi�Z�c	()�W�:�7�JgwPj;2t񬧸/d2��sY��/��M{�C�E�X�yf�b���n��2 �K��0c�-&!p��$'{
j��b�	aK�fC�o��6�Z�.3B� y�cU�K���[/`Gx��=�Ʀ�0[�0i/��bg�`�o��L"gTM�p��sP�ަUM>�MT+�����S�ml����#�kG	,F�<S�(��稉j(~�<<�^ ���Fg}��(�d)�a�0�}��U�_BZv���`0$�J]�|�Eo�#Y�_rx�t�"�,� ��^
�<�4[�-�k���'����򹧵k2	��{ <#��X�7�	o���4��L�@q���yIw�,Cs���g\�S��NM!����bh���ZW��2b�!8�g��K�h�>[���a��X�(�)��� =�`_���
8����2���S¹a.#[$�h��c�*�����Sd>k�D/��=@����r{���j9�$���`QW~�	�����=D���KҔ�4k^>�� ��иTE�9;���?T
JcQ g$j����G�,�	P�/��%��:�Оܩ�z�_H����Q띴)�=�2a^_��E8�1����6���-x��v��xѰ��P�S�T��s}�1A�u3O$�O�x�G<z/Ņ;��-%�
ؘ�OD86��[�1z=̨o����e"4���)��aF_�����k����˴�MJ[��l^����ܹ��(շ];q�C�Jچ�{{sdJJ�-I¸����\t�I.b^�=��ij��;z��As�㳦j('rʊ���wN�i7�c���pO1eO��&I!��}{w	䗾��hQI~�� Vt�sp��l�4�`�B�,]Jb��ghK����
<N�&+d��A�o���
 �j���}�]�b~CZ���$ۤ���w�����CJ8X�*���GQ���%R�\��$��9і�N�H!,�g�X�թ��@E�K>��)����2�.��ۃ3A�D*t�jR���S�yP��'?�]	��pA�y�M@���2��i�����f�#����$8Ȕ%[���%�J�e�(�p�B8w���.�pݐA�^��ާ���+�*�{^�_h�*z�;���B?K�Kd����x�;�U.��ň��\ q�) k�L3�bs��j[Đ�]����}��K�p�6{��}w"�v�m������d�$��T`}MW~��3XL@���ػ�d��%������BK��!���扴u�͗���� �w�P�k"V�x�Ku�n��G<Vv�)�1�H�v�PYY��P�+���A O�S�I��~0������b]��S�r����g�[cm[�崕U��E��l$���oj�4���D�._���[Z]\-�������|�|��v�tw��m�|��m�^C�����`�3򝿱?�t�� T�[��K���ҨӬ����z(W\�'��.��%z��أ��6�P�2�#W�U�~HEg�����zپ)P=��x�A�ԙ[k�*0msn��#�Nڻ�cVa~&J77�rQ�Tj%�M������B�8؀'����䐅�W�(��+��'����C�tw�=����8Y?o6�骠�~zP	��Ue���P��D�N��m�Tڞ�+�TI�8	���H]�m���xF�[q*������S��N{���Nj+=q�`3��v9"_�W	Q̺E�2�gg�E�݊Ѓ�?��JG�A��B� ��kB Ư�J�_n�L�N���$ $��T�9B��.��E]��O��l9�"�&�OD�T�d�>�2��yAs�*�&����H<�v =Z�}ZnߡN��{�K �1Q���ȣ�<���_{����c�8 �t�	�:���:ʡ�jǒhZ7� �K�&.Ӄ�J<Z#.��5�������nO�&}Voees��Mv$��C%84�_j��l�0�
?3t �6��_'�r������2�](�t&�8j�ЏC �ev��T;�*����`P|�%�(�y%`�=	)���r������TDC�|@���֜�qfO)�V*&�3�Fo��s
u�zC������Ք?��c5q�����F���Guդ�VȠl��!u�~Be�`�f��m���
�4�Ԕ�&�ʦ��>|��BVh"���4��L�TdY�s
IR]	|�d=Cx��+�K��\�"��u�6��'M����!���ɠ*�۩�i��mp�� ;<�ZQ�'���=�������[���Y.2<�c)K��Y"�P��D��U�.�� ���~g�.�����_�P���j�6�V��%zX�	}����FDm1!�bN�p�G�\��8�v��CS������n7+�/��P���UE�>�t�g���,("�.7��d�����	PQޕ}��C�R5�,A�PR�G�MJx2S�v�$�R��M�}����+�i��ԙ6 �0H�e�^���,$��ҵ(>.� ��5�\�ܠ��-N�P�(Ռ?������'RV�1�'K���gKt����LAzِ=l#�߰��ͻ�&�;(���V�5ޣ��H����v#c#�8[��
�Ǽ�2�%�JXڬv{:nIߢ��(8��MΑZ{�
DN�W�b��4)���X��5i`��[l�G[���?x�3����.�ݟm�F��SjkKD�ѿX�\YM0�os��4����6-��Ji$&���X^�qD!��L "�8���"�?sI�A���1�Đ���0�}1����:�^��|�(s�@j'{�^/b{yU�����=�=���ͽ[����u�$ �
�-U���,Io#��E�W*@)W���F-1��~kR�q�4H�7��6� D6�*��u5��e���E�v�`�{?jb!��H�3k�yFm�ȂhQ4ᶥ�#H��}q��}^�N����e����w=6
�)c��ϣ�w�bu�=��-2h@��M8t�3��xO��~uձzS mU���i�@G�E��;�51�j�V|lb�d��?��[r
���[������q~A��r;�%Ւ��� �l��AHmS���v礍�%��p� ���U�W���:��)�SUv&�\��H_P�^�u�.�X\�eo�H�`)vH�o��K�<����an�52(�a��B��mI���U���l��@�|�_�%@�[G�'v��Q/�%m+D�Od`�{4��!�v�lO��{1�-!���?�P��ⱎاR�.Ks�Z\�8K�����7]uQł5��%8^�r%rv<Ȋy-����5j��U8���%���3��&�/-J6-yU��{��TG9!�4MG?��O��.��B��h�����QPt\�5��gJ5gw���?�~Բ�xBh����(	J�ɂI��y��!#`�O"~:�iqhj4���2�FX�)�B{Ѕ���3�w���!��=��0(�h�'��2�l�U��a�ȷ�����B��ũ�X��ݳ�����Yx �vq$�o�o;��Q��O"&~$�`��\.���@��s�T!�N)1r�x���km[�Ʉ�	�?������p�H{Bg����;����na"�F�x�<O�`�e�YҔ=�	G7 �oץg��亲
ٓr��b'�L90-��������v�+A�Y��m���-�������F!z`�Q�{�$�C�C.�):I���O��5P���ž�5`� ]^R5n��;v�ܽ�|D�D��֮�QqAjH�T޻0��PO���=�?[�g�|S?tYl�6��@�p����}�k�#F0uJ��L�oO*sQ&@�z��D��e��������lN�ِ��*���K���eH	�y��a���
�Xտ�g}n?��HC���-�|a_�{|N$$�*���]��\B��ۃ@�?W�&I]+O����6/�7��~������;7P(rP�e9(\��!k�(ȩ�M=��T��dK��Q=���?|����G�$��g�g5���W��V�B}-qG;����JbU��O��w�O�^yw�w�#�[�A�g�z��qd�B�"��\ϫ�t"���]X�=3}��>��A�Ͷ����������}kN��U΄u��Z�����9����K�&B��Z!�{��q��2B�B閄��(���ICӡ��1���4!���� �.6���q\���c!�����!~��_h�����w�1��4E�J�|YZ�(M�(���g����a�z���#�s_ީ�V�"� �Ϥ�􏠠MC����������9zٜ_<y��p�R�&4Q�j���V'�f�����C�5�J퉻�A�U��iu`~g��SZy�-z�#u�]e�[.AM�_�mNx���w�,�@��������,9p��61��x�	�+#}ᯑ��ȆN�=�K*e�Hs�h�@h	94�p u4+�����
T�Q���{����A��n$�=��(J)���ߒr��b�6��p
3Ұ6�]���3���	����gZ��Y4�0���/�FLZ/l��8����i)?��O�b%8�_H��J������{���$���N��B5�������0��a����9�Q!b�[#t#~�<�yh|��JE,l����R��_M`n��TP&��K��Я>N� ��h���L"s�d����#&�rv�lE$�����
>0,�+(}v��߉1g��֊	��t���?�-��t`����o�'��T�	N;�W����`@����!�B�_vzx��ΝO��é\"sgG�a�&���7�t�"��P٥�Ҡ
$�X2[��i���L�X���\�n���?�KلQ[$i!x����xx�$���{S��!���&�r�sʽ�Nǜ���"�ST*�y��Hl�������Fg������j�u�� F�s&GFRc���MD���L���8�B���r8ǜ]����)�cH���Wo�<i��~������f�63�*aH���G��p�[M/�i8�A���5���Q��2ݥIĊ��\:_�ӟ)�@�c��E�t &�W�y}��a"7���)�/�	��)yEN��:�[���.������{�p��K�����������<g���H7+O�󦿐f�����4:��o%����:&i�z�����V:4A� ��P�F2������ e�M�к��Z4�ROHt2^$�B�~n!4��kS/�:���|j)��v8T�2��h�����I߳a���EW-���w)5*�%��	߳AY�,0=��F/��ġ0+�7]0�Y+�j$(��@	$ga�{�J��|�2���B�m����e�zI��a�|�Q+�8�;�:6lO���ZMO ����)��$����e,�B���
^w7T�P�����,YKw���!�c���f^9�! �MG$]]�ii�a��Dè���]�|�D#R�5F1h����W4�͖�q�����n\�y�"QaR��W����x��m+=�F�_}�/S�U/2�酮b��>�ֹ�N;���j�p�O�'�x>���c�9�X����YFvc���Ǽ]F�\�࢛���3�;z�*�]�6s�;@��&��l��B�3B_��Q���(3���k?�]#˗�Q��'\F��9���t����D�Ҏ�/�B ��7c����7�à�"�ѕy�G��n]\�Q�mD+te�,��Tcf�%�C����"U_~	�/Mf��Q��/ۢ4�l-�
��������qֹ���N�� ���3��npR�G�b_��L;Ņ�9ہi�Ui��"�/�	���&�/�C�%��a��,�v�[Uz'M��ؠa�ź�2f/��e���^|2��ǭ��?h%e�m��}Nw�x3)�V4A=�!���7j	{�a�-O�NCA��i�E����I�q)��&� rF��0Q�{w�a��v�`F!F7gΖt�� ��CZ*pV�}���������zz�>�*��͜=7�0�y��؏��+��� ����1N2���sa��֐�b	���C��kEg� #�R㗈�Cɨ�սǂFk.Q��bZ��;��"`˴�w���5��x���#��0�󔮑��������kY�C5�zے��O���{C� F����8��+�TiS�Pc+;/"�:�����Ö�YϷ/��{E��*�{5zDM�t�h� ��إW�ʫ�Y��S@�y!�>����w��V��-�p��u|���A���*J�fm[���/��Xx�����V��̈́�i=J���r��ݔcH��{�N�sY(ZR^ʺ4���K���<�`H8�)d�=2��kཁ���\��ɧ^~�XW�o7�s�;R�+cG�[��MRr+mG�͏�{٧���Mm�f ꙼:0˛5�̍!�)M�,�8����C���A�E��r���pa��&hD(JT5���X{w�r �}����4��]O��Ȇ���Ѣ�� �9��P�!�q�0a�$o�_�}Ҡ��g=�'�m҇)�i9�s2�B���P#�lq(^��Eª����:[��u�����;=kC�����$ޭ��v��Q�kXm`��ɺ��Byms	s2,�lHJ��+�z,��RDd�l�����x�~+k�|!T��G3WVNK���(3��p�;ǭ��� c����\�/I�_�ƳV�M�E��FU�Ѱ>����-��J����Z�
Ʒ�,��d\�r>zp؋����ΒY�&�c����F�ͣ�X����I��|6k��t
�C?��&<��s��Z����2���z�եCe��q�z��.�(X�
�"��+��JNl�rcJ;XW��D%Y�͔�e*��TSry�i	o��c��*���N��Y(䔃C����T�E��@�� �ʿ�sh�9�U@3�X��9{˗�c�����1T?WXK߈q�Eui�Fp.��9����Yi�
���+k��Jd�����NP�z�PWӜ��1H�#͛/�[��� �nˡa.8���|rB�N`��́D2u�W� ���J�y�+�xL�Ep��� �����HB�,C�SW#yWC�jL�vmF��ZH��1����A����t�5��(�:/��Gr^z���=o�Ǡb}洢)Y�2�'AE�5(#+�e��&�ެi��=�ƭ'2|�2qi���������B�iq��H��9�����	%_ػ�������+�#e���uY��nV9sgnTv<ꊰH�gE<��j����N���]�"��k����l���P�&4�*AA��g��1�Ч��P��W�S�������=�g���u؄�]�==��.U�̌�spE���)�;�~�J�5}�̄����hAfE��(Q) q�ƘY�b�W��9���5�Eg;{B�'1�P�2�N�
 �6������qV��a��w��~��&Lf��L��𱫄{7Τ����@`_ˋ�I2�/�����ȚJ��q-1>	�pVXs'_/yfX�$�>p�q2*�݂mx�}�+�\M\�]�U�f/u)����?'i�+D$�FK5���Pd,�>�Q
�h� �$XC�0����u��`�~u��7�m�??qr��>��!���V�bl:-��7˷5+o�;�O� �M�ƿ����Ȣ����kg�P��6J��/3��WNchΨw��Sg�5���V�G-�d	����.����_x9P���ǝO_1%A��t	ƨ�_n��V�_`�'�N��g�v�h�8��KE�d��m����{��p)�`���w�3�"��rb^��'� �=��P��iP�8L���FF;����P�eCF*�Q{3ũ��s�~.�p򈾒��/j��҂%l;�|[��
 [΂;���������o2�Ӥc)����Ħؗd�u2LF^x�^����(��{�ue�
� ��v�6�Fz8t����%��#�e���? 1I�E��9��d�/���S1{�a���dVqmJ�\����q���C &����f܄?���7�?���x��I!zATFa��^��ቕ{�V�j�����]��H�7��2�xǧk���S�ۊ5�)���Fݝ��pG�kE(ѷ?��^=y�CJo�=Qcf�ܛ��c&W��ӜC����?�&���Z�mrGW�qd������-�0�tv�l�6z?g�g�d�!�j�,�/-���q ��dUgi�j����.J����ʺ��:��;���ͨ8fߕ�\:�����8X}����?1��^���:_�y��^@��CwWƧ֘>��87�%��^"&ÿ���y+���������~�l�?���9�V�����HK��R|�b5��t�O���,���Ϫ;j=�k`C �.���2X����zxΙB��o��"��Ea�q�_س�	_�)�ɞ0�'ȝ�WJ��j`�ȷ��6�
�Z��l7�ä��i�~q��1z��u��T��ڇuƴ{Q�r��f��Ծd�bG���Z��,w�P��p]��	@�c>�U������z�u�	}�rdgsE��5�r��\���\�ؾ�mA_����:8��0�a48t]S�N����O\;s�w{�=)5Uf1'����r@��my�<��:T�\�ᔶ�cj��	P)>���y��D��a�;F��p;yv7��$����"f,��]{XC��3�1Q���C�B�b�W��nE�dĆ��9�D��P1�][L4rx�m� �w�O[�Ǿ�N��R�'�����&nJ�OW֋�5�&���d�4�������:��տ�;O�ˮ�J�Z�U�,�ވ�B�X��8�ċd�+�m�3z'�f��8��}�	��ҏ��Nvx�jqG�������nL��D?[g�jP/�)(R׻�X7c����4���_Vu%����+s\��mr���{��*J��5���4��((�t�e���KUG���&~n!�$>�)� A���
 h�[)*/VP����M��	}n��l���!��T��ꀯ�4�YI\iX-� y���l�	�8�Uc3.�n�?哪�1v��'%�VW�xbv�������ڗJ�c�jS�ح�TkcĳgyyY��Bg���u��_g�>�+�T��wS(��<��3�.���K4*R��3�vpc~Y��!�n��Of<P�����%��aw�M�L?!&�ݗ&4�Wrw��鬺~��2�ɗMK2�܋d%г�+��[� @�c	��|��<��9�q�$�ס���+#�����h��?55vnՒ䒴�t��IqB�Ɔ�q�kxE<�33��3��}*�sB�dH����?D��Q��x�1}v��j���}-��tL���Jr�HQ.P H�5�4hF���3NNes����t�wT�0;�i�&]�)�l��(�tQ�<��w?**лT^1HN��L����R$��n�Pf���{��>��; Z���ER:�ɀ���H�}�}V31�*�r�`A}��i59�c{-�I�\��3{��
Բ)A�u��V�.���M}�Q�fN�Z0T���� m�C�#�׉�C��Օel��Bl�:&���)Y�P2�fl�8�ܧP��֧�H�l�����ea�c��ϋ\��U���5��j"�����A?��dm3ev
d 2��[�P����	i}!?Х�3�K�M@���	��(gj�6'��������e�)�#�_1DN��������U�hѹ�~l��U��43VްE��-Y��+
�Z5E�8�f�~��O8>�R�������*(�~{�i�f2[U��qG*�M^ےs0E�\VSpu�?�h�/Q��ι�11�a�Y���@�'	8`!j����Q���7L����,F�ǩ v�=})�}��5���	%�����/�tU��B�T�HDR����*���p��/6f'�>bP=Z�b���sS�i��T{4�S������(|�(�v�67�U�M3��X��T�n�b?��Z�xm2䱳W H���`(��sD�b\ / ��~����&� �	�>W��P��in�E�.�����u=�ƕY�53���}���p5�6%[[��J?E�r����q��'���:��/-�!»񒴃�#��8n�uf�`�~n��O/��h���md���*���<�!\�����ƺ�p��O+?�,â|T�9Zˌ� �|�\�4���.=�,}b�͆��{�-���-<�p�[���կ���2�͌G�J������
�r�Cy���Ȗx��[a{qcQ}2�2 m�:fq�&��#ʦ{TM)�?��o��C�%�(MU�Z�h6�e#�}��6�q�����W�lXw{y/�!a�8�5��[����Ї��M��~0��ɽZ�B}�8�E*�}�D�
�J�"Ɔ3�A��ȯ"��۝lA��%~�W1.%�8Z��T1yH���ぐ����)ԧdk��P�����L��[;{�Z%�Ș-��F��9T���0���Fo�D\"{n�5�fd	��3�ec���}����Խ$MA� /�n�hx�G<�WW0L!Xȴ3��_(a��EKIeQ#��ϐD��ɾ��aag�q��Y��\t�q��3e�CA�/҂)��{�|ͼ=?��;6ǈ�|��#f<��՘xg*/�/��_p���6���z}�])}}䀙.Z�X:%J.^2�F�R��BT�ߐk����x�L��1�<k �.�D%��$tO��AZ䂚R<�������^�$��Ͻ(x����{��sR��\Gp����ݯ�/C,�'鰌s<a_<[޲��	�c;~�<s�B˹�W:�M�b��r2��oU�B��$S=3k�x�j��6̯�(|�L��Ҟ����di�]��Jm���	{Y+��m���|�4�t37T2��e3u�*��Z�/�]��с�{���|
�	a�^�C�^bt�g%��ڐ���\GT�s�3��D^2`F���}d$&*���2kh]-T�lp����iO�9�jѭ,*�QR'�\K�geɗ5��.v��oc�j_�����:��_|hU��Dsq+��V�ny��nu_�r�����j��W�Ev;�#,Ù�B�7�5L�<���Ml� 0�e��4���D�n>Hۣxa
��Ǫz�ӳ�Ig�߇�����H��/ެ���Ša�����ܖE����4wVu�$���C���κ�V����eIpz�#��3iD$���0��a�,Тa�:%��[�`�S��?E%,���b�Y�]�}A��â�O��B�ł��B�nP���d��sw��(�{�;��rj
��;��Ak\�c�G�Pq���TF �Z�P(0��܂������	Kx����H��?�q:Ұ�-J�q��ҍY�q��\���ԋ4�G�稅%2�\�~�L�?�n���xRxOMW��![���`%�ӷT�J%��Yv�[��P�s
���a���H�{?K{��Ӱ��&KĤAE 
���(��~�o�`��%�Z�-^��L�,�u-�3��%�Z��o��T��B�q �4���$1�+Hl��`�Ge��4�F�M-�|xm�9��d�Ls�Y?�z�N��:/hb�o���^NU[3zf�T�P߬�7��?�@��v��eSo�P���O�6b�+��I�;'x�%��3�%r
�f?62/����n Ir��{N��b��l���E;��Y[2��e��z	j6�Q(�z'@��c�aߚW��\"���~	O�jΈ���!s9_/zU�X�����a��%[����%�%����aU�sbU'}'xT6Jc���ظ�K"u�}��7
�	�*� ���!Wp�KJ7u�,�~��r�m�~k�j3 2G��Kg��r�����V�ih��%B�����NRl�$u���u�������[��e��Ϡj��i�;㽦(>�=3��%◝H'�A<�Uם~��~1vlv9����ӄu����:r�Wwx���_��2�tE6#5H��v���EM>�(<�7T�7�L}j_ufc�;�K�ygb�Qj������5w>�y{�w�����A����Bx�S̍"&�zS~��N���m�ui����v����xA��{��h���"ԮJk���
�ɮFu�(2e�[�9Hռ|�8�L������ղA��8G�K-<[�EI�=\LY�k0x\�5hNԛI�{<�����Xu𼔤dM�!";(�C���ǿ���m��'�P���	A�_��w�\��-'S�KF-��I��8j�Ű�z@�i�~�=�X�s����bm)����#]/�k�/�F`�4PP��o�J$��h�S!�D+N��W�i+L����$�<B�Fs�dz`E��VA������
�	ɬ<(�p�{���=�h�Ɵ��0zY�
�&�aS����	/1S��o����9�
&ǭ���3���8N�oo�?d#�bX'
Uu�{��`�(�Նw��yI�F2�g4�A�6�w�xjDH�D  ]�T��<�+�"��8�W���?eʉӁG���j�_�T;iG#��<�����GF�6�ž*�r�2���;��v�f�J�����qD-�M�yc�Ml;5�z�i�]iR9>��O������Q��|�le^�0���c�&%�Lt�sAUv��V��:c���V�<t�H��S��ȽB��$�s��&�,D�ֻt˷硵�(�40|����ㄓ�K�uF��AS�l�]�t�5���JM����p\�0V�}q=��r&�����P䲾R��t�@MEӗ�S�� � ���^5i_UGA�B(T����B�iJ�����Z�-){N��C�>��}���	�k�.��OBU�F�2N*�b����^���U�ؤ[;�g"O.;�|�3�b�j�A�r��Z�b���9�f->S���ϥ6(+�q�i���ժ�ޚg$�݋0>r�b����"C�R�t5�����������[ka�Ly����-��#�dE�:1�!�)"\�	�����G���2Z�p�*�A)���gB����l�w�b�L�{��o�K����~�Y�!�M��r�/�*����H�rxtm+�l���[��e�7z��K�c��q��Lf���+V�#�݉�v��P
r�k%�iw+
�9�7]�T�/?Ae3M�*��S�Z��*)�?G�"���g�	ͳE��^�C1�3@�ڵ긪�l�z^��n���A,�F�_�8m�س���M�����U�ۯ��(�Qg�j>p�'XA����m�$�!O�0w+,��R��\��y0����g�Ր�uy,
��Tg
��ȟ:����!�<��.r����=}��������s=)(i.��$|���YG ʣ&7�x� ��=ѱ�[ެ$+�32칓<��}?^�ѽy�Z�v��@U��;;P��-ʑ�jK^L��6 ���N�	�^��E�8������l8★��5�s:�%1r�����2z]�����[[�C���v��?�  �*�ꅺ�􉞒�q2�S�؋�>�I�H�%�&��u�vN�~b�唨<�� Ewo;��������صL^�*�`���_ �E���3+�d3��+�Q��?�)3��D����Q�پ<7��.���HٝE��m�LY�<x�0�L�\��e>H��l�<�ȱO�'���Z'g�605�Z�����=�(m�[4�jʾ ����Z��ɽ����0)߹��ֻ.�Jm��7⹫ �ʆ�W��En�^��k�Y)~C�
��(��.pR�F�N��!<���c��X�ʶ��qZ�|Wz�|&أ�M��JX8�c��ǉl�d��U'��H�]�'�Z���VA��5����>��T���)�KZY�(`*BJ�
�e����P�7�xzK,�2���ӧ�C�ڿ�����49��j~+$��w
�x�=�k�Ұ�;�.	���>�O�ln�?��n��&�t-��6$�xJk��b�D�u5��ͫ-��O7k�՝��*U-M�_5ҁz�(M������VzB��~ڸ�у*����3��Krxa6O�#������9��6+�x�̆FPM�� ��L]�e��	�'p�&P���@�}�|!!�t�a#����� �W��V�\]�_��
��ݘe�T���x��#L<���A��X)+�Y��k�h7�L{���a���?$2�1`x�p�ͮ��0��:ƣ�{:��oŴ׻�K��O`O�
V��i�e�
�~��v5X�^�=�!��KJ�Y�2��l�n���#���I� �4���F�%/�E׉�����X�՗7������ܩ�z��ƫb=ޘ��/�]� M� �<�8�@�|0d%���<��\�"N�ѐ�����|&�0#NV�ng�MSY����\ϡz�*g�D�ʗ�9'룤�@S���Ί˸�2���P���&���_�@k��w�m�-	�{n7���`�R��B	iq�?���ߎ4��+A�8���t>9:ɍ��YŐ���E&[�������u�'M��(�`�$C�,�'���,��JH�����N�A��K,_ԟ~���Y5,��D-�jAG��(1#�̿�Ʊ��<�SV��}�P@�^�Rp�h4�H�]F�����!'�$��t�C���K�o}W�!L2��b�r�{ƾ-�%��o��#r"2Q�A�A�׍�qxsz��Bn�P��QF�/g�����p�f|�M��j���BZ�L�;�A�g�E�'�Je��qZ���'T�S3�S�trЍ\y�]���]u.L���o��(�la��@�*Qdq� mF99��)�ے�%�i�����n��v��~�9��ʒ"�	�)C�WI$��4���[I�җ���}���dծ���B�<K8u��uD���!̢\)q;0=�A�Z��Nx��E��~x8��cL�d��:�(�^�mq�:�č�~YQ�xQ���g�Ԃ�w��4:9�)�G�a-��:�2�޶ۑ�NA����KA3M,2�{=��g����8>�3���~��\�aʉ�<}-���Ӆ�'v>��֐�{"ʬ�w�I�(Μ��D���h���-MD&o�-q�j>ƱxlU�)-��8�)�CQnh�at��M�
�䊰6�{r%��}au�4]
4�j��ݎU����0���\�)�Â{*E����ɮ�0�z����8�64MI"���X|,��z�J�����ޔ�Q�0�AH��a��Zg�"b�~[��-k���	PNJ��R��+$�B)�s�	������n���(6_�\�.�q_� }��	74q���=��ѝS����U�>������=�љ��O��ή5�/߉��o;�dP6�|RG٬����\*��O@l������;g��u�oLR���[Y�SE����a~��$�n�?1��E|4����Q��ps,�]�����V���_���2m�L�I;Iҕ2���ĸH�0�U�b��>-�]CY����]���Ȉ
?�S�ѽ9V����,e3|���++�"h7����m��Yߦ�K7Ed��T��-����5����8�G7X�����G�8�0c����}	����|�0��;N���8sR���;G��n{�(�IiANl,�A�3�� �_LR�����À����Y\:���L}ayp_a#� 1��BTJ1H�4tfڞ�c?y�L���	�h�{����qt�J�������S��pD��U�L���^1�&c��d�J���O�yɭ:Y9HHj���\��Y"l�3*��~P����l!32�Y�J?��I�1eE�*]^� mT�[Ȃ��)m|O�3~�`揳"�M��*%CU���veȻ�����o�#1U���ikL�gP��1�ʹ��C�,am�{`�ԃ�<���@�p�ܵ���{�4�%���E�,|�̉�V@\����VBS��H��[�������e�P0��ov��eFcpЏ3��A}W^����J���&��5A�⼚�� �F
n����Z|@�*Pl�2��W�z�LZN������/��aV8jV���P��K?�{Em��*��l&jxk�X��5�P��\�4�(a Խ�W&�Z�ΑT�I?nC�}�x�,�pR��z*��L����ٺ�yo:�M{Yg9v��꼗�j���Xm
�&�����պ3Mn�-)�l{�3M	# #��#�f��H�d�`�O,W5�y+�������^��}�[�/.���#��$����d#���{���tJ7	F�z�,�s�aw�z*hfAd�a��
S���e1�P1<V|NU�W��c�q���+�z?F{��M@�%̑n��}��k����ڦ�|�e{H�+/wI�z��˴�9 �ߦW��47?w�'S�H YS����0d[�E_��W\k?z����89سWʀ�=��'H�-;ϾjP?� 8��e.����{����L����y,,����|�rf>�Ӱ�P �c��&�_7���2C��h���
.N�8���'��S������Qʑr� �����ͩ�,	}�K�,�P�K߽� w����|9퍳��o�uh��/^�)0�{�
��D&v��������#_.@�a\-�ZH5eMzrY�i{>C����dъ���}�?!?'�������Kv)�GeQ�A�5�]�-W:?̽��q��b���;�أ���<��e�����r6؅z����Fr����C4�S�f��f?�MKz���M_��v���|U5󩍋+.O�����c�?�}��俈ׯ�#ʼ9����)B��W�����V�*���雸Q�� Hfo��֩�5����g<�X�"��v���E׉�l��_M^l8�:��QA(J:'ix�c���K7Y�F�]��-�� ��L�k���-N�rv���!�gi��k?\�#���R%��Y~��m @�>��Ʋs�ѝЍowcNw�`���_L�(���'e��e���ZSGg�u�ۗV:�sd���?����=�3�U���ɧ�q"��G�[)�~8}!�O)}���e�h�/��ӂ�[;�E'���\o�[#����<0�$��dj����^'�	U`(9��
�H�?�� o7
�6̤F�8�D�g��$e�6�!o��-�J�5������ۗT���N��駌���B�lL-�2����/C����6|Lv)U�KQ�i,���͡��y�&ȱ��2�2{F�腫�%�%��5�-�&�bԅ��i9P�AVh<: .���""!H�EӼ�v,2#t 4��� �3j��n>�K���c�)�PyE��{���_{>��7��ª}�R�)-j
3�*H��Ө��i��+�q�	6�\��y�#;���4�5JX30� v��.Q��(3��V�B����O`�S����gߒ��!��x��5���т�i%LC����ej�6,���xS���X�z��<��!'@e��`�i(�G��͇帾�w@����:	�V��F;�+���_���ᯜ31��u�F�=><$%<EᖋA�b��g`����fN<�!p��<b��1s@�q鮊�5��
N0GO$<[�'���$uՓ��v�p�	���2��r�!�E ��!)��)?:Δ<Ө#\4�i��+r���.��8�����* ���<.c_�H�?�Z���y#�jxC�HAr<u�ű���W�;����d���ֈ�j5��6�z;x��;P��e.��T�Sp�]I���T��Ѳ�b��,*���K]i��p��S��pY�O8�t��q@r��d�-�Uk�tE���p�Q��'�2�ۑ~W{ҠyDF0�5�����o��n$h:9�\�jd�����fS
a�8_U���	�r�Ǹ�NCi��0��	�����"F�*�Y�_S7��Sj�m���0.ʹ~�m�m�S�B=P����J���S�b��m�r$g\�8�6M��W���8 ��`�j�'��ڏS�X����0�ギ�Xf*.s��3�hpH��)<�,J�>��!��IE4�����rg�C����Y����^.�{4�p0|s3XV����֫I�6?���4?�:0<>���FPk���F]���;UY�: �a�'��\D���@WY�_}��]��ۦ���5o�O����N,�u�l$R�8�<V
��mMy�w�~���Jq�Hr4~���@���x���K
���s�,o�[~��>-�l+=抛�����g�K��)lw:�#�� a��U�uU��� _r�V�6oQ� W�G�eRlX�s���hu�=U���r���R/uvG�߉�i���]᧢I�dl���2&rPpU�������)���K��y(2�[f<���N��A;��	������;�$�x0�$ ��B�:$��:�˥����Y��u!h�K3
P_�H�ɵ��ekZjp�0�_�~4m���Q���5���:rT�X������~@��XH���52?X�V��2��F~���׌F�c���g��1�b�R�&�E��݀��O(�e=p�Å�j��a�m�P��L��6gݾԨ���&��X�dJ�ei������e�M���R�<$?iK�Q��C;�O)��g�d�
�����bD��Xn�+�ި�}^Mh�7�X�(��w�Y����f�6���_mt`r\�E��`~V���1}/�(/�L�l� c�^�j����l���-Vl�.�=b������P�K@��ׯ^;X#�!} #�����"�{��+��#k�W`�J�+�<1�̫N�Ļ�W;K(����:��Ev2b����U�
� ��i�[_i,�\.��k���8s�}o͹��G����*�+f���8�-~�t��ԃy �>�7�|���kC�a�"����H�D��v�뀝bgh�kpow�ۆ��6f�eUoE>�Љ8�k/��̎>���9Z�+�E��L�į���ֺQFy%y�̸iH��H��0��!`��φq$OLbg$�]��]�m��ZZ`_e��τ}/�<T�����+����=)�Ͷc�ջ��r�,�͏������@�+�_��A��"��I��(��G�6�l�����b/�;����LZ~���U�&�4��>v�go@��^�P��ũ[��YwY�W ?C��:���b���Hi>V/�bFވ��1ͪ�_��P0�u:S`X��R\�*7��w�W|&e��Wض�j������-���ULyHK�<����}:a��b%H��ʳ+�4?��d�4� l�6^.��=S�c�Z%.���qT%��1�k�JXЯW���Z|:e�xA�
�w`0��7M{���Ok�5�(m��.�:@�����x���i�%'���g�S@���@_nsƥO�Sb�.���-�%k���tX6�:>N�5���wo��2��,Ժ�����w~������K��B�QӖ����kFWC�V-]'Y���$n���p��r
F�!��fK~��^y�n�լ�Ȫ��D�ݷ�~L�k,�����X���/�y�Ɉ��|K ��;o��457&B&�|�J�Q����zږ�T1�;g�3Guuz���/+Y2E���vJ�dA	��s<�Cw\��z�,�C2��{K��.�Z�<b�&Q�'ʼ�OI��S�U-vu�G��Ԟ���)������3��,��̂dJY�=���F$�5�9��uC@86�\�nˮZU(�S����Vk�/�*�	q��a.�p$�S��h3�ip�n���F�,�tţ̹�j�W\]z�q���j^��^R�� -����A��5�M��]�������������8[�
�}*CvD5��d����Mx[���%�h�´xcx:^��wJ���N^�h�����W/C6=�gû �K'�P/h��G��`�	K!���oGA���̿a\�W���9��iȵ/��s��E8f��p�9�K���_y/���pF�C�T�DS�d��MĆ
�RR����6�sN,_�]�~V��*���|3��ߐ�A,Z�UMVKѩ�l�@���b�d㴻��^1��GnN1��w'e��巰E��1���a9*�|;��P�кI�G%	�9�L�>CO0"��S)������$�E��Bތ��!~�}Q&:;p �h�њI�[��Zf@C��ݗ����7�������S���?��.�T��g��!�l�K���z~�k���!<�uH��n*���\ڿ�8���J���&�Y�ͽ�b�J]'}<��ѱE���ק��u2f�	7��S���}��SK	�g��F���&�Bv\�������d�m�&5���ߊx����	WOl٫�Kp�6�ǔF�<uQ�+'c�S���&��#2���&��B�,#��@^��q>��nDibq]���Ḭ�i]9�FS�s��%�^�*����|8����_���ӦZ�>3��#��WUr��8��x*tkU�b�m?bȉ��>\�
�]<�4�R&�̱|	�S��<�x쬂��k�|�웯�j��㚜=71��N����_�����yvS�!�E�]�QJ�ۡ0�QS���� z�Z�N����Þ-��
���:��1n��ށ�e���^kc<~������K���� 왬�����U�yx^��3+g��H�ݴ5�i�h��_ ʻ ��O��j�IR�<>�5�9����J�$	�hxY�A����3W���5�Zv��%����I���hX���P��u��j�/�a��֛����S�s���>Q�^�����>�>ሐC]]2������1U��e��i�2�*�������v&^L{/�z,��H���DX(��	����o�Y�,�o48^hC��\����_������_��+L0�k��l'|��:r��yIue*ξ��|[�1��q�R���Y#�#66��
��@8�}V�n�������Fp��ӳ�x��Xl���*j��dr�.J��wL%��g4C/���^:���}N�c�w�q,<�jn��o=(��c4e��Ԋۻ��Y�2�
`KFce9�P����o|
�{�n!	����}Z��8�b*�{��Km����}�DK�p �^����l���8�[�=�(����^����j����f�&�/.䦂B
4W`3G�����wR�P�l�K�b�I��4f�x��N�̡�q�O{�tp^,��6)��s_}ƍ�5x`��.G����7�OX�~ச90� ����n�4��E4Ĵf�|o9s�i�m�g0%'}O�S>u#c���5.�3@L3�����؈J:��s۴�߻ZM�"���ҍ���H�l�׾�T�;��B8��c�x���VB������?�R��z#�U��A#����^��y��d\�}�R����yP)�kR��-�w���f�剕mCX����͇�$c�NT�%�ͺ�72ul��7�r�$_�	��m,>aBi�`?�ࣻ�q
&,��k�d��t�J� ��vpJ��}��\��=H�TX:g�a�V �Bw�! �}��p�#Z <�ux�QD��Y@�)��Y%,��jh�Si�y��\���I����A21b7�[Q��`G���W������� +J�~��40!�Q�G�q��"QP��YG薜$3�2.��B0q�YG���^¾	�vr���۩���M5���D�8�xnF�����c�(��U��Fc����w�鱉d���������(	����z����<[)�{�,�w�#ß��8�Bn�������o�HM�e?�@�b�ņ� ��<<�7m��ET�#��Q�7jY�9j��f����l�Ziy�dE���9���՝���a���f���!~�[��P;v���u�7���OD�I�q�q�?W���8���1��
"E��%�q� uB���32�|�[^�g�	m$F��|G�=��X������У/u��AR�X��'O��9�,6���H��<�̵3���Z�e�D������Ɉ�6�ӓ�<����!>�Qv��s
�Ѿ� �LL������q��p�Bر�v`,G������W���I�!������3FRF�,KoD3�Z7M*�@�2a�>�>�SN�V�D�v��w�j�+�m0i����g,�e~�F�ദVK�/B3y`�Έ[�.�*�r�a�.�߿��vKat��h����L�'��D�S�+^j�k��[uQ���zL	g9:�N�.�1��!���\���$@�x�	l%n��ibu���x|���uE�+B�l�T7�'�;�07�m���5_[�[�R��}	��x�S#Ę@3���u��tN?����~V�ʰ��ԭlà�Ϝ�w=ϭ�YQ o���`���?Յ �l}=�E�2�.n�u�з�bE{2�E�/�{?��P�b�;�����)�w���t�Klĭ�l����uD<"�����^�� 13�Jq��$}������/��8hz����%�O�nt[��z��_Zj@���8�<��14T�mb�smD_�r��{�M%7�:���Sթ31��՗h�}��D팻=��coy�v�ժ������Gh�؉N�g��"��2��#��
0��*1�j6FWͮ9� i����2u�B�N�!qd��Aep�)���L�C|<�u��)$j���uҲm����zk��Es�_������ �(��i��80!}u��~8B���k7���M�$g���
��D�0�YH�Bh��V������L=N9�2Ӄ�lF8�|� ����>!S[2��hU*\�;�2NkY�4dɧ�k�O��&̴QЀ�-���B�\��ńʼ��۪a���!�SZ��)n��>�q��v��&i��V�/�K��'��
�C.:<�5hK�`$�VA��g�O�K��]u��Z֭��y��+/��&���N��G��5�.���>��K=�Nҭ��eef�;�����gT����c�uq�p.Ѱ6-�;��
�<FW�c�V�pe|�)8��
�v:�$Ή%ތ�=X���lU̝D�P�����v�?U!�|���z�%Ɨ�`�1�	:��3{�w�8���_�E�F�Ch���ٓ�9V)-Q�?��g�؊�hYa\�`��qco�l�-Z���̍�^�K�����	t����f�����^�Ivp��TvVE�L��C=uE�4l���udO�+)d�)�y�7��ܧIt�֍�4�,#��#�(l{��k���`�#(�"��
�G���^�;��dj�!|�Z�3�M�_�������ڵ4��0���;ˑ����~Vu[LlR�}�%q��B���˜ ?�y�$1%d���=��{S0)'�pk� ���-��/5IkۻYJ?UFqw���VT[����_uӬgB�b|�`Y��r����2;)J�qr�˾�� |����)���S��g�#]X�F����	�y^dN�#�/n�c��M:�����݂����>��R�>�̄<1I�|��c�K]��p}�]b�p7+���Y2Dv��
G+/���Ȓ��
�m��G",��#���B��7w��1�WbdL���G���8R'��+ӝR��^��&u��C�f�{p��9X`A)�Si��P����� M=>�����d��U|��;'i[@,+")���+B�ڹ�̍y1p�M}n,�ؕ<*%r���r��,O��!��T�Wٔ� ҕ��-���W�HL�ܗ6�s��8�q����7ݳ� �b8)��������N�#��R�5
Y��1�������$�0gu8pU���)�;�y�͖����.������2��2%	O}��?�V�
�d�����e���ǨS�RJxuPF:.폗[}�����;\�<_�̮�&#��5��ku�)�����&�4ٓ�%��KQ$L ���4��kT�6OWS]�P2��C�� f��۩^k-���� ��
�)�;it�b삹.X0G��px���e?9}|Γ^�vi��o;���8��W��1���1�.����яh�8���;�<�����%fG�[Z�p�����(��Z�����6Y�ci�2	�m�"�W�P�Fي]��6��y�	o9��PP��W��5�h�DpG��T�6�k��٣r�g+��Ͷ��.۾�������0�j�{;�X�ڨP
0Rx ��V=JS9�V�k��m�a���Pw�!��{�o#Z/�]E$nww��_(�U!�!�[r�?6ZQ�t�է]iY���G��N� ��{����:��ȅ��ԥ�ƁlK{:�T�A�?�\� ��(xz�
a��e�خ�z\7�rm�	�B| 8l��pPQO��A�k�"^�;�l����)��]���smO�4l�pn�:��0Z3�vj�͌6���X9�K�.�jן�'\w��һ5��G).)Q��&��p��9�ލ��f^��8Zj
� (��[�^���2}>�]^�GS0%�H[җ&p�P<�����}�J��#<�ک�bq��5�K������S����&���,����`���0�˂2�}����b�q��0lQ�n8�I��K���Ψ�����p�VƦoߐHQӗJ5.�gE�+������Y�l�̉����P��քC�tI,*Vj�5�3�>��`���4����eP5$c�G��uZE��j��9�M�1���+�·��`��_�ŷ\�*�LcP�J��qU�+S���0kN~Ɓ��Θ�u�N�d��Q�������ķғ�wA��|�E	�a�Y�\f2yn����U�8��U>,m��H��W8^�8���}p�ш�l,�`���f�/�=��g���"�3֏�_�9R�-���"썾��\�/Zн���Ax��Nh��r�ƆF�k~"^�I|������	�{xA����c<	��Oױ��R������;�ߥ�(� t��3~G�����M!91+�Ə�
�~Ǜ�U��Q�_�C|\�Nc�ʀj'\έ`��9[E8�z݁ 	��[�3�2vqI�`�����A��Jƀ�
���ڝ`��X�J��j0�w,x�s�I�ؾ��N�Y|�o�z��x���$t_���eٴvbWs$����4q��Sp,����w�PVMc�+4Ck��5���k�O�Kpj-~�j���<*H8h�_�QR7�f��#V��ք|��$K�x?�Ϭ���Dk��#Z���� �EL�Y�� ��O�@��4�5���p8D�k�]��	>�OkM��3�r~��;�}�I���_�]��;�>�1`����A�KQ��5�H��I��&��`oBg����<���/�&�[�J&�'�	���;v-`4���_ P W��I�4��qf�(����^�7q�>]h�n�m�W:���S'���n�yW����:�������Q=�~uj�d�1��3�M~�>S����Hun[��B��o���ruƌ�_[�ki�������	I�=GWYOpD������Ǩ.2��
��L=�r󿨋^��W��YՑ�F��\@�3���3huE��a�[����]�2��'��33(L{);�J�,*��@�{���k�}��@Lg^]�Q�dJl8K��@y�����ƽp���_g�)8!F�PuXh�o�Z���Z��������8���l��Lm�P���Xa�|�5��<�A�V}�\$�����L���0��֦9�2��q�@����̥��RP�{��q����� ^�!-c|�K�E�D]���2uM�!����`�O1��]�E,Y�gm�Li�k_��W><�C�q�%�TuO�+������I4.��ӳ]�#)����E��T�2���g���@h��G��f6��A`-�M�0��wdUvTƽ�qp�Д�`��R{)-,���6��ثPB�8M�".�}���~�N���#w�F���G��$7���?,��eH��E��j6n����Ö�7��.ƪk��gM��,rڔB�AnŉUB�0�+���#��0��>�ڻ`�P�8V�h$�C�~�6q�i_%]Ϲ�I��'[Ԙ�'\�D��ȯ��e�IHI�T�z��5mrV9���N�sb��	F:����b�#���M=VB�O�연" ��?�����=䧜��ӹ�� K�+��f[��K9�$E@�XO���u.�ې�����+#׻|�I����{\q�|4:�c�l"Q��h:����G���4�a�r�y5G��}HS~�	��Ü�6��3�3�(�@ET#�����}D���3�$d�e)��9�
w�������t��<��C�D��QP�"�Ýu�{EBEK�F��珌�A�� <�rϣi5GWF�����������芔P����U�!uW��99|7:���Y�:~�J�TjT��Vm۾fTU�R|��)w�O���\p�p����:z'�5������0)�Y�3���ߞ�=�+�ޣ��W���v<?�CW��%������Hi0�!HR۾\#�O��^�2�.`����-��J��ul������$�(�5�Uݣ�O��5dCw���2�����#���L�A���㥣0��<�������z3܆"���{�.xgP=��Bx|I���"��
���ۯ�-��T�3~��j,�����aG2����\=�R}����p���~�eN��*
-b��_�cĂ��ȿL�xq?����h"�F��q�M�j|P B
*I��U��G��Z������L$/B��s{�C�# �#䩱��@Pֱ{{(����(�K�C�Ϭ�	��[PIZ�3-U�i8�ɋݢ��j�E-�T`%Vzܶ0����)7�	\@�����>^[�!�u
3I΃�Kc�mᖔ��D�v{p;o�J�Y�F�8@b��`��k1�\{q�{Vlm|I}�S��J�#�չp�F8���t����\�����5�\��C~v��Z}��Zl<���ؒI��������	����މ Oi���tp���������^� �A!�?����$Xxs���f�$���w�%�Xk����_�Z�XN7k���'_r�εƬ�3��3� Eҙ%���',�C�3�����K���:7��W�&\ �;���n�� D���FlF��g�Ӭʛ"�&Cj�&2RY���>	�G�?�˰�U�k<c��h���#ݻ��r��U�L(���%������C�2W�Jj��Vo;��\X�-
�sٷ<ަg]ܒ�Q	��2�P�.F$&)���6L�A��)
�����f_*r����H�4��3����٘|��6,]rSäϯc(��y����2)�L�Ț��6t�cw�3�uF6i�h0G���d^�ǁ�W���[���l���PW��Vף����Ӭ����{x�W��2����XR�H3Gv.��PI�����H�<K<������ ,q}����e�̞q(��D-V�ܬ��3! ��F1�&����i�%�&|�!a�q��x��v�z�%Co�n=J#�-<9c��6{��9BD�j�����<����N#�$E�^Auz��:���4�حU��4D%�����5�d
��lS�/����}����X*)5�~\A�	�)j0d��<�ml;;�����z�JęOGsyI��M����*e�cG<o��i4i�N�jy�͎��_&t�t}ATu�>_L���[9�R�7�U��C �I)[����XA�(�UI���� �lҔʈ/z�E�݀��ٷ����H˒3�����;[��7&Z�z�mL���m!��o�w?\Gt��/�E�f���Bo�'6RD���m|,�[���|����d��Suh��6��~<��}%7ʃRP�xt9��D���.Ǟg�U�Ա�5�}��(#_ŝ��EҼ�� Tj��2���ʬ���u�ωB�*���#d.qG9�{�Lk��Ӽ�h�0���%�_�"��n�'�u.�@���������D��p� ��c۠K�Tآ�7��~��UY�"J��^��k����H�0�g�����@���T��+�	�,�8�DuI��2^]M�h���d�S��ZU� ܣo4^&��Rx0Z�S+�2�ـߥ��W��_���V���L3�8#�t �/n��X?�Rf�o�;�lUg�z�P�ρ�Kվ��g�͡`�����g��� �{�Kj��(�]�5@�.�Wi[1]ڹ��S��ё�=��f?R;�擯q��Ns�NV-�;5:4�f�#����!��F�Dm"\�[0�Q�1�J���,_R�W�U�}7܆��[{S/^�C���Ĩ���0���$��Ԃ��5Q��+�K���t��=|.X@����-}�c�Svb�N|*�!|�e�qՙ6l��Ol����C}>��q�y�����(����uo!��_�`��m��T#Pq�aLln�k< /�O�2�{f�
`B�"�d���O!���ԓw�\�t�'���y�&ڴ�ߩ-�܍� �l6��xI��%�����(���\���"�1��2�����&M�R�#�N��~��>/�O��QB'4ƃ۟(`2	
�h�*����{�m�F8O������_�MV�t��*��c�ѣ�yc�K�=!�#�9 <�3�	�TL���.�A���[�m�����S���PL��	�χ�ʦ�p�5O+#�az�2�VG�'��u"�EP8�ޖ�^�	�?�3�d7`p��'G��l��/��!�z>6��
"��>|� �9���N$X��:Fz�A����U�ؿZ�%��3�`![+��m�?����)m ��#3��0uh��˧�'y�s�W	���e�l��O��*�E�az�]țẜ������C��u��	�A�^C�dɟ����c*���ɪ>$N��G'�I�d^�����/dY#}�)`����x�"W�!��q�;�����AL@�K0׈�C�b�}��<�߄u�@�8F��C*����v?C}��l��DIʒU��#���Ȋ�0���,8��-}ʆ����%w�è��̰5l�J@�58D)��v�G+9�+��X�.��`�@xm���W��?���[��t�L�G���4!�,�v��z���N���2���<X��	�q���i�@G�����B`�s�d�f?鼸�t�_#<�ܴ=�;uڭw� Y[*�<e�lU@�����l�ٗy��d��l�M��}�*�[���������!j�̿cr����N
�-}>~lg-_��n飝�͊���;Zw��Q[�Ae�g�'.+G~U�0�?Z���Y6�����sTW���%�W͵��#�p!�Н���wm;とbn�&k��Ij5>�4��4X7]�l��R��ܭ�Z:ν�w���~�j5pt��$ʝ��o����0�3��˿-޹�����Hf���d��������L= � ��y@<*�lJ��C�g�a�v�(7ĝ{^\�b��%mu}'z���d�s�N��IQI���*@�3�L5^����Z���M��m��S�/
���ĝ�����lS
S��K�7��&���� �I7�ͽm���
:�)�KobV��N5G�<���x���aBW�d\˅�bÄ� �b-���Mc�7�	�C�D�ڽ(n�)�٬����8|ϔ� ΁�G�K�n���{�Y�1�����
�P7�u2-ݠe�k���l�S2|�K�6�����ICQ�h�^��[�*��(�S3�o'0�V@����xp)\�kw/�����j �Csa�8#7%F5�MK�툑y�����g{�*Q4[�f>Z�׈���%�  �_ˎ���
�@ݨ_E�IY�S��Ka��N�����C�6��_
��E�`7��Zb}50D/#kB ɱn"D����T�a����euv^���mI�!
 z`���=��d��JQ�H?:��r�J���1�T�S�G�!y��o��"��Q��W�geW��A\��9����0r%�XKC�m���P����������&�[��P�UF�3݅A�����Gd�V�1!݃��&[4���2HQ��Ґ�{~�E�eъ�8�s�|�ѐ6p+�L#8��� n����whP'<9�����Fz�����hM�L����0���8���>wG,=a �`�fY������̱)$
3��l��ݖ'�������������<�E�o�p%r�T-G�{���r����TI�%\�C2���5�n�JF�L*\��AS�cV�g**���h�V� ��7�vC�#�|$�:����#g�����"�X1X-�X�r/�d��M�T�I�gB�-�Fz�%W�X����z(�9�3*��mk*�[3}۲m<��)P����|��9�v�;	���p�<����\(� �gq{���T�$�
U�*04bSEH�d�3C�,��LTED���{�nxe<���m�s冞�0ÿ�f}v��e�$lf�Š�h*D�5l~�c����=����5]�v��dg�W��bj-�֠� X9��6� �Ku��/K�� (����L/�h��S�2��`��Nr�0R�:���n����m�:·]�*%���f)��/WҕQj���r���vV ��,��>/o��5�=�&Q^`ێPk�y(%C���o4e�FtU��_b�N�G1��T��;c�+���U_����6u�$�~7@W��ڔ� s�̾We�ȆX�@y<e�٪]͝vX|u^>-ZR�K�F��(�����F�$okMG���aJ[�T	-bzi 7�f��@�Ün�������F�g��뽬��
�DkB��4d�ȅ�%�/]��'d]�=Q*t���"�	��&FC�j�|���E�K�&x{$�W�[=�C�`����b?&:@s��9g�ֻ��%����J�@V�h�s	�4e�����,�D1��VR�xr�~9^�i��L:�X�-��� ��b2:@����JQ��o_�{$~���R�M��L$����Yf�I�Z�-+���g,[I�"�Ӡ'  �n��"B;�;-�ˠ�v��FfA�'£YL�����ݢͼ�$*�1a�$�w��-����
�����ZJ�Z�;��?���p�C�JU͝���A����^-��"S�<��`�[,�\����P¿o
&����ӗ��Q��^o�D�r9'����S�<�!�+�������!Ct���He��g�B-��6D2����;�G+���p9��w��G��Ֆ��Qc�<���F=��7���?_{�F�;@̺	�O���{�Z�~�!L�I�X�4�8�Oh�ޕ�ט��I^-���Ċ��0�a��"��L2Dz17mq;�Yv:�,�~NNN��,�*�� c3�^t�"@N?@�i'b��Ӓ�*�٢X���~��x�
��n3�*f%��@��?�>��jþ��X�g\���2�5h�M�d��ˌ����N4�c�7tl�e�^�"�cq�L���I�n�����ޘ-�hI�q�ȷܪq2�ZC�.ԃh�, f�\�h����{<�
���	�#�ٕ�1�g�rKZ�^K�3ox���ǔa/��ߘJ�0yua6$0�Y�hp�� ��7�e��_N��*��-�#q�+����n�tM�j�iX��(0X�p�WS~���l��c�F[�"'(N�l�C�W�~|QWyE�Ĝ�XA�w/�%�
=r�̷D/��ѵX�{���9� ��b���Չ;d5���5�^��T�A��Gh:��N�r˶�-���p�	^I��^�a�E�Z�i�Z�5�Q�҆�X,.�"�3q;���
[y���9��Z���m}�ǪE})Iz�Ks�,=L͐L|��ג��u&mE�����'�;�2x<G�����kÃ���D�cE���IX�R.
O��n5���t�7?�v���$���(�P�&6�S���o��#u�ކ�����i�I)H��A��Q6��cIU�^��tR|SE�����&Rǲ;x_���&��;(�.{��0��1���Z�Û���۱�N~C���Ȯ���d���?�ϔ���AU����Q�M$=P�53�qF��V����	ۦ���&�^���-e9؄��F����Zٺ��z����٢ ��(8�M�D���;얺�tu7�9�c��d\g�I��a�DYJ���fp<������8���qQ���=*��{��t+$p1�b��!�9�v��1����j�2�2�>g��ʎ��	_�7�a`��1�Y:�0����/�3�AA�C�5�՗����/-�K%�P�>��zyM�Nʽ�]v�T�pv��ˎA}����i�Sh�rA	�3�[�m���3"�#�B�w��H����_���։~NI��37��X�S�ux��nRV.϶�X���)�αf:[m�(������DR����]�G9�5zK��xr1*'�!E�7��ςk�<,��Z�L�͕� '^���%=re{�(��m���K�W ��U���W�6�ʹ��m��ft'0�����f:�����n��Ӛ%����+ۦrt�`���$��6T���s��B��VF$;�u�D��@��V�b?��$�d�O�;�^[���PW.�sc���cn`i ڱ-#�Y��H��#�j$��6T\����;p��ۨ��nX��6���K�j��w�����H�	��ΰ]�^ W�U���������d{1S<oq.��2�|b'��mS�l�ǉ���]�M��ߞB�	*^���KF�%�2��6"p$�)LT�g���U��ޓ�)Rj�%E)� �u��﷥���m�(;�뼎��wc�}u�Ċ;�G�@8�P?��ޞ<	�<8�g_�0��(�s�nOL��Mgq�C4��w���9o7�}Z�C��)s+��:��#��;��b1T.q(Δ�9�L�b�C:��b83��iU����0��,���X��a��	�Y�1�)O�j����D6Z��6�6��C%�1��l���D����)i+�#b�E7��5�`��Ą݄w����||$ޟ�w�v�����>O�ޮ���r�9T�4P���²�Tm�tm��W�]5���}��=�h�}���]�!8�[��±$�E$��b�\pSh�D��Y�ԗ�H��ռ����q�j.�T���t�A5�Г�j�Ug� 	]��5���N�Ѽt���ږ�Ŭi`��[KY������Ow �@zBC��Q�ΉxuB4;C7Uئo`�9���Bo�}#v%���dzӑ~�D纇�X�]r��Y��>d4Y�u>�GO���f9�>5(@�;Y��匚H#)Z� (���8b�_���F+`������)�@�mıM17aY{�*)�N�y��v ��8���Z��]DY#6&Et�7�`RMZ`6�E���ϛ�oer�"��bQ�Z��]�^pC��9�4S�O��jV֫k��װi�:��<�p|ϯ�1}�p�N�˯0�� /Kj��d��E�>���T#�א���C ���]��ίp���0z_*�� �1��9О�+�"��ӝ�|����p����M���;�y�ΉI��b�kU�an�)��.�$�C������{A�I#�T��tB����t����5!4;`a��fze��{��x1el����K�R���4#/���1U�+�n���;~NH�BY��(����|+��j�;Y�CB�5�b��~�J��
|c�H���|�%e���u�qt~��L
�A�|0÷m����"D�A �oU�#U>�s���^��<��L�����*k�[��U���ĝ��7��Uz�D�A��*1���K��,b�Xg_z��+���j�j���ߖEGti��=����`��pЖ��Ps��҈)�/FM�b�G~wWu������QV�VL��b�-"t�6T�v���J��D�2"SaZ��|��U���j�*��U5pH5�XU�²�O~�.F���L�h�b���α��H�� Q�CQ?��Z�;9@ E��e�u2Qq��,xea1��D/�r���K��K��z�<��]����T:�#i}��"E��9�'�Uv�8WBcV~w!u��aΏO�Uw�n��?��O�����������3�h!�@,N���,�W����tr�C#��J��Rop6�Ө&��5��o���% ��9�����i�#l������2{��Ul���z������Q+���m\1 �=�FSH����A�IF�0��Tٜ�.���)$䢤��69�� �a�h���T�%T-�����v5�Cgm)o�-��_�l6\CD6��5<D���_����<�/��WX�����2���=3GI��{!X
͡��o�1ӿ�eb��jv��{������)|�-��-�`e���4��Y	���c�B$�t�AJaV�~� Fi��N+�������L���򦷃�qo�jR�@�:Y����Wgm�oy���$��>-���~�x&�_-�$U&�LEJIZ�CqZ���g�g����6r9��T�i����}���~!5V
(��-���ގQ$3*���R�!6o���b�|~��dHhn%r�V0�V�h��BTe�޵�ۥ��^�W��-2�$�q|������<ĚN25�N��D.߀���W�UyB��K]��,�~ i4j��o}3<4l�ʋ�����R���1'2�����.��*:7);G*4�x`	�Y���}~<����k�(b��!V�vE�Đp�x\�+jc�f$���M"̒#��(�7T�ж��<(N�u��rWW� #�E9�K"(��TF���?�T�پڟH_�7��@�m�Ԉ(�6/�oԦ�4ӛ/7P��~E�������x}K�m�G����8�:��hሙK�s�4��R����Lsx�Q�귊��h`�wxq�YuG�Stq�wì@�@�X�y�s}�������.�]s*������Ɔ���>���fߝ~����2��Y����:��?ޞ�"׵$�Ά�����dkC�\�o�R���;��^���E������<��mk�Õ�Yߕ�Ɋ�I���^߇Z'��=�j_��2������H�y*���L��M)�q�At�����[vo�71o�\K�98� ��a���jL���|�̬2IOy4�Qy�>P��7��
�����c%��L�j��`�j�kJuk���I�R�t�*u�晞I�Θfה~���Pܮ�7�\�QB���s�v�Ipj�t�'2�_䗵gQ������[E����$�r�+d��E��Q��7�Frr���J�~��B�Ԙ�5�ǣ�-y���8���8��6�߅�	��V���/,���|�!,�0~:��M^ۣc1��j��BH���5��!y������3�j���V=����W�uzڭz	��=���
�� 9n�!э�q�T�SΤهg����4�n2P�Ab�wn)��W-�PP� &�ݨ���R9�u��uR�}�'�a=t�۩���9�֑{��;<�D ����|@��q"�8��0�3��i�;�ಲ(t(�)�����"�?����Xq��%�^w�U~�D-]�S8��uR�:�r�?޵��N-�դ�z�Z!,\�}@�b�O?�=�B=	Qu����(�2��,%/%��V�"�Q�ޢ�'ԎK��hZ��A�0��:�9��%�f���](F���m���E'YA���~g�	iNl�`A��Ͽ;� K�xx�v�@��\#�U[0N�ص�ޝ���v=K
?֩��z�m��	5����������<!�� <j�m�/���:f^-*Q	�g�n$rC�w������3jLg��CܝqG]^�O�ٰ�P��Y?�"T<氃q��7�e����� #36K�Fi
mq٧rd�5��� ����UtӳI�
��:aj����6p��&���`��bF�z���������#�>J �8�rl�,�	Id��"�����'}I�,bop���~Mt���C��d�m����Ψp�!&/>�q�=t�`�f�L��|N'&4�}��>�3��C;H�\�#�r3����}6T~&i*�Z_3E��{��uwxo���
��
���	�)� `�Y��$����������CPO��C�/�xݙ���ry�G�x0���*�Y�G3�Ӷ�0�]�䏌�	z�58L���W���h_��Va�Z��5��
{rs��nw��J� �[��k��c�dʚmӧT<��xr�6QYV�a.LS+1�W�s:�#-���g8ugB����E��:�»�����FEC9�w��$9( �0'���u��
zM	8����8 �]����������$�Y^ܷv�Д
@�)Ap�$Xq�"�@CSj��n�3���o�8�wi������6l�!��.�б����:�5_��萊��oO����*��ߣ�����}�IE��gJ4��T���Pqdf�c�db��U|qQS�k`�;&�0�-��=va�-�MV�J~Hz���E1N�$�$��.N���v��9[�3��m�KFGm�"1�"����7	IV�J��c�g�[h�c�O�{�1����h�>/N	m��s�.'�r���l���s�$t�uwjQ`�3H���7m�D�x{�I^ӛ�Pz��������*Tk~=Y1}HdY�����Mg�q���43v=5v-� ط��u���W�f�b�fV(�����T���ޕ����%�WE�[���%1]&�����=�}�V������ ����<��7��15��M�]|�,a��������V�c)����A����bq�i�9e��<
��1}��9�hx�FίX������C��F���d��}A��C l��G+���.ܔ��2p$�������t��y�{��X���%�i��!Y��֛l�8��0b�'�y��RLY��9*��O.�J��/s��
L���r��ZGW_����n���0UA��?Rrfv�������R�!�!�2��ɽj��U�q�ZN�l��$J�]��>��)���Dϕ������-x"3��i���i)�eO�����Zy�]2~[���7���3���D��� i����THa����J���$�`㶃F�ʣ��S�<Z��K��O9r��@p<�Oc<��R	,�f:ڙY;�^�u+�C�e�k��-�5|+�6#A����█�Kl��o��u��f&碯���v��_�V61���v$��r�����.,؜�Ї����"��u4���j�S��RT�����4���<�̍`���/재�I'�k2�l��= �${uu�(�dVzx��x�ʺ��1��/��������`O��xaV��ĦX�|�8KNx�L��9{ʡ�+�2�q<�w��r�(`�6���q�(M©Yu�-է�I��;Ԅ��Q�?#��,O�����E�|s�*��'H(��;yMg"���=�v���;���X��iF���ϗ��5��ם�M���p�w�1�(q`�z�>KL��]LQ*3�ƌTV�}U���9�� z�-���U��A�C�nm�oh7T��g(���CWeq�ѝXXݐ>j�_h:��)�~�C_�$�����R���d�M�2}o�(�|q������r�NēFP!��t`	���I4 4-��]SK�w���O�rjM@$�|v'%r�{�q��aK̟O�¢�@����MuW���,�5"��}��@��;B��'�B��x��2�~D����sqC��8�]��/�[���$��ABi�������1 �$!��v�h3[s����	&xR䜪��uh,�`�<���.��_D�:4n��nnlL$	9�ƶ�	I�p�
���xmQ�C�mi�R�1�.s���v��aQ%�s�+��d�)Ą��=>�J��<h��Q� �z0L3�N� wP)l<swC�������q��	�����5DW�9	xtyM��wU��:zMB�_$����+�^d%.�]�q��@mu����cq����הK�ԫK:��j��7Py��3��;�W�!���:��0��qn`��&P�{�5�?����>�gOê�I��	4'�,�t�G��BA���]�B��x����1Մl���`��O��?�u�ʐ}��t��Y�TD�|�g2����� �Ψ�8о��ɼ+W�>|����Q��U��0Lxu�4[��F�%P"0�R�b�������O���'��HfF�B��+��X�|� ��h�O��0����E����[ ��!.?��Y\#mC�rh�m���K��8~<��BH�'X5a=<��2�V��d���,���"��	����#O����L����Fl��ɔ�ɷ�gj���s�1�&.H�����"���ѷTɂ^��u��������|��A�%Hד�����?v(gx^�N��F��b�nA�A?���n�l�@I=we�އ�O��R�lk����~�9�3tNu8�<mw4ı3/�3K�����j#�>��4��R��T��6^��ػ��˼�_%+C/=5F�s䉿����U�Xi4.�-$�V��%rUR����f�$���- w;	U���;�&�M�g�B:�w�$��*�F��i�^
��u	���5�ӢØl3���9r�6\\��|z��О>*��t��gO�Ƌ0�އ���r	[v��u\)����5Ɣ�M�!lFV��o�{�2�6�n������Ŝf�c
e�����p���s�M�خ���R�4!��ɰ#��JqU2ʵ�BÍ�'�h�����),_���� #���{j{��?��	F��2��1d�%*=(K�:q�+NѨ����h��_'�yJGn�JV�{�+����B��8}���+N�V܍�ư��~�,Y:�+�|��Cy�/i��䫀"l��'?Ȗ��
�ԩ#4��@Ki��P\E,��I��m�jǖ�����dbk�;3����B*n`}���N�֍P� E��6GS칬؂ȍ�9aL�� �NA<���!"��P���lε��~
nO��2y��� jG�/�N��;(ˀ�$�	�u���T�u��ʕ����?!���������k�pM��<�`y2;_ز�,І�y^�?,�z��Բv�q1+ˀ�w����v��FWEVL4�&�nYM�`�2sN7u�ֶ��|�� 	�de\:Ͻ`Jʣ/��
����_ɇ�~�]:M��G4�{g���{��9���Й2�[z?P^�1�Y�1�y,L[��M�� �5uB�	�I^@ŧ�=�4:��"獷�ř3rdG�w
aͦ��$g�u��
C`f$HC���T����f�U	
�E+}	7�C��Ndj}�x��ʾ%�Ss�A��f�^��h'~N�z�O	#�+���q<Iou�^X�~�����Q�ㇸ��C0�=:K�}a�z��$D]�r@�.$Ǽ@!cg�p��3E�Wޗ��y�؛�s�Ha�b����\X<�@����q�����ף�D��[b�`��Z^�88���8"�t]�w�|�17f��'�u�+<�![�VTB��xi��Ƌ���������_�_�g��
Y���p�����A�%�5����=�;,	�V�ۙ�G<T���~F�;s�`�n�}�Qj�.��*Q|�+(���?���O%��1YWC��cEI&q���A D�VVVu�ǯr��v��OE�v�x�0S$	�P��D�2��=b#�D��w�'�4:����Z����
�D� �83�] >S�=j{���������r��x�(��۶𾺫��
�zX�����b�E����SK��pt�#�Ks����1����S�/|��+���k�h^ 7(�4���]���	�A�xt���#s����H �	14ܙ���}V�f�)>&�F���^yg�D���Q�#_n�ӵ�?���f�X6�����!4��0b�/��~|Ѥ𴳬VҜ�N�əX�ܤ�K9Do�"U��v����
3�W��6Q2wS�i����&���:�3�ܜZ¹�#����[���]Y�v�$�,#�j�?lTg�¶��ю�f���p=D�)1�=}>�R��pq� ��j[����`z�t����lsRx�5�`ETC-��K��)7CL{6��y���<��7h2cC�	�d�d����� s�w�OFC�W�L�s�+�Hqי8��n��y��I�^���z�d�ŪB���K����Ꮔ��G�&}\���f~ u�n�0�^�&�h,J�A�m�,넷��`���[��6W�4P�D7�Lx�Li��V�ncc��O��朧�z��s^�溽�Qi��n�Q�V)�˜q�g�w�J|�B1��Egnp�-r�U��L{���e�o��
����0�|�Z�z|�3�l����Sϙ��b�� �90h/���ho��,���������oܲ��̇<>m1�@�5�����A�E��JA8��|�Zp�rI@��Z)Z1�����	�#�ztS�p�kH�Τ/��G۲~�5]���`�[�ee�<W��d�*!������KY��=ѓ��p��m�ři
Hh����=���R�t"�'��-��j�b'9D����H��U�Ķ"m�ôI��i�nR.=�7@��r��A*��L���M�v�42�9ph�G3{F����T
'Z������m�D�1� W�_W���~�������n��Q��y�3���ͥ,p�鸅0�Z͖��T������@E
�l�	�]����;N\̻tE%S����e3M.6��?@j�;0���M��z��y�
,jҎp�:}r���E�gĉq�n�;L�CH�7��"zyu8jN{�	��5�s$6��E�j�)ȯ����I(!��i����o�y��zt�T�y|%_�A}9�}�V��R�� �
�O)F�֘.쨕7����~����*�BN�β��]�Pzq��vBBTZA���'^�@�B_,�r�!Y�d�u�t�LF/_��T��T-Bf�Ms�I-��2�i�b��ҧ����I��D	��`d���R(%K�j�F�^v�it��(��`�E5��5�aȦ0J�j���ӂ�[�3J ��k��vƓJGukߡ5�/1���՗���n���=���f�/���@�;�2O"���y��A�]�@P%�1�&��2�ʴ0PGSܘXH߶VO�5��{�II%�\�-y�\���K$��W������5�)	dx���i�{�'�G���x-��(�nt���:�KGb�/	v��,K>��-f��]k4'���+s��O�*;e�vEp'9�y
�t ^���B/^�p�����V�}6)��Ok�i����qh�����=�	_�l��nhBڙu�8,�����k��K�p�Z4�`V%����Hܙ�-�#����P�($�Vh3?�ʭ���p���8����#��p_�d_�|�t����I�:��3fF����K�n�WS����'��'�,��$����T�`s+�1�	Y��R�ęQE�?�
"j2���UG31��gD��1�E5SA&I�2(�ljc%?�jlr��XB# �6�����d�����͉P�B��qV����w0��d�W�ya��"��B:y�,�R��X@O�d�\��ppչ�n9��|D���:�Q���\��Y�r{�p���(�{r-}H�z.UtK�^�O`C�17�����Jwb.�.*Y>v��`%N��D{�}�Vk���#e��	)���.N�������3���ǹ����蕣]�~3�ҋLxX&����Y�ժ�`L
�F���h\�FS[�	wD%E,��?���3���}a~�!q��`ȩ�6���Ȧ9��«�%M��(��"�{Ú#ʢ�Y��ŽfP�MEűo8;?�!t��FM�N�;=��Q��1B�ލ;��y����T��I�H��V�@�m?y����^b�.��W8��z�G>E�`��L�"���O���d�A�׹���U��)Ք���3�����䞤f���4yݷ���cNl�M�
�y�Ip	�4:���ďM�����\[����_𙵁�Q��'y���Qh�˝D/�7�(6K	��X��o��M��\%���zV����_Le�m~,j��s)��=`'=���<|Ar�9�Lq�tlg�s�K��S���"���u�%��nH�bV0oQ�&E3m�|���qB",�3)�C��k�'>�mk�C���Ԏ|%z�	����cp,6�R�c���ǋL$�W��>�[���V�wU�W�M�<�xD'	��j���c`������V�㉙�3�La,ᣃ�tC-���,mQ�F+�D:�h��n�Q6;�U2�x�\�-f���-�Q�v��S��B-�F��f�v�I��$E��p��HxG�jY����e�;^U(Y�]o�/�%l�#uEo��'�-88iށ'݊7ی�s���X
��팒ؔ�'��9�|��{*����L;ֱ�ґ�j�5K"B�r�ߜ�:�,��y�ˮe���^ �pH���yZ�ӡYn�19LY,��ώ�T~Z����mZ]��3�)�S`&P��WO����ms��bQY��ȶ��U �{�p���#��;��ᚓi���4�!��El޷�/Cet@K�R��o^��aW����&Ż1i������f����+����"�!�lki�����Ϩ����Y�f����
���Z��?D���[�M�zKd䯞ɋ}F�oN�}kK&�l��o���80�-�7��v��z?G��i�U�iԙr�餝H1��ǀ��zx�"x� 	e<��N1L���_ҳf����^Z���!���}�{�I���L��IW��	p�vOF�|H&�Nr�~��������®���B�>s�S���O�Mj�CrgYٺ+Bڨo��#�o��o�g.�;��N�-enPn��0�4�^��ļ�N��`Yc}]c��|��9Z�r��]`_�۟��)̩�7k6t��f��z����-�m�M,.�2kg�ʼd$��o�?̼���U�(�^h`$�\\u�?�[��L����[H�
�C�CS1�[wL�=�3iA=��F��0�U���+A�#y>\��L�x%}*�N)���XM�aE�g쒀PD�G����]�G<��<�i)ri0��"|Q�?MW�\��0N���A(K፛k-#��9E��9�KV��+l�����E.P��m@�/���qZ�f�]�e�'{DP����1?g�J�Q)�'>�Y�$���.S�*}�g�~}V����>��49��|X��r *��ʌ^��Y܍���aMK.ti�
��:X���<mJ��D�A���R����Ӳ�̆���bS�KM�΁�b+��|��4%����<��q��7"2�g�Q�b7b��ࣂ��A�`���\�+FN�2��O"�ޡ�nZ�h5��H��������>�2��_�5�yp�mʢ��A��]�G�_��:�W�̰�<%��kKGyr����kR:���)���N����f�L(z#���c�L�VA�buCY��fG�b�������A^����r'2�ߛ%]�M��gC����ݺ&��j����(�͹׮��9G)~l+Ǟnq�b�ה����.�
�4~}G¿����Z���?t �Ma³��P3I3��^|���`�?H��X�&���s#�;guȠ�%|����/�������m����CV�&HIx�c0y]X}�ޜ-�J���`c�F�R'B~q����?���W �R�� ��1���L�u����*�/�xV���16jL����Ȓe9�d�a�@�ߏ>��ˋ&�pk�	�qJ ��"%��:j�!�W�nHyC_�7X�4rʳX$"nsI�����o��(y��y}�����$�ο���(��i�y)��e^~�f����p�ޅ	�S� L�g'�#1u��2�kD��b:�u6�{9��ߎ�xB��R�:!Y�%�ȒPT���`#�m�*����Q�4U�E��5@�ǚ09��Q-�4$���-�K8~֩���f^�z�5����e�ɎR^t�)3������?i�����"�YLM�|���wԘQ�h�0�r}��L:��dn_;��9�M���m�-xh�
Q3������͘�G@-cH_��┌M$�M�T1�m\]9y��=�0��Ȓ,��n��(X3-��ix���@ɀ��o���7�@�MV�+m���a��H��P��~��gN%x����?�\���tT]o��DIDL���i�ڢ�hn?���|r��ʱ����Ðŗ���:3�'��!��O��Ѷ�x��.���{r�C�h��w.3�*��Jb���A`ߟ��
�)'}�q&'x�j�őO#C�(�Ee(�&t��=�!�-������u������n����(Ѡ{�l�:"ޕ��Sf&���"�}�62TN�a��$J��z\��w�69)NΤ@~#��f�p��g�b�����Vv�d�Z���@�e���	S�iX���EңA��Sž����NPr7�^�@�(�R Pd�m ����e��RN0��,^G���L��o�%6Ū��P3�t�M�-���&���S�}协��	�w�q��w���}.�K�g臾p+*�}<UCK��Y�׽j�j�8�+��Q'�^�<s�BE����,�]Hi�'��H��8m�{��p̉�|OHr�������ԃ���n5�1�����wP.z0H/T4�=���ً�eP�su��Ey�ݯD
�8��e�f�鋝�#�ߒBk���o�mN�.�b+��~;.
:�ƠM8|�3�ż M ������UA��J���>ny�02���zG\eU��yУ|���;�	a����DbD���ܠ�u |�Go(>����s�CY�ya���Q���;A	p�GQY���9M��o���H��Y��l*���V��?��W�|QxЁ�4�qs�o�;��zb}�!�$4X��� �e"bv-�	�e�Vm+B���0탽�#~�A&�j�r\�_����!����t|{�ԧ�it�`I�G��L�
`_�H+�(=#a��^E�'��>h�&��%ucb��䏥�^�e��O� ��-�婨�./N~� �Dq%O��0Q �~*����%d��D���-Ҡ���!'�ԏ�8�_"�j�,�Ҁo�7|%�o��p��H3_ba����,�K�W��Q��Β�1��g���GCL5%'Z���,D"�AƅYi�hig����\���KV�8+��A�"#��7�n��i�(�F�|3�o�m���ܣ)��_��Wٲ@�'x�K�B����y_�:���9Ɉ;h}���!���mC��h�DX��fH��VS�b�{<�����fjC�m�֔\n���J.5�2@��I�%da�t��-���3ϧ)<Ey���!E��7�̾q}�IKs�9S~�w�� KG8�C�`�TU�y��2�!Nx�1� PA��6�R�F�^��͘>���>�Q�˅�	\9�i'��W`�^�@�4ug�`Cс��*�e�Q>���u�uk��4��L���n��$l޽fY���ʜ*�]��#�Lh[�d�W��	�j<��8 \<�wU�zB��d��L����7�a�Y.Xn�'��b)��p@r=s;�3��w�h�k��;;c���AێA;s�>�@"n���Lu23���UU����NR3�}��۞~�B3�L�+���/c'P�%Ky�9�
����v�z�<okjG���Ȃ��.�vRo9�2� י�h6ۛ}h���i��{�Cv�����w��ޑ�_����݈�t��ZPP���4�N�x��Q���8�'G�2�F����G���� �V� Z��Ԋ�fn��v.�@��`�����쬙ZS_��R8����,��YF��Ʉ��?��#�}���8֘�!�t� 
�zA���Y8��&|�2��|j���Ns�L���p�l�(fC��΅��;4Fj:P_��"�w���]����Q=	�7�&�ߚt|�����\S$%��G ���{~z!��]W�ey���J�ٷ�}5!�c@ŭ�X�j�˹�X ן6�.4��W�ukfP%�D�&,/sn9}F�yV^�kulnPevjAl*�sC��G���c�E�o�8�����ga���]o<E�J+��E�����.����Z����{��8���+u[:����AfR�2[=�۸M��\`��\�YT�]-\��?�t8q뮱�pxHv�L}*+fMEI)X-�픘��+w�w�敗��Q*��<s7�.�1/��C��aI�([��?r��E�?_�.�5�U߰�x0�K,��%�&s�o^Sd�T�·�W��#��S�U��Qg��Xgnm�j�K@���k���zQ\ܻ��R�4��E���_o�Jp�+����*����%�fU�4��_E�[1Q�Wa�4�zCҪ{~��T�a7�-j�c=S᥮B�P�'�Y6�e�b��]�If�E�?��6����RVÊd�ފ;d���qS�\�pG���n�D*= �q���G�Xp��U��t���}�Z)|̈81���nYiHR�R�	�`�b�P;�Ӊ�M�MEYm�Vyf9q\x3���ެS=L�������'��̂���&�{����QN%�Z k�OL�A��Ʋ>���t�?��!P�)v��bM��_@i>%9 �Q�˥�I�Z7qX=q0�����-������"W^�Db�a~���ӧ��n�C��K�6hfK،Cx��<�p��kũN9���4s�F�S�gU����͗�n�1)&>+cS8���z���E�xG_gj�o�v�Eo��rY�W��6��Ga��D�k�ȱW=j�G��j���icҘg�]��h���Ej���l�����dߟ�[������L�ɥ跤vk,���	�hC�ę����d�n1\)oT�Q��!��a���3�K�b~!�9_+nݜ^J� �����٢��������y��u�X�s��x���~_��YURbhm�5p�sN�6�f�HC��h��ڮ^)X+j�i�-ta�� �5�V~�Yd�����az?|Ns��@���6�9����&�)ZoW�9���d_�L�9F�������3���C .i�4y:{L�%\�dwo%‑����(`�Į�Ih, ������nPO���L_���s��������qi��*2����	�D�q�80h?׹j�&ưR��Q��~,��o#va�Q�«�[��H�}fC�#-}śx�6�E���?]��_ɪ#�A@�ߴSt���RMn,m�Q�R(�a�u��s�ý!���ч��zr\�ӥg�[�*���i��'�Y��{�W��9Z����줥��M~h$�#R�i(L_*�C֜X@`Yr���0{�u�r?�[c�q�h�L���_�eD���*���?��,�7n��Č�S�����n�w�g&>=���L�qͬ��D����\֚�o�)I�ST��&�Y0�Ҩ⻱xpy?�oMݲ��1 �]n�u�,Hжf���G��榆�Sk&p}i�y�\Եw�^����?�w���C��"p+߻���S��#����Y�-R?;�3���~��\�!g�_rt��q3��JjW@�6(9H�5L冀�x�Uޫk��^���'W��rfSw����8ov�&��0_3¢~T���h��OXP�Yt�fϑ;�x8gX����)5�I�'O-y�S����<w�r�� ��nm��k������J��n GU8�@�Ƚٙ���GZ��@{s�G����t|5�S��B{�����HL�ЗhZ@�XU���Py�Q�z��zq	�QAb��7I��_��E�� 3Pغ��f�[�-�qA8a�R2,2Z�F����c�$���;��/���GO���l7f�?�hp��L�Y{���+�hè��ă��:6�|�ܲY�z�1\�"+w
��nۤ�!�d��BJ\��!�W`YW��)���9�4*��A��T����8�6�Y���1��_X]����j��Nm��b��|*C��+� k�-I#��N8�78��n��.^�;d��"9�A�x-U��s���H�钵����m{�k	��7.{�~����T��$�������_|�4�*�K9A0��?�^�".B�0H��,P����s�jL��f ��Fo�h5���녈�t���������=؀!��A��������Ly��ʲ���v���@°5�!i=�h�	��&�4��}G5/'3PUΩ=pI%�*u��vu��Fj 7����1v�$�I��a�r�M�����iB�	�~L]Z&5�ڎ\㶟���;�5��Mֵ�ϋ�'d������{����4ǃ�Rֹ3x�-���� 4�[�,��g�~�і�\�l^��"+�Meӯ�&�VW+i.�w>j ����s�L�!o��m����ip����&�B�Z`�8�U������[
���x����Pr��	e^��N�n��� \D�=T�zp}^��j%Z�ϤP��@ov,L��3�V�'W�e5�#Eι�f���!�:|;ǌ��[ ^�XK����F2L_<��;�NK���.��4��+#��`�(�|��k8�X�JPo��S1��T�Z:�7/�0[p�X���3��Ļ����̚R����Q�����#7Ȧ1FA=Ƅ�0RrM6��_�8,��n�9�2����;��wDd�9��nX
�-�֖Ǝ��j��*k�%�\���1��7m�;�4��	Bz��wş�����! k=0����L�8U0�e1���W���� F�\F�3l��h5Ӌ(U�y�92��3ۏq�%?��(6�_BH,�t��9�>�-?�J<�nM9\g",W^�����D�H_�|m�׬�W�|��?���f90B�x>&��9�h�!4��_�!�;k�4�\ߵ���z����`Jͻ1��y��5�-_C��f��7@�H�2��/��r���?H`�s`���O�b{>o���j=��!4������=�b(���J�Bti��`ax�T�;�$�	����u!��G�r�|�B���zn1�M?�����n��_c�0���)�q�= 5�ژ����>O��=UL�����~���	��K
~�R}j!(�A��	�^�9n"�x�A<��72�ߊ���LR�:����x���#S�қp
�Ec
 ����Jʘ�y�՝s#���,�M�f0��ϡ;3�����Q��Z5�K-�T�!s$��/�W�џ���w��rV�j�v� �8��	������\[�V�d�k���{��&|��Ka��#��ـT�v���z$/�����6�;��3�|�h��
���I���K���״\�� ��Y����=����݉�#ިbzq��U�@��k����!!��(Z��P$�\�9�t8�pKS�@ =���T7�
�#���Mᕮk���� ��X�*+5N�kݰ%��Ѫ�yx`������p5�	pQ��-nhr�L_jG����h|��	ԝ:<+r�8h`���^
�	[������766�����|�R��r�YFc���9/�t%��k�a���Y�z����C���-?���uE?+��Z\R"��U�ɾ�r��z���8(��~�Ao��q��T�(�i9�¬^i�=?��V�4C�XM�kJgͭ"6�Z���Z?���!l�
� �(5�S��B&�e__��ױ!����*7>��_���>Xcz �"�B���w��9�P���C9� n�q1�i����6:���$��xh��=��s���΂�u_�+��Vp��L� ,�j�4�
�[��?E_�����c/��p㬞���-I�&UPJ6E�l��q�ސ��f)���2��y�s� ���|�8ɏ4Ͼ�%p������ԣq��ѪNv�s�����������YI���`�&8�y,Z���	�2��O>]k�/�f��:��'��AW8����Xs����)�.�r�އ�X�Y��)y*p'kUc�ˀ0���+��+���W9C\�xs?����������q��@gJ�l�|��=�<�{������Pķ�(�	��;u�_���r�3�+s�1�u����t�L������ؓ�`�M�8~ʌq�����Q]I��=E��!����O�z�%T��쓼+��%�����cqE%(a�(�#\79]��͑�����/m�r:��w$��S�I��5w�/����e[�������h��h؋�{��0��%Fň$���z��&T$u�@���{����pدId��vk����wV��o���mR�&��Hm�#�Kr��[<���E�����{�"l�=��;�5m!�U�7M�I�������I":e��u�f�<Q�߀��Jt �p��{Kg��{w[$�.��k����@����L�~��:�nC��oT�g���8O8�A��ð�,�Pd�h-!P���U͛���{<�85B)���}�� }�w�������)Ǖ�m�RI���!t�8����	��9P��..�"���C�̿%�m��>w�.M
��?}��Gk߁:�i{�!Z�^��<;�uL��_����x[5����Xm����n�2	{��(!r"r�9��?��տ�^tSh��_wL�@��|gQ�Cƍ1�z\�&E���z�Smi�-��ڴ�z �ǲ*�@ �C�Mk��[`��$ly�����ۧw�ȅ�@�Ǵcy&E� S�/�^�
�����ag�=���95�Eϝ�9��|��)�*�ĿK��;���0�0�y�Ȳ7��<aM�g�G/I$F�������`-c.�K~���\'�2E�v1cX��p������X�q�H!Z@]����wr8H4�[��`+ y;ݘ\&_��Г���Q���2��J �y���ZU�>>F�u)��e�ݒ�r
4t#�K�H4Kd�����Fm\{�v�޲���H4���V�56��i1i�`>S5���M�N����bUc}�j����``p61��5::��Y��.������y��^�W��#�	�Bn�׻2�.ll��=!�<�Y�
�V���8 �������7m�`�.9 0�kT��`�͒uL��G� �PW���Zv|��V�{ogC[]>G�&�@jD��P�w�
��#�W�
#9]ȉ��5:�)�2K.�#`��S�V�·#��F*h��KnI'f��eخ����0��5�C��ip8{4���k�!����2ޅ �灇�v_��XF4v@����*+<vb�q��~����}�f�1��It����Y�gCVk%��|��0ܯ5�\�:�*�D�-�S���S�)`��U�H�z�AÌ=�Sw�6���lI�9��)��ꌁ��� �H˼l��pL8l0�r�H"j�,p��.�AG���u�a�>�.�~��P�c��Ii�QTI�j���c3����T��0etb"Xv�ŵ��W6U:�X�\�/1�~�Y�$}�<�d�+}�r|��]��+F�4yn�\P��Q�m�;iL$��&�>F&�ȧ���z�H�*P������A	�2C�<��l�d���C��=KJf�4]�5�5����n1��UI_~֎?�\>j�9i�P$8P+P6�̒��3X��D}���=�
��m�U���xaR-��Q��X*Qo��矱D�"f'���>�n�W%^�X��_2��:��������]����U����4M�Vv:q�Dn��F�iY4��7���3	�.z��	�����N��'y`�,l�kJ��fXm���9��tcU�\mSq���\m��D��F.��Ej ;�b{>~}Q�C ����K����bS��˕%�Ҝ�VF�휹tz�<?��Q֬d�/ �#����c��)��0��v��1ò�Z�ce��0+y��_��&XM�Z��!0䰔�Fa��ұA�k�T�G�[��
*�L��U�1<���&S�� ��?h�rC���2z����<�U4@���׉%���{eE�;�&�_���,��U�p�AhX
�F g�Ax�W�i�9i/�͠Io�J'�D*M��eF�e���1m�$�\E$Va UE�v�Y\@�F��m��?0;�Ա��BH� X'�S�Et� �x�^(����숲��o��vs �*��%��O{ZC��r��.��Sk
�Pk�7�A9#�����+�n��W�˼�q����1N��������Ƽ�ҟ��u|�t�ʸ'*bgs�_x�S3��uVS5Z���0�SA!XV����(�h�\[v������/{t~���#x���^]��Z������7cE��;�t�lLs�jfM��
o~�����w��¼�\�'ĉ�^4�^l@ZM������dVr���/SG_��UP.e���ُ�b���"�\C$��j+j�&�֮�)e�D8�hKs�'+��/5ϕ(��1`#����i�p�p������[��D� ��S29���^��Q�gN�D��� k'^�ߋ��m�^�	�)�t?�j�LU{;�:0���,ԫ��M�<��ބF��*�����	b,p���,��'7 ^��W�75���7���y7w�)��b�����d�aJ ���K�/��F!����e��o��(�Bt�7fl�;Z':5Og��*ht�O&���'�x���in������V��y)YM,�X<��+�[��]o��2����Vr��3ߠ��.<�����q�Pܹ8��gl���(�D�aA=gމ�˒HT��u�w���}W�2o��/vЫ]'R.i/�L����"{��k�P7�T3�>z�)4��g�2���x�y؄ɋ���;r�\҅�����#��.���_�ɬ�6�g+�*yK��3�' l�a��ޙ�5x�Y�f�]���jn��GT�Bb�b��fԸ:����N�۹
k\�3�Kf���c��1��3���u��i�ze ��>3�a^nu%�+��^��D��1bG*�_t�na7S1�?X�^�4�jKs���W1Leu�aB�,�jk�p>�e��LgAE�+B��\�#y"��q��݉Zb��4�����O�k�9���:��Y�g�EP��4��%_W�J�y�a>V�2i<��-K��T�6�ɂi�.iy��#�$Ԅ��z-' �]��Ɉ��M*�f���4'�peG޶��=4�y9������M�yD�|[��vw��M���ⅲ�_y�f�F(��8���*��@t���x��x����n�W���6�S�#w͂��S1Î�/�6�5��E���*�ы�'�m`<x�ү�F:\�fw�MK�_��pf�!f���;�Ɋ̥J@�$���l��j���M:��6���y1"��}�<�G���5��**tQ�$"=���q��|�Y��i  *x�f�mU;g�uAD�4]�%E����Ƅ����>�����L~�c{~������Df�en��Bo
�ߊ��B_G�(C��)��x��ȁD��Zc>���F����Ky����O���W�$W��N�t�g�"A~��+0x |nd<'���m&V��-^,rS⹄�_r��0h|X�:�{�n��jwp��|�P|��t=���F(�Qq�W.O�f;���{�N\j ����h*Ь�X&x����~�.7Vx�qѨ'�-�D=��{u�;E��m�X_�G����������I�6;
�C~�>q �Ѡ� �>ϵ}/�Y�Kcֹ8��ܘ���L��~�='���mڨ��@{��Zݎ|G�6z��#-G��G��{��>Ӎ��\dU��f�b�[ ��@�v�R�p.Gp�R��u8�a-��b�.�2��S���{�⯻��j����|�6!����Ud�4}�H�n�T�*�J��3�ڲ�I�N�ć��/����DD>��?;���dщF��c��C���+�t��i��o��Qo��t�����j�z[�2�ؘ����'D���_�f%��s��e��d�*[s{gk�����յa��I:�t�����9G����<��h��H�Q�J~�s]�J0V�B�㟷@#��
�'`kٞ�ѕϺ^�Ks�|��]�]�;�+���_��ħs�Z%�4xF�9��Ֆ���g��H�Yԓ��0���7��Z@@�!Î���B[h���"_�����K=;�n�f������>!�W6i�·\�ա�]~�lr���3\aQ��{�UzZѢ15���0^�q����<!�}���R ��銯�}��bØ����DV?���K�U���z���SU����5�O���)�W���c-$�S�s�� �1EC:Q��p��O Xb�=��^1v��iLW���p��>�(��m��`)�:�O�R�'GCw�%���le ��D˟o1����aj�W��v�����)!����XΝ;��<n��*�I|݂<�x䀛L�.�!���t�|��G���FlxC�a'q���V�@Z'�~y�d��%��Ts���E���#$��g�� ֚)M7y��:�,As�MS����--��A1%'�qƐ���)�x��uq�r��&dd�ʖ9,�կ�)�5������H?NR�C=S��,�!pYoO����@��>�����C��+ ���m��b���a��r#�*���45D���J "EJm�5�"/&���6n=�wQ���������*-���!��*9X$�������[�c?5Sa	+�p
�;���;�Ł�ps�5�S���Q����k���i���9���-��U����~]1�$�.;R��,�m�tt���N�9�tO.ĉu#c�s9�dX��Y�|��_v�o���V���x`1V;��5S�F�>�އu��ȵ���:�"��}���1�D��̠�=��Q�;�x�#���WU���y�>�*z����{%��T^(��/�v�¼�Kz"��~�<Y�5ʠ؍�$����OO�ۃc�vE��bH/�vf�֏9�(�4�U��M��O��`��7��F����0v7^8�q�ƝD��b�*�=;�F56�E���| 8M�:�kEB���*��v����ي���a,��<r6H����|�0�0v�ѳ.Q�d�T�z�8���%�M�t����Kxf��H$g!O)�H�����*ܹŒ�mN�7�U�R�:�K`h����q�ᵩ�E�Cj6N���ewvy����i�jSR���N�i�j2��ԢжD�x!1�&sS��H#.}�D�1�a�b�z�5�P<�FE T�&�c?1�x$!M������E#/INq���s-+�ZJ��<���M�l'����2qD|_�s��Y���>�܃�P԰y������O\�gi~l9@GN;����'��gVU{��y�ʷ8�z�L��6g�עDe`�T#P>������~厨X+B<��4���/�K�`F�~_����Y?18�ڤWB���.MYyhs�*�J҈dр����MetLv訕멽��l���4 ��{lS�͸��Ů����l���H�σ�ﾄ��/"S��j�l$�r�l��Ǖ�n���{5}G��X�%�"��J��s��T�� f���[>z,�� �K��y:���˞�!�������+�����`U;�[)0�����ru�mov�+s#x<�nJ3U��OW�W������_�;P�z�[�L.��ޥ�Ô&r�6�\��@:��7����yn_V��	AM�����7��}�E^/:����s�!���G��9�Zc $�����]a��G��6�0�i��#���ә��Ou��5w��s��*��QHZ~NR5N��|ށ�S�
n�rQ�=Q��ىsж��L��r���Q�!y�ʶ�A8}� ЋϢY^Uܸ�Y0˃��=M��?Q�f@�W�@�,q��yp��D� l���{�
��x�IFT
��C1�w�p+�F�Leq�0�ʿ�	;�c(|�i�l��(:��zn�;�ei��W'�i诡������p�4��{ɭ��S����Mj�ؾ9c4��y[+�G�
?p��7����PC�Ћw����w������IB��-FU8rh?�9%c�Y�,r٦B@�ìd����[�㫚 ˘\f�G�~P�N-����H� ��Ds��%l���:�uqG�9���nI�9�q�><�`iIɶ�lCE��&{0#����A�y���~��/�;r�Z����x�l^ԍ��	�q�G1����J��X���_l�$((�,_@����A�=��- ��5xV����`�b�c�c)P F3w������/��M8�0f��	)� ���
&>	��K��f�)^��PO�Xc���`<��x�b�\��OS�������y �OP@�"�%	��� �o!&�#��Dn��[3�z���e�b�R"x@|7���U��_���șB��ٕ���U�N}�&"gH�=^mt����96��"�g*��V�������X�7N�;mǴ�����MR5e��D����G8(�W�9nx���ۘ& ���)/��+�Ȝ�7��v��.ڦ��� �r$ڰ��dW*v+{An�A� 0ߦ6��ݎs�*P?G��e{�z,����R��6�����Ü}��.L�LTl:��q������bh�CiY�K �tEf��7���`�����~"��G�_Tk���0�5�/�T�7��jok��k�����؟n�~����kI�q�ъ��}�x�K�Xe
��rD�,a����B)	�z*��F����Q��U>ދ�^T��H-Ī;����P1�@�}�ءy�n,�f#[&�A)4]��k�!辐�
x1XWP3ӏ'��U�E���R���$����9�kF%V� '��^�/��Y���x[��d���(�lȮu�E,��;����7Y����}zU��?t�n��S�y����i��j^����j{d��)����9�n�&+5�Zmrf�ḥj� %��q�%ɻ{{j��l"Yv���0��-�3�DređQ�D6�F����Èjh�X�*�V�� 1��A_�iv����6$���P���Ҧg-�z�|+��@�=&I��n���嚲�a{]�a��Roe82`��rI6���������x�?�1(G� �}e7mx�ܦ"x��<.���(zFkm>����_Ф��8|���`)��齼L�	��"�ڢ��u h��kU�6{v }>�ڂMY�}nň�0�ܱ6_�O�=x�����_��u� ���8
^���E�����#
��d���[�A��0��4�(qp�B!bL���2$����5[�����ڴ�z��kJjI�PZ<',���V�%i������T˗��/F�9�(����g��d㧅&YZ^�V���z�v2+�d��S�y��f�ek=�{j���bN!Y�0��L����&��(�F��t�#~R04J�Ձ:͌�װ �v��r�z5M�ٌe�m89-12)��z�V2����j�t�)%�����{\����b����� �H��,2��~+����eo0Y��kE���Vf�_�F����&�ŰI�.� �����ޓ���^�Ö�6n~lg����k����z9�W���s���!$�%��w�,�kc��ک)�(Tr�/��������>�\��9����9��Pj��]S]�b�G.6®�F뺻�������=�%�o��f$��쿠�<w.�����~�A�f�e2G�aX�_I�����a�u��V��k�41e&��u��qA#��V�xC�!k�Y^e �O.�U�1Ҳ�N� Hr���舄�R���J�~��h:Lc��	�b!~ߋ�*�����]��*�LE��w�M����+�����deq+�;1�vm��h�Д;)Fb Dͪ��H�����~�� ���2	j�S�.�Q5����3���-/���nx
��˭"<���G�V�6�<𥐮X!�J��J��>9
��9?���N�!��[!�ŘRfw���	�	M6�fkGVk}��~�%�Ue6}>}���)U�#R���0�k�`.x=�9/�o��k�k���˓d~�?#bGF��4D��'�Ч�R+W����t�]�Z��D���X�r�<^_%��=�h��2����^t`�-�����D�o�|Mn���"�s�_��c���Na�pH��m�i
-�B��=Jh-T�^�}	��Wf�Y(�^�C�ׂ���ʦq�r�c�H�<�;B�.�?de3��+����^�)7���BSm�
�����TN����<S#��s��T��I��t���(�1��.Ľ�m�픀L�mţ"�˷�kAvwV��;wx�� �c@�m�.9�`�$DC:VE�ջ�E�p�� �m�
� �- �N'��Q��;�Q��cEX�+��i5�<���f�K��F]C��5ܼq�����1	�mr��I�5m��UD(5�Y3-/ �x�� N�;�O�Z��z�?-����]+����۹Z9�[E�g\���­v��y�*�0>`X�<�T��;����c���ߑ�C�NOl����H�S��0�i�9�MV��ݧ�B�,�bж'-vz�x��I���(�{A�s�K�믳�3��:��I��܎)���~:G��b|~*Fk����&ݕ�����J �J���
ۑ4�F$ADQ���Ģ���.V`8�ќ�"�vx9}�7�9h;]��Bj�=���� ���z����#�ɵ���(�ڪ{���zg�ޮ^B�W�L���ν#RE�=�"�vPK��#�N��yt/�*��Ŷ���Ff�'���������Rf7�n�w�"���$��|.2՟mohE��3;p
5�Ɂl�e�r�;��F���4�]�xV����.a"!��:����N�A�$[q:{Ʒ	LC\-�1��Y���0��8�U5 m���bx��S��K�wdV�o�_R?� s�q��Ͱq����6���苕�_c�n
Q���S��{��m�*u�y��<��/bl�#�zyb�mft��k��%���d�cz��UF���6ߦEM#��|]e�$Tv@�g�u�S�d�]w}>+��y��D��ׄD�ݣf�[���p��Ӈ���� (�m�l�f�5���ي4��'�(��2��y�fe��6�.����]�w�J�XEc�����*Hi)�U��:#Ă�-@ ��鄔���P
|KLZ�ΐ��(��S�y�t�!�P�V;�����L�\�5h�_�"�JH�B � ��M���*��)er�齅4��K�^��y���a���W�j�T���Ԟ'.��d�ы����5��!V���d��mYq������y���jX�Y?�����%�<��j'U-�5L�f�6���=j��#�+=>=ϵ��<c��i��p��N��G��J=ݺ82ģ�k����v�H��T��S�PR�@=�~L&V��P6Y�\�}����sbN�ɇ�#l�48�j�#L�{���߯�!%�h�3G��B~��C�
�q}�{�s�m�)���!D{� �5Tv�Y��B��v��-6Ͻ�B�%ŷ.�f�>���w���B���|��S ~H���2T����^@{g �A�F�]��eN>!1{�~+���G�|h��k�cw�O-�����w�	Ga(���ݵQ%�\S��6I_8:���UC68�� $ݕ��f��_J���J�$���E= �k���#�$��^�pU�х���F�Qq�M��<���+B�+��CVB��ո�8 �/�k9�A5�pE�87.׵?����J
7bB�Mnm^�Seǖ\ۅ:+۞|s��O��p��r��.�a��6=��݆5� RK���CZ�t8�ǜ2kn�(�4Ŋ���5Tp� �B��s\���.+��}�H"�Zm��j�����9���k�N�����z�Bn(���P�v��q'���:�S������m��W�ՅO����"�΃���$Bн�e�i�P��5<;��L�<p����Q=��%�J �3�ݒ��V��c�n@�߸�v.Ytm+�o�������2�^<�r"Rq�&�ܹd�՚6Xk=$��^m`A�yj���2�����ٖ�v��ᓝiI����M7B�E�=̠0V��<5�'0�d�B
1�����5��??4��3,޳���Sx��:�F�6z)�H�Q��KQ�=I��w�cq�t�U�V�e�*d��C�̷�H͑�Ѩ�wm1��J�?�C����O������6�R��z5|�VXSuo�
�q¢��R�t�	�GK�EF���3�U�Bؖ�~�C����z�<>��z���͛�A��$P������y�1���Xo�"�_�u���H��B|�V�P6Up]fHwGY8fg��ʶ�� ��.���[-�P�.��H�)5�/xa��P���!+
G�7��NW�.%V�89�=m��^Z��cE�;b'yO�=�s�4MXUZ�V����hTmH�-L��)�������9�0���5�����)���b7�����qI�������"y�Y=?�Ag���?g��2͑�"�z�c
�l��`���~4��e5vOC7�>	����Õ��3:S.��OF��\]s��㸹�G�N��]�[���O�2l2��z����۾�����Y�(!�z��q��寳A4�O���
�3��D]����b<���"�R8�A�u�
�߈��6#�@�Z�EI�Lxյ�!��)B�xl��Z�Y���)3 ���q�&?�g W���Ʋ�d����l!C�٦չ�"%P\�����<�0�(/�/L=�I`�"������MG#�&1�ZeiD�%s}��.F-���8^��c�xQ��2�9��{�<- �`��E�,ʿ�mOf�أ����D������)�#	�I�g��ۻNh�}�ϕ�$q1Y��$4@��;%���͊#/���)�w����b���:L����PM<�xIYј��$Y{r@8L�泋����Md<3�
�]s��F�;��I�1�g��ڰ�f���$	�C���G7I��0�ԓa�Le|g
��x&h��$�/'-cR�<�
*��L�S�b��J*�J�9ϻ��j�@ZV��.󟇏_�(�gث�ͧš �#jb�����g�ee��^����A��X�	y�����F�r��������|7\ȡ?�D6U=2i��X���,�Pc���?��/4 P?�yGW�F��AO�r�l���
�hr�k���A�p^y�z�c�G7_�KT�ъ���J��x�������5)ɍД�:�J�A9*z6�x�pE��uSwya\N�vauW��\S,��r���.��Ҋ�L�[�p�[g�3��N���x8D^��}2���il� �ir��{M�أ�'�ZT�Z&{���I
�	?�Ub�k���ң��uK�3w�v�N'J�����K�,�x�x�x�b�] {�1�_�0����ɦ$*]h��;q֣H5�u�[)�o'��rO�/'��)��,��`��3�[c"6�':��Y���+es��ߢ�������3SB������-+�5/7�vx��b͗J���3p��x�"�T|��xb���svY�v�V-qr`~�	
���I6|a�z5	�����������M�%n�����N�mk����_�j*[zh[6�\ni�a��g���<�S�V�hC�)�\24�'��m�.HKh�=z�s9Z�P��g砑�٠�&����$���E���G��=V�`-{2a�돳O�����!�D�a�f�-�4t���D]�L����� ���'YY6�O5��2n�������A���痶���F�j�����!v�8N��	ǜ�5(⎱���M`�Yb �¸[$T.���ɖ�0�z/ktH����rr�D���T)�X�nA���h�d�ÙddF2�l��� !+�?w��k9�ps?��KG߯*y��_���?t�*Y��?>��EM�w��q��M��X@ή�g9xԕƬ���W��3{N9��Tr1����r �HC�=|n�YK��������w}�/x�H��|���6��=��Er��c����^l�g�4�����	+tOY�O�8Q��4�f�px�D;x�w��Yb��
��QF_f���=2�U̠�r9P�|_������W%�ntqd���6�8K�$���E�7�<��5l磃#�R��3�"~3�K�_:��3x��r��i���#�'r�}�,  *	��[��	|�	)�D�?���	6����Rm�0v�I��h�/���������=�~�V�������&��'JO�s&�X�L]�F�a$��l�F�J ����&�6䶝yl��<��}:C�o�} 
��6����$\�4]Av%���X����'���z�ls��C<��+�*�G�`� ��e���L�®�N}l[��
_��J��!g�W�H�j��BE9`�[-�!s���+���Œv-9��i$��eu0���{������{Y��G��`�%�s�8��l��V�8�S�O��Y�9j��|c8��봮���E�A�]Q��~.K���w�t��>lV���c�3^����tN ��xZ��������c�5Տk���E��7�_�Fw%�' ��B|=`��xF�����Q]P�]@?��\�Uzr�&Yq�u�G&�S1 ��Z̴pp=�W���]*��0����E�0c�ˈ��#�(FYT��h�~D��"=��nU �R��{�/�Fy�g`��n��s�5hF�Q�=����4�S,sP��Ƀ�q�8�蹉���k4؍E�cmE�>�� �P��:�V2��8�*���P}��=��<��p���I#����`�[q��Ik⿷��N����X�E��Q��!%���E���&fc0:���oYj��Ü޷w���IK�:Jj��2���	���_lK��/T�fGz��/��ta߳��5��V|S33�j�$,[H&�.�>���bb3�
�7�S:�~,3y��Rٗ
��{;P�����ͺ��!�xU�Y)c�����K�=��C�Dow�(�j�R _�����Gpo>Y�'_ַoV��?��;K��<;�}�:-������Hֽ�m�HC^ ��\
:˹������B�,�r-�M�H4f��]�����Á�s�Q?/�#��S��*���|7���b�[��"�{b���q��)����ڱA:�������1�����-w�ܘ���#i*I⌮ys��Ҽ�,/�ȸR��۴�D;u�.�Ax�,<ՃM�-1��Θ$����]��y�⮬��-��}
Ax�?� pL�{���$���O$.|ʼ��CĬ*��H6��/5scL��.i��?������{�3�8]j��xꕷQp_�mѽ��6'M("8�sm�wAu<L�)�遺oCl(��'��D���� }ȗA���믄����7�������(Y!�8����q5V��X9@����ΰ��NZ�$�-�z TĬҷ�|`8x(�����!-ŏ^��>�~V]��h牮��fp��y���r�#N	ɑ�*ط��"NоF��;�i��Ƈf/�����8ۺ� �1����ɹ[͓�y��,ɵ~��&j�wŜ����x0���5,G�ZlD�|c�GX_6��~U,"���~�o�|}#���4U�����:QJ�	�>gAit/�tL$��HK�����������O��A�7F�����y�4M�3\e�%ü[QNF/T��0(���`d��2�7��FF�奄����?�����Q�P�>,��u��	f����[a�,�,�D�P6؍G��7'~��/�oI
�,g�sZT+�/��/��p��T���E���ώSz�17,�&�@ SNu�Ye�a>��"��Gxr~ywK��۩�U8�d�	��7���'��\��_��ؖ��SJ�Su.5���7���������n�|OyI�g� 7�vߪ�n������NV�����	�4��6�ap��y�2ݔg�e(z���[=��ﴍ�#kHU�`6�����L���?�C��a�rwJ^��]�r��8����<d��Tȴ�-b����5�f���q7ͱ�;qp�Xy�����򄟆=����������I���Xp��kNR�f�m6�<ke{��9��yi3.�ؼ<J�D�-��(C�"	�\O��ś���4l/3�w���uKSxA�_�2���
��և큷tk�*��=L?B���*�Y�hpֿ�a��z�RƌJb���ٍ�)�?���P[����!)?{�4�"��!��&.���A���>��ث�Y�1P��$�+,�A�F��SHɩ�p�;���m�؜l���8�N0X� 1=K����4�����e8tk���i�#��ۍ<��+��-Kq_u�d�}4��Jj�2O����l�,b��g������.�Ɩ�������FڽМ,�J0@��9!.�9%�:2�⣧Ի@ʐ}avcĈ�}N$��(��Kcj֓�(pƻE�،�M�3�3N�(������Q��c��4����@�^�e�k�]X?	]�|��Jμ�������	W�eB��"?ٙ�1)%3%ӛ�F�TSns�N4�e����d�:IPJ=�Xb���6�k�V�qٷ�wVj�;�+6�SR��Z�f#�W}���4S�[��z&PXL�J<ﴅ]e\��˝��t����2����(z�yJlm��/�(���3�V�A#�-mR���9��C��y�t�P\�%�P�m�˰ uj�
I���,�rb���J���S �C����akG����H�5�Ӛ�#��M�s*
�m��V�|�3��;<�i����3lg���0��<�}����R�&���o�q��uE�/����1���P���x0�V����Z\'��{���o�ef����X"�/�ݐ��؜�Y��&�r��k�q�i0��-i4��f+����i�v_�a�e�ǕVB�q��ƻ���E.[u���]pe��`���6]-�K���U:Wsh�ƿlځ���Ɏk��r���Č��	Za@з^��}����k�!�i����<f����U�6���;���fv��T�r=�K���Pe��Lg�36E�E��˜�����s�n\�]��o[!�.h �[�V~�� 2��2��p���\��M�5�|L����PS��
���.h�!�َ�R�8�����^�s�w3���%�?�$5mb��g�:zD*hU�dI�Iz���H���"��B����� �<�FS�Jv����XxH>�B�ȊWXfq�g�1]y�q*��_�o��҆i����)aב�w�r�G�"��Ί+��E�[�ώca�Uz��Ehe�e����c�rBA�S�mx�|�a/�r!�x���� ���AAS��ѡ��.����&�K��Dْ��J�N��*�$��]Ź�qf�t�g�p�I���d���W��u>j�BVx�W*O5��6���1���fF���[�Re��͕����kФaj_U����0�P��;緑Đd�I�vN*�E�}�1��	_zg7���ꂬr%�{x@�ϩ��|ܳ,�}u��O��d��i����Ǎd�/������7\�������L]�(`bhf�)q##&Et�i�W$)hf:�`06,��ˆn&l��cγm�e)�Ig�-"�HX���C/; <���
)>��U?�,s<k�}��׍���?���,~�����sOr��?���g�E��;ꎗ��#�8Az$ی��⚐��?.��d$Õ��ø?�r���CvNxOW�Ї�bFś[OwS�O�d����O�-A�?�նC�`�B����.#H23��o<�UE*E2c�2C�u��޳�e���5���r#h�m���
��w��e��t��C�ɧSɼ��E�E���^C�`�t��j�if��0a�o��{�S��HMZ}w�L�)���/�X�D"�*�#e�G�f �
d�-�7AufB���OIRb��{^WUg��u�~L|�q�9����?pN��1�p��9�p��0I�쎲�?�5�A��Z�mJg`
�� �ED�y
WNg�������l,H��j���,�3�b\�Hm��y�0&�NO��@�!}}Цq�o��˴]yid�Ȃ1a�Y��hx�x�י0��υkƃy��h��W=N䬐�6�F7]y�V�Z�ٻz�n�9��o� W)�D�]���~�A�,w��(�[%�>k{������V�e�zDQE!���u�9���%�E��L?��1�ʇ���� ����Z��}[3	�TǏ�,�x ����_-�{K%�8L�f�OTcx��/8`蹇#� N�&/�I?��@�%�ߞ�S�K�Qj,�N��7@�_�%��XH���T�jW-��W6�O=���|���۟K���^��F��hB�|����,�QHc��$ǡ ^*��yt}q3�T@��+��k����p�thC��H���	���|�P�n�Bk%�w!�O�����gj�w���+34i.�Г�������s"�hJ�|mY�Y��&��r?ЩLY>@�W�5�X��Z4X�I;���͍
:2�,��R�t���E�����"��.�`��u �/g;L���h��3Dg,�W����'�ܻ�[��p_���mv�"3x0��`�.�ˊ���xn~~¾ *4�Y�?�9��?�r/�z]?�u�)��pQ��6��vË�	��a��ʾ`��Z7���e�[�X��	+��c���d&�ɜKum�Zm�#��l�:Z��	`A�{�Yu������ݘR�'���]ŵS���K�������+�t�,"�ը획��h�렻����/m�6����@3��#qƬ�~�2�H�Avk���Sl$�P��h8@M�\�Z43Ov�G���ܾ7����<Λ;v
Qz��-�/�ǅu����Ц����&�y�#�#^
4-6��L ��e��S�9�݉o�\��N��[[�F���j��j�:#��#�k^r�3 ���D7y3$2e[�ԍ3^�{���o��ё��n:z-�/'�1��$9���V�=�u�G�v83�m��_��$_�R";��F�o�Uڽ��Z�-vb���HG�1l�pH2Y~s��uo���3C����`̴�OAl=&1/�q6�n�vY/lR��&��&�Þ���^�kQ�c����Z�^%)V�	�:�4�}�ߎ�Ap���v 2.8�#����9�hji��,�xo�ֵ 5���9N���-�@��`��Z�fUDX���	���}}l$o�s�y�?5�r�4��B6��N2E�����TwOsڏ�����8���ku��b�Gj��V��D5���n��<n�Q��-��[�um�l�K!��x��-���2Eٻ C��F(^$��W��R��D�l�L]D���"a%N�N6p,�:�G��FR�7��^0�B�
h�u3��jS<|�y)'����+�D<^^����J6BQ�.ו;�}����`E�Gn X�����y���R\L3
�&W��~�}8����r�|:LE.tD�m�%�\�>����i��4P����̹���6K��?���_���,�"w��}ܶ&7�F��b*��ۘK�kkα��Y\�R���IQ�2}�H�M�ɀ#��5�?��32���
A-u'�%GIDy�]�6mf�i;Q����M�K�e�2ݞ�M���OǛ�nScL#uT�����p��i��1�vZ���E,i��-��Vt�m�����_�{�X h�����]�������R ^�Q���h>�z��8Y���l�[)hh��߷�c���1z=��%Kv"�K��1DjCl��_���44iM$ d�VɞME=�	`��3��d�a(>����P�q��.���P`fl4`���ԗN�ݮB�ܕ�/��3>�z������e>$`$�M��K��]��� �֦MT�F��Ȯ`�ħ����V�[�q��e�j�2�z�A^�[Y؈��{fd� u�^��W�i���b	��@�i{�����N<{:�L�/G��}`l�u���.�[����
r�HNFt'ːe�ЏĐ	�;Yz��=�(w��@�N�����a�k���;�<���9;�<6J������g��-�%"h�N��7���ir-�>kY�x|�j�yL�Ċ=�Yh��2�'�5�3C���v�M9[�� �^{:�;q߭�o����ԋ�Gg��D��-�E�����KX��L��B7�y�V� G�(_�k�����o�U�B�	/����B0���`�F=�&�\�ivx��j���Ds0b������f��w����}Հb�Rɋ}vj�"��4K���4�I1K��9���Bm\�~oj��Z�G�2���_��+�^�Mό�Z	�rZ�]�y��Y@#Chy�	d~b��.���g�v[
T��P8~A�vI�Y��@`K�z��#}����N]Ssv�&�*�36h����78l-ޔ傹�L+�K�����y�.{�ӄ]ܘ{��`in;P�tH�Z:��ð����P����[���wʴ���r��Jk�_j�����U���&Hw�����/c"�e1+*i�~Q|ē�J��ǋ���Y��nd�;I��bƧ'J�R�<1J�X`i���5�߂��ej�v*=��Z�6 @�@��uJ���%�h\���Aw%��g��a�[�m�i�H�Qg'O�+�8��R�z�,�\��?�߀�f1�#o������߯wo�WPI��������P��D0v)0��:I<rv�v�+��'��yG=B��n�z܉���}^�^"L�D���#�e`¼�%��%!�v>���z��aw����bFg$����1ܝX�/$�7	ca����������H�i���O�eOMN蚷�_NF�0R�
��P��U� RJ>4���ެ~�ה���V�tޭE�'��Us�N���^���m�	Ԟg60^ԉ3*���J
@6*�O-��f���vUE=��,|H�<�|�!&�pykO�M��}�=`��W�8��K�Rg�Q�M�����nT�칭�����x�d�R҄����^���m�b=�^�V}������s���]+Fg��$wYg[��.���5E&5���J!��) HSC�Z_�v"T��8���oȯ�U+^(D��G윎E� �j�;��UDH!8U��eL0bW~�d����8�9 ~���ˤ�R]�N��%�n��/5����F��3������^���5^.Cƛ<����
���w;]�U~t��U��X7����δ9J��F�i0���}o�{@���6�e%=xc�f"D�����>�{��T��5��N@��p����p��U������/>����I8��=�)� H��� ۤ�[�e~L�)r�E�T���S>����Em EZI"�Y*��Ҋ`�I(r@�L���F=�,|�rA�M�M	u�7�/�,}�a�K_���-��G�W��Z������]��!�~��ͳZ�5�r��7���/�=�|O3g��	����2�Q���΅ـlSŉ�~�����]�F�=	�Ƣ�]��,'vsR�y��� ���J7�iS ŭ�M4|C>����Q<��}�4���y�U&S��`Vi��+���(���K8�oK$�T/��a񩄨���o��)aS��E�����߀���
���e~c�r#2$�J�A�Ei%�
���-��W�㖾�'n׋r�WZ��@��7�[�2ɫ�ֆ�F��o9�Vm�w{t�{���x�����`�h��u�p}J���i	nol�WnJwP��������#bf&�AJ2��0C�����Mc�!�U.�xiL�3�%��!����xa�����ϑc�G��h�fTO��F^��6�[3G�3Ds�v㊪7ty���0%
�)@z��(@��|;����,�l�T\GΎ@\�������d�K�G�Di���򘧿���oOΏ�hʷׄD�MK���!���ڮΌ}OM&!�R���b� ��d�T��M2���)�V����h`���ǲ�!J�#��|mfP�jF�-�K���o0�C��
V}ʺ4���&��:�%x�E��|\������������i�25O�}@�	"nφ��i�^�CV�ܪq�e�#��Imp@�Y,+!���*I}��>�/w�Asf wT��R
%E��N찧Ls�D�ǫ�;Z��2�K+י����ŊiNK2�+�A��csaŪ�NI ��*����x@�f�n�ߡ�Kg��VJdaW/�ț�#���?>}�����A�n��}��_��N������_��dM���b�Z/�-�j�֒ѥF���"쯔mnv/�y�wQV��x�d���4����~�e���{b��,z�5y�K%9Yx���
ɣ��^.G}aGr)����B����0�gp�M�(���?�\���!��\��!�Dz������F�{��.4%c:=��'$X)�/#j��V�>u=��?)��R�W��k+�|��H4)ⷚ���O^mx;vv�h̬>FP¥k�
�� ��)7c�ii͖W�e$9m����"Z;���N�e���
⩁�ڍ���g�	����^b��,��ޣ~�Bͪ7���m3��ʐ�Jo�)yv�������Q͚�6e �WY�t�{�(��p/^(�L �q��g�,Ɔy�z�(���ZwD��b�5�)�JY�v�����it�Ҥ�/�
GDqMD�	����vUQr��� ��q�I%���>���SF��ͨ�I�*����mj��j
����%��<o��8��p}���X��i�X./
���rn�H�~��]��F�\8�*.Bǽ�M"�����_�����d���6ɘ��B�m�Uc�`�K#���`��?&�_�;Zү�ڽ�r3���������6��j��@C�t���2J$p�Wh\C.��(�J�V�Ni��L*����0����Fd�2�H�\����e*k`<|�ޭ���s�[J�8�A(� ~�l0y�yq�E?k����ꅡM�_�dr��H�	[5D"�)~�Е= �N3|�p6	w��]:\�W��:,?�1�K������#�kK����&��Bʓ�o~���w1�Pk�r�g�t��\?Sa�F�~�1@w_�NA3���\�_|��vHĚ�䜊	O;����I'(� Q.+�'��{s-�!����"P�"=\�����c�?��+�/]�*ds���3�G֫M|]�ʓ[�o�:F�ē�+O��'��-Ө�S��2�\��f�+�=��Qxr���|�~�k����[r�P���,��F������t�ݫ�}G�����>.4CPY(I=o�(y�\{��8#kD�D~��0�Z�G�'�����)3�V��p�X��_���V,*cmaI�_����י>�,j��)�R�j�u�M��u_��;�0�hp=�����	��"L����f�)�Oa�ֽ�Xz"���r��b�ٽ�P�k�)�9����i��T���\8G-n?�-U���L�BU����{����I�`,:��Y���\XJǐr��R��
�=��\�xy�6^�P`G����9b�=��?�g�Q����H�����,ۅ|�t2��j� ����L�	�׈��$G���Xc�#C�B�?�-ږ�B�O���Ј���e��y�=Qǉ�
�ln�o2A�j]�C&m*��U�J�O&��l����2*7U9��y�O��!+~�g�/�ZiB�}�(b�؝�R���ǹ\��R�V�miY#��8%d�pu��ߔ�"'uj�#��W ��[E����W�$��!g��VT�W��[4l"�2�pR�o���)�ɜ�0:�HH�s$s��Ls�ǋo�p�Ȉ��|ݨ)��x퇽�e{y��L1Z�E $�X�����;*<qѡz)�@hX�H��@<�h4��+���N�s���	PM1�Ѱ؞��F�Ê�Xv+��xJI�$n솧%ހ�]o����y�¥
כrBT�/Dﵣ��C��IKӢ��$��>�9m�W���hu�\s�a;�Etm��1��^C��� k7%�5*���U�!`�`���;��Tb����|�~��f�)`�M�
�)�>3�P"�� ﲂ;ά��ARo�R��
�L}����oL�tm�����v�m,#o3������(�8�(tr\!j��>|�u����������	7��}�[+k��]d'!��wP*�)B��-��]��hN��mm/�v��+�2�l �GԫV�O�T������qu�����sFG��?�E���.W6J p������#�y�ZA
!.K�Vy5�0C۟|8B�Z�CGf�gk�4s(��.�5M�bm�x��xv��ڴ4�7ծ��J�Y�`2md�+덟��*�����L��jr�����~x�������ޕE��cQՅ�{J��Uѹ�-�־t�g��n��ʛ���0S�<���J�c�[�no�$���	k��{�{ط@��P�z�*~f��Fr�KZ3��ĽDљ�Y�"�S�,���:��Q�:ɿ��%���j��ڇK�k��F"����N�.vՁ���qA������G��A��Ț~hIe��ɪ����>�L�j����2Wkm�0�\�k9��s.�?;�|�@��� �^e�[[�ģ�Es�`�D� V��S�X6V���sſZ�b�	?rC��(�C�O��&fO,�,�W��͠��ɜd�
������}����ĉ�Zm�q�-WR�CF��e�_38����c �G��J�׺J����iz T�A�L� �*%�sX�H�M�J�?�Cufx��z8�g��u��ډ��-`��e)2���6��:�Ӑw����D�����(\��ᑎL��~��C�tD_a*�T���������//�1�Hr��;DM��� �:�M�|��_���8k�/�����&��ğ�&0� sMT�|7��C���w?�����O}>�TI�jnC��[�c��MQ�X�t�Y½�R����m�-�aH/���]Cϩ2�4�R�'	�f��V2��{D�w�+�Ď&ޛ�/AY���1����!�]���Y�t3���U���ar|{��4�c�c�SW���b�}�^"�{�#tifX�<�/����&b�O{�"��
N^p��͞wg�"&F������z�Y������p�mm=LRa�e�1w��M�B���Wƨ���~?�j��N���xa��CKY�D3:CG��)�Cؽ*����^t�j/#cu/�5��������꟭l���y��"���e� ިBYF�󙤫o%�} ^R ��R�)=��!�Z;��{�j:�I��%�St��J[��E��w/W�r��1�U|g���_j��!i�"k��i,�u	|F.��E�JTk`Im��.3oB����ݳC�8f3��Tl*��H�Ռ�'PPП��+MAs�ѣ������
ag�R�����Z2�S%�����6�&����������p��a� ���ۼ������R�v1G������$;�����?�6��3k)��F/mDM~M����X%�ř1.�����C*㕬��-6]��~�}ؾ��"|�j�6�m}�����m�9��y�����/�:�H����X�9R�^&��xM��h7m)�_�r�M���.����26����{���A[W�R�`T���g\�-�Ku�*��CƗXJX���4���?γ���s=^k��U��ʢ�Lk��:\f�G��e{q�a��+Z���&��B�r,F��7�ۊtXzW�V�;q��x���5f$.���d�����:�Ʀ*�0l��j�@�&�oe�e鸕N6��H�1`�HA�f�� (��Ȧ���S�D+8��f��䭴��r&��Mӑ6��0�c?j�.�NG^����'�.8�7�s#c��~Z+L��Vɮ�}���Ng����$�$��O $��uo��4�
�4�����ʬ�kb�.s#�6�/�m����83����D�x��\�h��zXD�Rcb�ֈ�f��W��_=�k�* �����]y�u�*zc-_��G
ˏ7j�4(��c�m��+J{gǓ;���6��Mo��A��=��*M[OV^�6�&�����h��uf��D�j�/ʔ��:�a���9�q�M� U>2�6Y.%p?��v�?�t�����LΞض��aV��7�W�٬�o3/J͠�${�U�xn��?|�c�a�����
� �A������+����?S��+�pްqۏ6�fB�Fl�m��W���[Ǿ�%l� Ze��a�����V��װ$u5��P�,��*[$����~��HCb�b�a�f�R�r�#T�
���Tkg�.������#O�Z>��_/�GZY�=��Ξ���+��m<;bcZڐ��{�LW�� ����^C�5�M�;y�)�NeD%�y��R���v�u��й3�?�7��z�<߶�άL�D2���;��Y�H܋��^��;�9XnYcx�G0�)(�>������$.�_�K�վOQ"ʞ:b������cp{�$��dۀ�ǉjB�a�`t`j@L���M]jT��@~�Űv{%�nr"��j:�/�W=5�3��$��w���!��Xw��$�Y���{�)��\}��ȷ�q��5k��ZS�P���d!zJv�μ��FaM�c���L�J���ǻ�"EhH�g;Z��k��0��Xv�()��S���� f4/��Q�p�1g<ٿ8�6뙑3�������(S`ڪ���5E'��%�(�8y��t���!��+����s7(��hF�"#�W�[�,Ck���dΑ�A 0u�{I��ۗ��2�� 5-��'��	R�O��^E�T��j+�)
l#%y'�̽x}p�p-|_�U�D��`�r���V�P����Y#8_wu��5U_�cme�3����7єL��ǾAa�4�m\�vy}C*���˰+�I������A)	V�t��*��L�5�.�1A��w@�b�o�U��lI�U����V��I=�Kԣ�d4�Ǧ���"���e>��{���GBCƿbG�f�Q��FT�A��?���J�P�'�~JEM�ԥ�t�!����7Ae7���u 4�
`]�P�O�P0��Қ�6�2�	��&�H�>�6&MV�lӜ>��Տ��}D{A;cn���tp0IZ>�ȼ�ELD*T@�W�Q+U��ӡFv �$�����{���QoqwI�P��o^Q����z.K<�eZM�Qk�I8ݣ� �v[T���l۰zA���R/�s|V�Y|�hD�J+Yr��+�6ۇ���E�W��ZV+�Rz]2T�:cd�u'3e\gv���#+��	�P;mnj'b|!
�:���XT�7%��};���������>f�+����*8�Z�+�L�AJ���)��M¤����� /G�/����e�t�$����;nE��RU�tI`��0]�G�~�Mk�� m)"�vbG�s&��>k;����.��Lm��u\`����
�S:P�F��1��>@�i4+�&U��v{��n����~��d'�d4��ə��1I����3��$���tŕh��cD�adʀA�z����Yl�M�xw���2딞�|���i����	�rfW!R:�a9�9g$D�N���:�B��Nd.,{���0��`���.F���e�W�2���$��7>�SpĩE�z1FE^��:�E��C�^=����mE��)�ڗl�<R���+ض%�4�T4��ws]��B筪��!G��mt:(����,.j�{l������g�M�s��@�@#T-�)�a�=숩}0��jF����:��u��Y7��n�U;hR�Oķ��lhH�� ��_.\%9����[��b@���#j��w���nдS�|Ε�R�hƹ�d�:l݆��S�5�Uhe�mk�����Q��s(Y�6�}Ll�W�6�"��Su�1�W��� JD*�$����AP���Ș�+�V���wR��@Y�eZ餝����ڈ6�"�����a��{1{.�fXӖ�.h�w��,E4�mF��DS/�G*�0���:�g�T:�E��tX�Ȼ»�Ib|�6�mviʓE}4y,1k��<�_�;7�u9hOq�UC.8p���D7�㰋��&�W'��֙���l�ȁ�My㺠�m�������l���P��X%��i����*L�/W�Y1��A��kX��у^�9���i�7'�ħT�2���T1Q� ���H�r�^
�N"{��9U��0��z,���E6��QΈ�[k9���O�<���h�kb�����f�����d[�����`r]����Rx��I:��b��I!�q�D�(W萟{@�C��..e(Y%����c^�&U��e(�T�K����<�����w��ͫ�#����/ҟR௉�7YH�ѓ�K<����q�������J	�Kws��${��=0�p��Ѭ9]Ƿp�=�u�́T�tV�b*1��.`��[y�gB�w�����v��/3�Q�F��VKD���<"��(��u ��
;����r���Q�	݃R�f	&pτ�F�1<	5\n
���կ��#׼����Z��|�c	*e�k��g/�#��B>5P�mg�9]��~�N�
T9��O#�ޖq$ѵ
�{ҋ�.o���Q���O@ՙ"`����ڪvi�4q��9gU4�cR�	P �\{Ox\����dw�	Kh�{����:��"RS�v���.*P�aN��'�2M����P���lT������?���q�_�@�_I�b>8qr��FO���nP�V0��<w��0X��B�BLwW?/h�?3mTCͬ9�3��S"�;�Ty��9�5�!$��6�2�/��˿V�P��hw0FZ��\w�)g��B��2Z�T�p:rN�����@���U���Z���W��%J�����gx{��I����	�~*�Ԙ��[)D�d�m�G��!^�EAI�\�Ǚp�'��6R6����� �g�u�M`��:Nw[�U���c�E}��; �|�E�%��i	-T:QK�G��V'd���Lq�H�R�����%rF10���i7O4rqo"�"��-�(z��)[B���%�q��\�h� k~����D����� �/���P��b&&���5:���}e̛�CD�9!�.�nҳ�[�7a������Z5�f�Z�y?s�IQO��W1SBϐ��G���U}�b�>3��+wj2VP��r��˧�L��t�/�B��5�&ѧ�}츭v������ 
��tX�"�]��@���>�����F2�;�ȉ����">ƩS�#��t��/���T��R�6	��o;�9$Z⽟/8|�K��t��`�}�.b�F�*�G@����+\X���1�@��-�j7N�������)���"b��Ҭ��q���U6�Ȕ�f
Q��}�]�#�2�����?ש+�x���X �mR�W�u%�l��A����?�́s<4R@���x�&(D�i�Ajk��M,)ia��5h����Q��C17�<�n�2�#9�.^A��%�/x�~��@���;"D���IWKVǛ�K������B��E�kANwR�3��_o�H+��D�翥�AR�K$�����70I����o"=׽VQ�H&�6���`��B4%���J%�TO+�Qe���ֽ�xċ<w�
R�R^�'XpSP��-�����"x�	��Ö��	���+ݯ'�c��tx4
FeG��#���!�\��["�=�4��U�*sA�٪�������5�����h�YZAO�*BM�(���|�R~�֜Q��O�a 8�P�L�tGe%^� ������J�K�����*&����8"�#[��=�/X.O���� 麃Ȉ*�<)I+=��Ё�i�ǘ�!�¥���A>�#��o��������Di$���W���dl�h �8N�jy9G���!�!;d�]��]�7����~���t��v~�a������f��*��%�Y���)Y*����Ne�zg&㈠F�H�k�e�������="!��m��{�ŕa z��	t4�Vk.�>����.D@�"!F�r�sƫ\�!,�V�{�Y�8�>״�ziB2o��'�8��CL��`�����N?oc�'�)<;�^\�Y)8����_��`����{?�Z�<7Ù��V�Wὸ>��tvL��9^[������6�/uK��k��SD/�Os�& Z�z	��9w�?�i.D�֟�i<}3ȑ��m��������>�����mE�]@���Y9�ц*��P�0����;����[P]�r�ӯ����\G�g�	��� _�b�H2��, �Y�1�?�9A��Z�`�ѐN�l\���	�?�ՇKwW�0�ߋV�{�hS�	}
<.�2�W�*M��x�Ҟ����/��a5��C����y��;i��l5k[]����*�Uީ"#	�w(�̎$��{�SA@�
|f6 l:jo��:M� �!��=��4�\/�G�fn���+�j��&QVrJv1"�A���qX��Ǹ'{���ϱ�����HD��Ŕa��2k�2@�F��<��y�����{UWD��R�7�!jΉ��Nw�R�e{�T{���L]V`z�FɁ�z�Db��k_�o�G~!�sL|��� �p�r 
�@��F�Mȑ���=n�>�9sIe�:���)�)�J�Wv�Ғ��������`C�C��.�'��XC��bx�=`���O�T�Gy����ca�ʴ�dYΜ0�ܡ���-���慀����������_|X��z�i��a�]<�i���'b,��}'ojTO�����"�Bk�]��1YƠM��#V������˛�w���E�ٿh� ��0{�Y�#����J�h0_9y-R�qF����������I�Y�����E�Q�����#�t1&������ˬ_��wPE�Z"l���iGC����ShXno�G��U��O=���%C�͌Ŭ��O_�f��k?
�|�UȑPz����	ymD�,u�E#��Chc�Y��XZ��M�yr��j�$��@"������e����;r�H�儵_#�`�(��*�4vO�ŋ�F;1΀���1�,�_�E:�P�IQ��3F��GŦz$q,���T�R���e�ጔߦ�	����r
����N��D!�i2���q����w��Q�ü�=r"�eA�ۤ.e�|��Ȣ�F��� �o8�$Q���6��Ӄ�v�-�}��"K&��5KZ�f�(�,�_l���@��ܱ,���J���D���嚕n��-��%LRAC���aDl44y��oa\L��h,��-���ER��2?��(�H��n��#��M�/TT�;�-w̞���x�T�Pl�2�G��V�����(��K�1M������f|���McT�:�/ Ɵ�O�ɐ��2��'�1�d=u�}��Qa�ߪڝ�e��_�i���r�zm�q�IJq�
Z{��]ߜ�jj�V�5�0��ah2.�J/A鷊:��L���D<����15w����K�1���Y�A�R6�ړ�1ȍڵ<�}�NJ\���@���X�&���?ژ�Lg����Tk�:�uiր h��Kh�P�m�U�q«��l�ݬ��oh6�A@ �������hH���Ǭ$��y���yW����l[!/��L����B ��G�{��q��UG|��LR	�wDs��m;���ɸҮ�3)}Y:2�� kjwM��&WK��)�4��'�/%.-;���L����G:�K׃��A[W5;Y7�b^)4���s;O�ے���
S)!�ur_Ec8��Q�vJ>X�X��DTS���趰������	X2=����dHb:h->w����uU�����\*@y|��nZ[�B���랕�1�k^8�&f8��� ��&)��v��V�����B9��F��-n,��?)��-�pKr�V`'���YGI�<�7T�X�iZ+����AB�Ŭ�v��т���k�,6�Qˍ�Z��מ%����������DY`��N���+�2��yW��Z1�0P�=@�������p[B��UK�8G�&5�^Uʐ9>,w���l�.��-#4rF��\r��w�?���"ב���H�Š� ���M��UN?���Jmί!�E�
é;�p��(�$�����R$�x���Tag)%䀖E���R���
��7�Tf��]X�2Z��oT�Ȍ���^BQe1��SbE[�˂�V����~�ҀF�Y�p	��Ю�z�jU���9���Q}��K������s�'2�d'dC�Du�*�+���T���JE9��ɛRp�P�d�����ͨ��KI��N���%��R�>>����1��P����sdn���c�0�0�0��c�Kj�o�K|��:�'n�'z�Q�e̄����E
��0����d��Ӈ>	�\�ё�ἶ�;�av�^Ŋr3��B��0�`:(��M�궉6���n�xJ%9H�N({~��\0�l1��g����T_��~�_�X䏤x��X�e�ߜ�N=�M��j"��'z��m�+A}�dFƔ�hW�O/߅^.�JW(�Z9P��ty�W���
FE g����kA�$��y��O��Z>(�6᯸XQ���ε�D�0ɴՙঢ͹w'o���+$F�K�:�$�_�SJ!I@�J�rb��"��)�<tm$��� ��Xwu[b�8�F������H�^��k,��C�>yk�<�j�}�r�d�y�+���/>�o�Z�C���=��2�et{wd;�Î@q���ǖ�s���Y�D-�H�S����d�����ZX��[����Q�"q�<Ŝ���g)B[9
���d$�Ջ�,������E��L�V۶w��<7�N$���.�+�BH6dX���P6~�V{�/�\z]�[<�_oyB�N��]1�&�ڦ�+G_+/����=c�]E1g�I�4B|�a/?zd;� �9�E��e��u.+9���M`n��y�m+OP��8
-IiI�3π��a1��,,�<X��C�4�T�ua7ILEۗA��xwh�)y����w��J
1��\���I�R:3]pMU�%~i��@Ӽ�4��� X�t�Y�8)KU:QA�����岢kw���t�]rq�%�=�xd!K?�!'6������h�(��be���uv�lgWѾ.����\�Ł��U�x�DjIR�����V6��%�,�����Ā��/�r��&y	�G�;�C|���R�*p�q{��}ɘ�c�ޠ�I2���$�fe:-~��%����R�Xɺx'��1\�%_E��vRg��®�6ʝ�����G���z��,��翥|�x1
�0��Y��	X����y*�i��D��Y�?��V�
w�����[��)=D�36�pg��̼E�¤I�9Ӆa?l�P���d�D����ǽ������n?VA@�"�������&!�"�	a��ݰ�;��	��d`�dęh^o"�&C��i��d_d�y
?����꫻N�O�>z�t�2��"}��|�a|n	Է%>}��+	i�@2���٦�j����l$bFA�~�XA}��)F-0�ׄ!�7���s�X�k$���[����Jun���r�������Yv�!��d�7��C���8y�<�� �]� ,�tm&.���F:�>�y���f�|(
`^��?grY/Wۇ %%�"SOp���B���!5�>+e�\a�Vq�<ɨ� ��%�A�[����r��wSN�;Cz��k�,�|O	씅`"[#H���-"�8j��A� �F����T[W5E�-WZDz$�-c���<R?]cP��.(}�X|��ܗ�9�w�}�L��K�ś���(����߳z-�h@�1��80	Y1)L���9CG��>���i+�'���,�\}��C�h���K��O�]h^�e�$
�?!���cf�%��v���#�����LbI"ɺ(E�ɯ�U��M|��ݦ���XL��U�	u�؈�us�$���3I�ǡë�A:�۰B���)�΃������紧�0�S+N{��
?�T�0��^�Y�+����X�L� ��l���ց_4����T�t���<�V�0��[�z�q��U�1/h�||�sR>�|?����@jU���%��^#�'�> X�eT'���g߆��k���Xw샕��w���߶.���Ֆv����5P28��𝮗@G/ f���5/숶ZP����͘g��t#� M��?�F����M*�	����҄�����T��f��:y6e����'&g��0��䶨�Ɣ��L�id�Ųl�F �����Ōe����O���'���:_�h"/ʗ}��H�v��w��"R^����,�<9MS���&�Hq�8��VbF�a��>uu%GB^W!�=D�V�x��z���Ń�FNS�?�
�4
�=�Hk%o �N�7mB���hˤ
���|b����U1\�v��Q�|��`vS�*����)�vRY�B�������EP���,v����}/�f]�߿1�0��n#Q�?�t�z}���8�ow^\�b�+K�@d@`��\�F����\�ƅ��A���H��"N�U;�8�����/=�pᵆfJ���_У�i���P��g���Ndb�#<���C�6��l��x乌�CB�	�@Ȏ=����I�P?)G�{Pa��Q���A8�`��r�~����ɡ5z�����G����H�Eqz�t�3T¢�P���IHD�XrlO"�#\=c�|��_���J�+o�U�s��̨^]G�V���y�'ME�i��l]�r�OF_�|[_�iD���V����R<k��=i��}�+��v&��7�� �yC��K��dx"~V�(��m�	�́����0ӵ�~�|f+�����2V�r�ι���Fq����X]Who����0��Ӄ"�$C�'��"+5���uN�P�Cc�;����l��/��Y�f���|K� ���GJ�ҙ���|h`�5�y��<G[�2��`�����%�(�9Z>�c�=Ѕ�8��^BYM�������=P�C����K�}"�_�Q���4rZ��^?TA��y��"ٕ�����'�5l=�7�,o�8霙X�.@D�����+�ص�""lC�8�~��r�3���J�-�}�����ObR7"R��BϵE7���(Oꇸ5ĉ��8f���t�d؜��!��4���lROԀnM������<k��P����Y����J#��p/�}E;;�j��6���@p�Q��7ƥ�9��0G�����(Й���_���5��a�49=L��{ӯ����{$�s=!���+o��" ���P��K(��N���|��b��h�9 �Y�r��多8��v�I)	�l�KM�n��5T��d��yEn�ϼ�6W�j���+iռ��LΪx%r`Nc�OV���3Yy���^�X�������S�ύw~+[�����cǣ�+F�L���v�cq�Ib2P5~_�;;�:O��������@*��M����a�� z�Ejg�7�03��h��u3�e Era94Y*�9�q!�z��2��ô���#-<`�5s,J�t ���e�ii�?]#��bX�)�ă�x��*Nj��^�Kz�7�K��2tp�S�6 �V�Ml��T�Lb����6��'pE��l�!#��OG���VP�<J��6�D�������W�����Т�e:�&Vb�Ϻ�FgS��j��s���"w[5��+�R�0z���D��Ҽ�O�8�����G7��I��)@��3i���^G+ű6�v\!�h�����8}���~[�K�=��&�4�9�\���2�%�%���%�ꣴ[�8�Q�9P�L�X�/l	%la�N�t��aw��7z;;ʄz1By�Q]�����?3T+9�7���s�x��2�81�ѫ�8˲Q�����u�p������f���1�k�,pY�pI#��H�0ut���-�l�_�����j����4��	*B�;k�G�!��*�r��S+�В�wB��Z�f��� ���i�Y��v�U��ei�O߲t7u�ÁY��˼��$]I�������I�Iݼ�����".5(�@C��X���\8���@}S5�N̫-^]�n�b���V�@|���Ȇ�>����Y�H)�Z�n�6e1ARJ����&F>G�}3Щo�p�?< ���(��6&G=����d|Lx������WH�����\��{��$�^�v�Nճj�"���mꬰ4j�af�Ȥ m�vR�I��,-S˒hFv�B1��I�����eƞ�F��������y�k�k��Y%��ɘ*x����7@-{G�#�����#xmP:x�&�m���E�\S{w$�U�3��O� ���!z��X�<ﯝ(a�I���"a��Kۿ��0Y����)jU�U=��ե"7^ޣ�А3�"z���^��ף=��`��ā���v�a�B���o��J雽����E6Q�k&$�����1��Sj�\e-ʘ�9ޒ��w8��'�M��Ca5�p�he�]��#�d|�d(r��6����o�	?�Y.lH�#]�?����`�3����䊧;��� �M��x�w�x���f������E��9M6g�;�s-^�W�*̙�-9��
dv��/?s^sKF�-�M&̴��$i�U�ی��YxA������>~�V�Ȩ%��]|&��Q�� �;]ol��e��h���5m�~~����o� V7���7�D�nڒ�	��ɲ������۲V"���C�tZK�:.������
��oh����y�l�� ,����"�*�b&�6 r�3����2ʕ�=*�--~a�\�OK��.�ޭ�%*���>�o�6��w��6i��h?�/KT翫T�jnmMJ<�H��b�?:����Z��o��>\'��zR J���rs�"	�����}���	&}�ګ�,?�8d�=Zc@*�JKY'�e��OF~F�gn��(D�;�hTf�e�iS۷2�p��:�x������#�e�A7N%e𶄔�d���?�f����жڇpy�8�9~��M
T�cFG�$��
l����c�A!�ӓ�k�\�	<B�TM��Έ�y�$�n����\�Ҧ�����(�n��,��44)���̚����l��ЖW~��,��%@�	!Uh+T9���U�!��ԛt�H�n�F���t1�n:a`9[I���D蠰���V�U��|x@�g�w�Ĩ	P
-�i�xɂbR��UlK�p��F�Ǆ�u��ꘪiWȿPW#�š�v�O��8�Ģ\��K������8Ae��}t�-"X��<d�W�Me���[U w�ii0��9�����A��	�K4LZ�`Q��#leߟ�;&I����]հ1?)ƽ:f2��7�ۑ�`_���E\r�ȑ��$��������t�ư��í�`��t�V�*�v��QQb2�L��ޅ�q��"Э�2�e����->�}�#[���(�\k۩<��4�۽��)��E�hj�����4dz�dJ`�)�~�=	d�7��Ty��Mzʝ����˺B�i��N�+�޸�r��0�]X�<_Wo�q�sxӸ��=.��&��2����0p����l^O�+g2�������h��Ö�H��uZ$p�H�W;S�X�6F-K�/��
m���#u�_ú��zN�]��ޡ}�JX�qe�S]aP�h���,k
����q�u��fZ�/o�:!I�l�6�����v�c�M�ѠGͶs^�NH��}�`��5�;���Ń��HX�P�;�g���l����6�����L�h?b���`��X��O0�M�����jjS k�U���׀����S�p�o=��|)�Q�*(E�ډ��D!8�4Z]�&��t�Nq�9	6,���y����<���[`�䬲Su�Pݤ��Î��\;���R���4��7�U��E�'��J_N������dqo���,'��7�/;�O�<�ӋY���Ѿ	��Z�l�>Ԟ�'�<S�9��,G �B����yh�yb����X(�`T�bG$�%^q�F ��iaF������X��؉1l�V�@��7�oeH�%�Z����JeLr�qe�`L�EbhJ_>o�����J�'pչ��8$�_�Q'���J���%4U�.�T���L������1C�{:��9�z0�<ȧrUt2�F�
U��r�������z�%�m������%��}E� 1���U�)�R�Z �j�Z�QD��\�x-�a%�s�%7�]9⑔�߈6nʽϤ�!�P�3W���b	��.���g<����%S��k�4��_��=[�X�~
��$L�18 =�"�X���E�^.r�������_�-�n�7����-�ۍ���e��q�s�()�����B�fc=��,?`�N+K�S/�gp�$�f��⽕�&����BR��0ƌ�l�eO��ϣ�J����\:A�L�ݍNpR�q��tM���/��@wT~�,n3��Ds��5� �k��[�[��׾��C����Ns�~�I���K�(��!���5�ʍ�ݮ3M31��Z�ņ��Ji�MA�&;�I���`�*UzJ�"����s ��ƛ &��gS/�$�S��?S��^����I*�.����CF�>-��t4���n^�;G��-���W����~��V�Pt��3�r�cEo����l��E�O,1�����aN�)�%�G��=D�֬�"���B�+𡬹�+��>bo���G gk?+��®���P��*r/T�`/�RH!�zL2�1=��\nml9��Zq��Cbs�(/��V��ސ|Ӿ��q3�SbH��^�X^��i��LܭH�������g���� �/C�0��S. �F��X��y��j,Zn"��ZDw��b��fM�y���3k���
?���d�&�:��d˰�jwO5��� 8F̼G$�H�C�S��٩c�1�!��)]sɺJ�Ѫ� ���n��� �B?�$���i��(��F�bs����)��{�v�"
��M� �q��1 :��_�K��c�V@M�$*��:�j���0�V�FRK���79r{�GĖ�w���6�i�{�6��aׂ��4T+��&8�V2UE'���*�J(�9:U�b��k��5</�-.���]߸GPH�1L�(k�ƿZ5O]�*-KC�z_�@�;Է�˫�cB��+2+�E�<�ۢ�38_)2���0^��_��2�#�,�������C�A�u�\�x�:�ç�ϝ6�P�V���=%��NZ�M�%r��5t΄
��������m�ȗ��t'�-azX�BU �rKj��m,�q���[����L�E�X�t�-�Ud���~NV��U5�elw�D=�E|�(E��D�3A(1�n�����2���7������o�Jv���kw���2�'Y`�Z@�>�1�mp�_ �T@�(�9+J����7Æn�`�&��M���J^��kA����{�2B����A:P�h��00C����(���6���Ags�5��W�V�3�Q����Z���^������y
9�20��R��~G-~��K�R	d�h֒��J�s�dVɬ���B:�2��2VƏ�)Owu�|�}.t#�ei�������(v�k�o�����}�5��𤋮R��s�"�K<th��3\\�u@�-�7�;H�[�}� ��W�Ϸ��ރ��5�y)�aE^��h)�<3�]P�jJ� c����1�d��D�ʕ���$R8� տ�˥XS����=��[��D���k��Jp>h�Em;��B���qpi���oF*�{�2k��� �������ê垢�%J�κ�aP�Ǚ"W\ɔI|ԕd�[��GVt'ؖ7
Z}�=.I��\�O�#vYder\fk�*O"$��y�%��z����$S	�6$�xάݑ*�{�q�RʭLiuSkͅ��\����W�3\��>���\ag4ho7��;�ڦ��w^���{� �=�� gUջEn�J��$�!5�+V<*�/;�
�f�3ض��X�Hv_}.�c-��ȜM����
|�Y�s����p�>y|�!��Dl;Fu+�.���C�7 O�L�P�i�(<GK T6�>��Qz�ښ�8j}�!��t)/A&af�+M�n�8%�R{G��I89������M)��u((]�wvV�H����_�i̡�GATP�1��F;ѷm}L:9ȒE7��Iaެ��:`�-oR�7]8$�*	��~"F�̸��)�@>�L�E��;�"R��
�0�^TC�~��$��o?tw�$S`z�p`"E�a5��"�x������c������Z��f[w7.��C��5�gp�L�*�&����� 뫄q�Y,�D�?��KBo�g@pk1�-A�aT�������s]��m�Z��)�7�&�R��ø3?�� =9}��i�<��Z��<��06���4�w�C}k�`'l�y0��n���"�}�v���y���x���~]�[�O>����6���W`~ �]?�¬��F1A����_m�!���[�2�Mf��L��������*�;�5}�����`�!��zZJn��w]'��Z@������A(���9%�y���GVaL�]��K�rGs�����3��c�����}2u'��7ot���h� .�|���$z;���]|����i�Jt�\���Pk9AM�.�|^�?�Ĉ�L����T&��9�s�^+�E�,��Pv�u#����gpl��F�A@Q�zf'2��]Ī^��x�0'
+�]dӐ�r������7k"��B\<)��c���o
j��~��_y��ʊݼ�����XDLp^QVlL�h_P����O�,S<��2��{l�OQ� ���3���0�t�3=��6�[��? ���u�C���5����{�D��>[za����9�z/1�O{2��O�S&��J�����Y0��5�j ��]i�������XH�%��L�uɊ���B%aԱ�������)������ WY�%�3�(���>�;yy�yj�r��u��L�A`5#q��c+��x�%��:Y"��78�X�)��������Mqә���q��qO�Z�]���ϧ�k��-��?����c�X���ܪb��l��9\Lɞ� �F��!�m�ň�1;�sj�_���#>EՖΐU#m��Cn�/���2'^��ź$��� �7�=n�O����y
��+ ڗd�
\P�ک@m��zELq�Vg���N�쓔�Ik\�X���%zJ�1m�)��M�u*�R3���ٜӤ����@`q�������3�X"�PK���
�e+��0�яF�݁���7<�K.�c�&��fRGxT�)h?���7*,3�E��vj=�D�,������5�k[x}��ҩ�5K�&|�--2�̠�B�S�p<�k\N��qf�#����:.^�18�`|df�EV�Lo� �����;���Bn,
�5Ji��ي܃%���ՠ���"ߝcy�"�N��宼>1�_ei]^�vQT�Z֤A��K�z���S ٌ�%�$����]���	�d�Fo�����1��2��D5�w׽5\uO �:��}j�6P�3���j��E�yp�q�a+�6�Ĕ�s؂��!�Z�'�
2Պck"�K���E�@����=1���K�H�!3�mWJ+�e�g/;(��%�H��AiU������b�"Ձ��"�z�D��lP�*�ղ�I<�2�5w��Xs�Al
�_���Woзʪ�w��,|�d-���>��WJp�BbeC[�L�)��q����L?ev���2R~���`�F�s4�|4�`�sH�(]�3��;��ھ��ve�!T���'��Az)����:��l��%�'zE���������g��X
{O	��r�\
;C��!�v�e��"ߴZ���ڝM�>��F�6�e����~r!Q�����o|@�n�����,ZLb|���|��Ӫ{n��c�C�J[��Rz͸&����3T�7F�ue� #6��٨�91�I@��M�6������	;��cp�b#�6�어�c��a�e��W�'~i����*$P�H�}��N͑��URqh�i�ށ��r6~	������]���,/��o�#D�UiI3��dWj�^�e�N�D���6EG=$r�@�"��5v��3Kױ���2դcz�J~�hjRLS�=���T��&�u�h��b�"s^W��&��$�Ƽv� @z�AM:{iC襽�Q�wͽZ��ʝ(�hXR����7�V�G�SA��V_ԣf�<�q�gD쾖!��K��>���BTL�my�~_0�D�	64Z[��K-���]�ye�	���� %5r�`
8Њ����o_�����v`�X��֩��iA�-�8;������U��H3j+���Q�c���~;R�����YWԙ;�i#g�R���bѐůt���$��.*R;��*TM ��}�̫cꌌ�#���·���!�Iꫫ�&�|�8G��;����'��S�y֚n<���վ^��`��Y43�"jδ,�-���m��xI��A{���<��D�:��)�NmE��UX��J���2��o�<I�X�P��Z�z��(���>���E伫-��t9�/��Yؼ���.XQwR�UG���B�5��!��#�z�b��}����_5��xR�'��1FL�U��q��rQ�β������5g�<\�}u�}�<�z�jh�*/7�b�T��E��J���N6��:Q\F���D�0i'A+7���"{�>��y�IȧY[�Mzp�f_.A��I;2ނ�4�=5�}V��AX͑����H
�-�%�KV� ����CR���gR=ϕ���
���8�BF�G͜=.nؽ���<���aצ̵Ex���};�
!ˏ�Vx��-*�� �S0/su���n
a8-1�+��؀��v0��@"�ҴB%����NŸ��L�p�����'-s���G9Q��x�2��n{�����Q������杦qL�F!*Cn��9���j�����仠p�v���>[4�~�q��U���;0��@�?�n��ȋ�0��ϟ��r:��&��F�����z����	w��%�̤-���kh-I�b����l�]�dm���V,~
}��Ɂ7[<6A�7�WU>�.y�8�H�?��|pG����3�iݝ�[���;+ H��QH4܏�����̙Ӛ����ά�>�>B��.�N��:дy�n�J���Jג{��֯�\dz�d�f�~���"A�@R�3cldԺtk�8ʓ܍%�:[�-5�]_���pv��T�`��/�24@�yxX�p|wmp�v�`��]<�y7p��>t\�5�|ɊX��x-���|[F�\�2N	x���Ѐsw��mL��!ɑ��t�(_��?v>%ȃ2i-����4ŋ���������R0��^<v�%+CΨm�C(�$Er(@���L|]0^���H�1�o�����@���/�5���+��a��.6]������1����f��I�\}^��-b`�j�j\U���,,6k�j���f!#������2�Պ m͢=��}Vf�%�%]7����X6�R�H�y{�	T¤�@��I�=r ����"/�	�|v���J#���X�.qrWa]�S���_���G�N`C��Z�L>�rs���s�up�ƺ��c�3��ی���9ÌZ�<�)�?�"�]��g�2��^2ٯ�z���#�*^�7�!,��2��Wxb�y��t?T#��� ��^�y�!�"l�~���/�Ԓz��2Q��
��0����F6z~�ڜ�]r����@���,�s���.-�3�	}X4�Ɋ!��G�M�y �V(\-
�X�p�'�C�>7@�X���s���Jq���rX�Yw^!�����w�1�SM�P�&�DW顩�М��A+v<����n�)�F�j�<�yg^Q�d�	����8:W�.��{�� �0Pˤ��Ǜ=Nj��zq�x9��9T+�� 'z���)û���P�X�RH��A�f�Pם|&�x��W> ��G\f�Cj}���{��(�� �l �p�-�q�.ѮF�B�h�c`��7Ibj�OI@�T� �}�\2�/����c�#��5@��bnIa�f�_�K{nT�����燴�3��h�S�{g�pzP�:f����5�ߋ	��G�_��4��g�6Z���[�<,Ǝ��DK&/���ikP���`i)i�0L-B��H�6Tg��-4j�ۥ��P�e��@��%*Ef
��V���&W�� �)����eN�	�%!M�ˠI!Y��-����V�b`O�$�RcnR�&�C�bp�29F��0�޵�+��т!�{i�A3wU��t��:��%uF�c�AJ5�����[,ܻKs��kH��0���:��¨�/����b[17����(Nة�M0��ytI��3�H ��1
�wE-\�Q�lTF���G������u�:%� >oq�["{3�_q%��v����K ��gu%Tג��K��eS@��Ö�5��D����c���0��OS� ����P������:�Q��Փ���#���7h�e#Ǐ޻�e/�@�FV��>dVCN�-5-�EiZ����xCh8b.p��OUر��>�����Su�d
� ��G���3DDG`񋏦-`���� �
C�UN�2Ʉ���:��9�Gѥ���"���IXs+����A&J���֕���ãά�X�4�X(%GW{����)'�Z`�a�����p=�^�Wyd]D̛kxN�J�?��:�z�N28�93��EZ�%��!��P�<~|"�TԧA@1Dܳ��jէ�(����K̯�(/g�n��������{�L֘	�G�ڛo-��s��N��FT���s�I��HÙm�q4�*')��G#3'��k*�4�DR;I�z���vu�ͽo�t1��qYLҙ���w�~f��bk��m͍15  �	�
�v�驺R�,ޜR�w����V�%�;�d�U2��ilr�����v~wg�Sz�b���4�??~��)�O��#�d��_���聍2����\��;�c� ����+B�n�=iC��3��ң�<�U�̸V�����Z��{���p�e���ǐ��^�/ _4�2�~�Z]%6N�#?�j�G&�J��u24�3z< �5X����)���\��<�N�^l<BY���$7N���O&��|�9t�����~�j|ҝ9q��o�������$�-�u_�{_�  �Iw�rJ�ronsذ���^f �N�P�� ���/2���-ё��+� ���DZX"j�N�;P�	���s<�(�W��5��Jp�KK9c7�ىu���~��H�7`dh�W�ֽ������!x "�Z�a�jq4���Z��ix���L���*f@ǘ�^��aڻ{J�ф][O�u�`���_V�%��9z`\���[��\��'tn�� S������M8�9xZ��ÅƨDBi�e����k
�v3�G�����e	��~���~"�Ը��;��C��Y��q���a���aנ8?'=�!J.b� $b�u�_a�8>N&�a�w��`�9|\RF��s������-���ɀ끐�fk�I\�gd.��+�	��D��T�7Vc�RWʠ�@L������}
Tem){�.͒�t�M0�y.�%�Fi����֖R�$�m��h]u?��aSy��Ԥ0�3��VA�2�R�zr����A %��Y4Cߠ�m�,J �~!{ܤ�/i⏎�'��=��,�=1l��%,��6#��r�?��Uu�7��=Fo��]I��<O06�(zMx#������4'����{�~Au�����Tl���������<�# '��$l�T&�!�0@�틀y�k�5��wT�oѩ���n�eW�;o�/^��i�JAo�򐮾C,�[Y�g�fFB's�]$�'#�Uo��C���"J�~o���FLP�3iÛME�ʰ�u6%"X�mD>&�N�5#�ۮ���\�\�5����P؇my�)�-DJf����&����!W��҃b�I�H_�AjA��;Z�C}!��`�|���*C���	�Vϋ�O���c.�;�Յ��Ow���r7�=��N')H�d�n�P�p�q���?����ݾ)¸�Z�i���:ܱ����Ƞ �_߾�Ͼ�xXQ�ߐ`�������^mS��E�d����e��{T��Y��X�C��P�"����0r ll��	q~�e�c�;ᅁ����{xDS���ܸR8����K��C��#�f6��}�L؇�?�r��xO�����{�^I������:}�+d�rՂm2n/��Qڡ��T�t�m6Qi�%=��j,�󩸰W���@��hߪi&���Z8�eٓ�<CŔRg���ZQ����(�w��3JD��\�Q�OH�ᏋǼ��O�m����ݲ�
�Wym�Z:4l�g��͙zH\�.,��8�8F;S�Trs7�n
r���_�S���8"`)�1�̥M����Q�ߢ�J��O>���x���T�A4���̘�؇2��"(���e��������l�&��'��Q�Ђ�9I��������Y�ű��1?'c+S��	����I� ���/^d�g�+ڛ��9�w�"���� t���t3��;�?�ٜ�!dWw®!��	��~�J&&p���)�j����>�~���s�ox�@��[Dw�6g��K��}�V1�rt�(|̾L%�v�i���"�5�(��*:�n4_<��#O b#�]vL9n~�*�7Dk�]h��p������A/al���r�����!	����$@�]|&uDW����2O�F�"�)>�"'MgxD�=���d_���ϸ�ׁ���F���j�)���(*�}ή��<�RW�`�+hq�]��[�)T|(���e��[����	>�NP�q2a����×܋'�*l@*Q� �o��K[sY�K��%��x�6ވ$M��v����8��Dn���pA��x5���Kx�������5M8�!;:��2�Bܑ�YX�e �.o�W?��G�l���F��Ǵ�KCx�y*� ���"E0W��i���t���uߚ�O���\�~�q��#=�9��5)1�"�7���Z�b��tn�<&l�,��gh_l	�$�b�u�4Gka���ꖖŻ`�P�7b)tbƭ��<�sM9vaW-n%r�l�A�:�i�R�y|���*(�ʂ�&��13�op`|S�K`�J�Y��c2�{U�'[hWiv%I�U#��yV4��:;G/�%ţA�����gҡhi�D/4_�+��H�O�4��e)!u�r�A�j�M��a��;�!���V����5�,,({��qb���1�j�1=��E.�'S����*i#1�CՑ���I�=�6� �
���U����H���L�/�,��X?̾+z!s�wD^��𘤔`�@Y>����j������ŷYkھ��/f�-�&}����P�� �Y�F�!��Z�c;7���5�&��Z��9�	�qf��"@�Ӗ��>�%�Fh�:<!=�c�M(�v3q֮�y'�7������ve��z�����(PW��˼����J���nMSZE���x�kƹ˪��A��������xwB4I��UL}�sH�~8�4'u(U���x�v�'�P�\J��Y��,���Ǘi��?�;%�U�.?�G(�>[�DBQ�~�2=��e�%�8�S�@6�O���+����	o8a�
�.k���#|�K٤�8;�0ݶ�ս5gL�Y��A���k߼�\u@P��h�B���Pcݍ�4� M%�W�C �Y��˿}�����x$|��Y[��p�
��HIy���P�a�l�?�>��o 捫/(�$۠�MeFͪ�s~�m���>�X��b���h�ѯ�J�Z�ad�_���lᨦ��Q���$��G��o&5���Ѳq��KN;.Opc�-#�1:E�^�v/���i��
'�����K�i�����<�Hf�S$FH�qüL�	���i�U��7��`\r�l�=\��yu���5Մ���� ���^7�����2�=�ʅJ�ȁ���Zb*�� -�0��Vٔ�-���Sc-��;lV$�-!d���-�i	���3i�cnj/{��_0ͩ�=a�����8D�'^���e��!ȡƷ�3
��c"`����w�g �	�+)a#���w�o�r�Ed�3J��K*j"��}Z�6R�t\yH��X��`�c���䜁�����I%sղ�˾��u5���K鎷� ���X�����Z��ĺ�x��N����$�ٔ�?�Ǖ�qݴ�0��W�;�u� �zu2�$����00����0u��e��g3����oP�J�J��sLz���O����,�s¶�R�g��͂��< �Ǵ�;��4q�'��si�M�Xզ�*k�=��,�zp�J%m �l�ϱ$k;��s�$苋Qއ|�������~{�Xᓰp ,=j{�'�i��ll��嗟�OE���"�'�;f�Cd@� �x<����ۭ%D.��\�UT=h��z���HZ��<�a�i��9�s��%�W���o����b� ���R�U{������������}V�j�'eP ׾u`%l�_��,?�X��P0�4[� � qX[]�y�&���W�3(���rZ�D�J�a�Qa(�Pc����:Cd��݄�`��!.�O�������i�����m	���)��gֻɼ��߉̤J�ÖW"fwS��Qz֤qS�2�Ma���Y]!�N�c��K�J&HyxKR��o�B�*�7�j���s]�y٥�
Q4��T�O��(�X�G�UU��$k���S��٥���;�6����x����W�D���-�*�Y��]y������KZ��:T>�CY��F\�p'`R�Zo��|$ce��n�&�s^W@��h-m�0^rl�+Z���>(���vϑs�'w\hs�[��ﲶ�G(�8bBoL����W�I�hʥ_�pC�S�"Z�.�����((�]�����vx_8?�l���)�OP봗"*"ˠ��ʰ	�F�f��?n(
�L��Ճ�pq%3�h�X���p�f�@<\�JL�gF���ѱI�_o�Q��x͐�f�Xz����,^��!Nu h:T��o��6��ZN�j�����%���Q�)��%%��7�����}#?�j�y��t��rE���Ѫ�c]q�@>���yW!�����5��3-��XN�ݿXȗާ\`��f����Z���)��z�؋�9�,!�Z	�1$�f.:������{�ql����>���|c�kc��A����:�H���0)D������ἧs��I��5V��SZ&%��9�Q��w���ep8�D��M�Q��#.�k^�e�cXT ��hɫ�مH��.��$6���/�2�m����v,Y�]BbP��`��@���:"�zsea��{"��(�P� ��*��n<��,����`h!��-Ћ�h�p���{Z�f��2)�q�d�c�m^0
�YDm`B<�ho�/Z��F��2�e?��]�7i%��t--"C��7�3�%�������åv�:�Q��_����{�lz�Ew��lS��2�X��T��1:�����_����w�5�	b:�%<�Jz�}~�N�G*)�buo9r{�`FA���ޅ���pu�%�޳/M~wzR���,a;�$]4�D�p�Z=3�����R��ƌ{�����	G�Ek(� ��1��KG��������~Q��=���V^�w�ERL��~��?	��M�F�Q�xq�Eہ5N�b��q�փ��&:��ߡ��ߡ���c-�͟]^�8d��z�j�w/�}R�|��6i߾����"�(c3������<$&��׹f��T��n�j���<��R<P܌}i� �����>p=���6L��������u�����E����k��-Հ�r����	e�0�U�XD��Θll��	�����=R��ó�ۆ��˦ NL���%�վ��az�.�'�B1�H&7�i�s���|��"s��ڟ�!���_0�&��p�?�cN�Uυ."�	8�n�|6t��&v�t�,RIҪ�bNg�;o4+D��PF���m3���EQ� ���!��ߠ�BO��Ez���6i�Y��%���CI+�Y�1Z����? W![��_�,�Zs��gˤ�A:���=1[	����,�M��[{��OK$��Y Crl���1-����P�_1>�x�z�[�sE8����|��9����Y�ؓA v-�
8ua<{3�)��$��g�	,H!m���Jc��/1�� �*V�e���OH&ڲUu�@�������.��%�!�Ⴔ����ZjJQGcR�_�s�7�X�p��d�\�|¦�#���D-5L��53�P�\\y�^gW(�_�&�������Je�"|7?�1��{�\$���J����Ic:�a�I�}����L��#�g������^%#4�6�DE����'Ĺ��P���]���HR�!FH
i}��s���/���T�>>��g�l�Cı��݀��v��M2)4���>���}�}6����]d[}Ʊ��g�bj�]÷y��~|:�Q<�����x��hv��a�M��aw�/������ȟ;�t�U`�xSR��O2�f�r>�T���N~u	���-���6u��� Y?4���r=
�9�;Hp�}����� �Cj�����b���6{�M��7"F&;���7�U>�O�����#��!g�ٚk�8q/�2�4*�p�uj����%��O<i^ٜc�6U�z��[F�	��<8���ʭ���"6�}B�'ry��s;���J�-�׍�yp���JR��>3�X/�c<]�܂��I~lÏ��M~
+j�Ä�S���x1=�����aV#��!z%�c��_W+Ǆd�u�Rh1br�� A>�֎��7j�׭4��9�:8�OMV(�Eq[��4� 6c~E8z�NՂ�SMAr�b�>W������tt"���v�5����Ǿ�V&���t&�����	M_joUK9;�PxYg)�L���s�)aj_��Д+V��?q���XBǝˈ���rL>�Q���75�g<�䊠mQgf�Dt�7�TrM��ԟyN�U�vZ#{�2���(�!�)� +,�/8_��ZV��O��$��&pU�gYZ�3mM�z�<yJ��BOו�L���������)����&�T���6Cd���A�(���^ZZ��r�p�!���x|�i.�/i3��e�3�7�-��?,gk�t�s�}�����e@����z�	6��Zt)j�i���{u������C`Z��I�˝񁰢3~������! �r���{��� y��it�Xi��^�%m;��L+JnH�{k�-.��%`�w� ��~.c�!�q��'��i%�hXI=��mci~ov[Skh;�H_��m�<��,谖��Rab1�Ac.�'� ��WQ� z0)��	��@��R�%�q�p�{���� �:��?U�oT�U��z��:d�*�q*�s�C
�񼟩����'�Hc z�Ҝu9Z�B^��y�B���+��"��h�E^Q���Y��HLt�IV~�I'#�/��Bu�z�*���n����y�W��H�t�B���js����%��c]F�hG�x�Ap2�Y�A�`B=�[a�)���s�]�3��W�MA�Mӑd%O�X�WBkX%��Efo:��"yx���E�^���67�k�Hm�)]w)J�:p3���sgjP�5�x�$ &8��1�����xRx�>�f��u%'�d��Z�`�%04���s"x�������[�)�p���w��۬�67:I����L^t�C���l�:��:��@�LD�	'�a�3V�zCYIi�qH�[��PT�k�Yz�KF�c�s�,fx�z~��."q4�2�Fn��9����=v��k���X�4�w�U/歟2'�U�A(���Z��G���9T� dg�r:L|�ۛ��'%;�^�:�{�jq1��G��b��!�)7E���_�~�W}��5�-�Dc(-����Ű��\wO_��"]*!C8raQ�?�6��B�1� ����ֈ���D�(v�i�1?�0���n^����S~-d���z�X�d�V�vCx����
�4�����Q}��ΙUEYa�)�3H�]ý;?�m����7��;|���E�J6�E �m�4��}$��x��]#y\`�hp܂�.�"��T1jSD̤::$|�ww�]_�&�(��q������*50�g��Q2u\�f�^����H��,��e�*V�c
7��t������l�9��"�qBə�>]-�.�N�n��=���=�����q�<�^;W�<�P��	�Z����
Q޺>+;)�nE��(��[ʌ������}��R5�`Y#�la����z��8�z����׿�o�V�k�
��Jy�8#ȫ���D�1����Ύln&��ݔ<�ܫ^�	bǔC#S�g�<{��0<�re�_M�#jO�_-{����آ���iO���a]�c�|Ԙ���F}r��C��j�|I�$�y�?H;�K� T�ƣ[���F��q��p��!�FLS��<�	�r��V/�$��ܹ��VF���4��if��[X��5�sF{�G�'Z i䖁�{mH�N�T�v��K�~;���-������!ם�k���#��9V�Dg��s,������G5/�B�7��-e�ӡP��\<�7}��=Ȣ���ҘF	�̗����Kz�P�`��=�Г'��FA}�W4&���8x�R��;~X����a�����i��ݐ�|�����m����yh&n�¬�g����kֻ������V�/� �,�q�:>r���p�M�r�W���!/&G�
���6c9ѕ���Ѭ^K�g�Uk�q��kP�������E4 �,E�����lwH:��a8��;��r3T��s����{�p?C�XH���
�V�[���2��E$T(����Ν��+��+"��Ɛ�g�M$-%�$871�;�0���JR�P�C>�p�Q��aE�q�ү���������yy��T=F{L��l���V�\�Ώ��q��~���Ǘ���'�d��	�d��$�å�乲𚵩+�����C�V9�ϱ9b�ۀ�1蚰�Յy��N����dw�A��J��8w�_�M��K��n;$�Ew40�L�M/�j�>�?u� �=� ��M�jy6l�A�s�������1E��H_7��4T�O{U�mtF��Z�f�#nQ����}���4��b�-��\I�~�H�{H�H�Jٻ-��@(iq�Դ�6k]�6w�pʊ��+TO��'W�����n(j��[�/H$���ͱI�ޝR�$+��s��9�!�G�j^���)O������B��{0 ԝ�mS�n�Ѧ�.�]��'��Cڭ��7�Ӄh�v�cv�7 4�+�ݯ|M�bK�o\�W����y�-��&_C>���.�ڢ�ݨY���������g�g����i�j��ϝ!Ӄ#8��W~
x�k"~�mu)&��B�ֺ��/E���,F�N�9#�4��!��*z���� :�Ο���fe'�Ճ�~��^i��}�*��ZG�l�{PdY�����JK��,��T�ߌ�W��^���H�N<5UZ�<��d5�~V�@�YY�7�4�[���NA9���w���|X�O;��,�u�s����5������|ο��h=1�|R�I���Ĺ3�cH��vI��#�K:t?�'((�c�؁>�����a`Q�*,\�}5~�v���,g��k��Rc>�@�q����FN�Et�a��ah��Wn"��Ⱥ]��hں����w{�:�j�{��o���ɒ�ϑ(�\�V�1���.C�G9
��m|�p+2z�_(�wy�ǽ���S��f�Ҏz��4��+ab�g)����s�~�Q�^/Cً��ݯ$ݲC�T�P�Ӯ�<g0=���SW�	<�Ov��� /=^��釨o�_��PbX�c�,f�~MQ�GX:�Q�,���>���@y�؊��k{g"�t�p���OX��K�>vO�E�_�neϏ�6Ω;�p7G��V���x ���g�oJ�47;T��~��e؂�i']���Q����L�P��m�~�!�Ή����v�˂��Fۨ<�(5I	f�BH����2��&�c����%_$�~��nD]gm*�k�����ICm@(>v�.Y�ޓ|tҿ',�u�����o0����w܈9�vʁ�Z�%f|�z1��F���+p��=�������\�m�P_}�"��	"�W����m��hMC$7�w2�w��d��y&�l�u�p�@�i�1ib&�m2!��D�	S.S��M��������6v�#��P�P<U�Zc�7��Pߝ@ǜ��J��RX��U%!�_�j�˿��C}�J����U��c��F@k�Z1B%D�Ta�$O�0�狾[L�C%L��RW����l��26�U���=�C��?�?! ���R�*͖��.��T|m��M���b�_�dfi�� ����߾QM���T������ ��3����¼�-���;���X��`+��K�n�_���K�O9tg
�~SY�Q�5m4�ۆ��P�C�0O7��P�临ǎ�x��Adb��Ɩ��>-:��� ��eo����:�;.�
�U��Pb���yj6��5��..4���"��������W��b�F'�՚�zb�����>�h��>H��'v��a�%
(��\6��S��~y�h��K�[�ה��B��&0u҅��^֣�1�3�і].��!��h��2�:Zpܬ�nz� �d�V6I6M{��2=����F 	�XZ�j�������:���6��<�n6~�L�iM~�Գ�H%��Q��� ��U,��@����d���#��(�=kE�u�J���o���K�!ք��J��r���n�x��I�h�����S��'�'!|�����b��Cn\Q�m�_�\����*���=NRcT�u�����ZY:�h��p#���_��O铧D����!��{#��l��^�_A���V���Y2�ͩfC��x�V2)Q&`�8����������+�k"2]��R��jm�]H�oC6`���T;S\����{�͠�f*�τ��/f3��YS��v���H1j~9_bP��(U7�M��d�kZ���>���m�穐j��G�!j ��b�w�.h^Z�x��eQ�/��I�d�$)�*5#��%�1�y���jk�+��y
���.�K]9LT�����[�Fs���7`=����y��ذP��A�2;�e�?���e؅�"AA��T�9�R.�1M��m� EU�4�עsT��1r��X�z;�z���cw�b�Mg�����:�������>:��.3ōz_IԢ:/��y�ڲ�DM���!-�<��wG�I`A6� ,���ڠ-�[���:M'��Ae%ֽ�
��ݟ��Vm#�"Ӌ��H�\���S�Q��c�ʾ����n�>�5��\��z���V�d$�.������=@��b
���ȽVE��J1���o����� ƒHL�9`�ˣZ&ob�Hx�ZG������4�h��f��T)8N0��d%)[�ކ�c9�d}�(@�W<�~͏7���oD���N������߻" 03(衙���a��l?
'����^!q^�㗰��^�P7;M)ż��j�Ӳfs�z�&�ƶI9�B����`��8�B���4WAOu*ߠm�m�?r��2?u�KZ
E"���q��Zǧ���n�im�\:��;�����l�b��^��s�|0�M��q��\���i�w�������ׁܑ�}��D�>�O�hK��qȧgE&V���;�|D�(a��:#�&H͛\����s��K^j�Q�N��F��Й�Q�"��l*���JD���]���x*����`�rn���.�p)M�}�3$��'X�`=���i�L��G֌��ss����SR3&���H,[^Z�j���[��$$�����F�ci<���7�Z�����`�� 0�F͓R��+��eĵJ���$�ٴ�6�-��!l�������x߅I6��m+B��]��Bp^�i��,#\�Dx��������o�*WW.��|�����`�Ķ���<k��ѳ��;�o���P�yj������u&jD�������FE��_Z������P^����.��ͫJ;��s�S�H[͹�%Hs>"o㥅؟>��� ��wTGi�S�ԧ���[åk��piK:n��������L��Q�@Y��,�wi(�n+oBC�!O*�u�zY��ͯ�/ބz����Z���e�g�!Z.������a/�%+zgՉ1�=��ԁ�̡&+��w��!w���s*� �N�M���G�#S��]Wa�fh��Ɩ�ŋ��@#e���U�����K�W��Ba������)2�y�s��K;���=k :�%"��:&��)��θOY=W�]&U��L�/c��֨�l�>@�C��1�* :�݅A,,4i���Y����l_�)<��ʄ�0�o�Q
�#���~2��ZOM��f��ޝ1����J�"�|�gp/�^�t�{xVD%|?�QL�\��|���T}>�&���^���k�л�U^��&�pK���b�?�4���LCؖ��Ψ��R�T�%��\������BX�*u52���RE����GFeV�H������Ab��$��~w��Ѿ�s��f�_�����:����c���ph&�����0�v�9�AE��m�)�f�v���3������ǖO'����C>���}9)�w=.1w�/���c��=$�C~ɴ�o��4��X���Ss��~VEU�gs,F�8�VNܝ(�xjE�������0�����'h��2p��%�;c��5������F��+�G�y��J6����C�]�욇Vc��L$�&
Q�UX��ņ=��S˰���8�)�f_��D�����jE����|X{2BA] �h��FQNf��=��2�L�,���e��J(���a-� n�<������$���I�@|�|d�ƲB*#���j��?�.�+��8�ջ��|3�W�}9���u�.X;�rc�(͛�����B�>���/�O|�t�%«�{/�!X3�h����hr#F��4�}VD��\��kd(���+��E��J����<u�K���	P�5���ۦ�
�B�S����r�� IQ@�o��/�V�q8�ڶ��� ��ޢ�E!{N���͘O������~1Ã3���xOJ6�3hi��ϰE�x�>>��;���1�)/�v˯�%��r�Κ�NF��M�_hHM���-��q�L^?Dq��#���e�3vء��2>Ѭ��N��,>'_}��ϸ#�p,����9K>bB/��Z˒�"6�L�'�G#��Oh6	C2ĩB��S��>6Vk�Ń�G�fӯ�6	[�1#l(��mqY���d��3�N��Z<h�=h%  նI���H	VR��b7������N �(�9tp�S��K\��T��a
��b@K����,�!L�[�ɟ՜R'���f�2",4���˘� >Qѥ��xk\���Zc���裓�&߈�Na�
y�׾�z�� #�-^�G��E�)���iH�	��a85�lIPRGDÅF���0ғH��i�$���i[ ������,�GԚ�m�V��]Z?*#�0M�h�����2�J�������y��zq�8&���IH��ovg�Qo��W�\/�8p���҈��RӥB�4��^�k��e��x!�s�>.�5T�n�(Ȩ���.�D� �yO~��Sc5�����_��DN�����2®_�k�@�ʧ�$��wߣN��f�/#^��Vl�sx�6:J��5_�!�~�!VBB�'�^�;�֘�-oϰ�	�=8�f�ғ�4֜�b���]������	hQ�� V�jUʶ�嵴�6wV{�V��\�
��/�F$Z?���/^w��&��*eS��-ab)��i�.FyX���	�+�tz5����!�k���(�H޳���I�6�*��b^jW��ި��E����]��kM�u�0.�BE�$���Х��:S)*h�5���X�9��\jQ��"�`8�<�%yh��&O����%g��ҠL�zȈbq�D�7n4syF�c�{0���Q=���<19@�{㬗,*'�K��&�0A]����O>g7�HӮ�z�J��v��-'I�G�m`�5�w�)Y�y7J����ꬵ@I�9����@n���63��6�ۅ��ez�ȇ��u�QS��_vIXHy!��c�3�2f��jHD<�Ҡ�#�����[��)cJ��;ޥ�}��$xYW����G�*�������b
<@.8�ؚ�?��!�j*�����^),��fv<~"X/<�EH}�Rܑ��ecWmJ��\��C���d�L�/m���e�)��Bۗ��*�?�ʼD���N]�gq����)䕨]�7S���L���l�������/yQu��|��í�rݸ����:;��%���.E��_��7Bi��M��J��AA؜�(�2D����?������_�
���M�iul�~�ޙ�Yk,U�浕�l���B�ࠍV�&���Ԑ��9>L�D������烹c[��\93�Ef�̭�ῐ�+,�����!�מ�'��#��h�(�\������G��HHq;���x��ru�9(u�7�i�)qYՔ��'�)��"8ŷݬ>���j��SDH�>�� }�`wh���ҡ��bl��F�����-6�4�8��f����	_�iW�,�¿{������\�Y���8�dB�����.�Ʀ��\�V�� ��J���B�=94G����x��I�-ʓنM;0D��k��Kx��;�F
ٺC���d� �sr�r]-hD2�F!��.����1ٸSz�Yg��O��+��.?$���ل���[����Uf��?"h���1����/a�ʧ󩁀�gb�9y��vb��=���M�\�P��8?�ó���u��w��r�B�����I����pe�юd@���O,3�}����՝�{Mp"C�U!H������AV��p	��)�n]�}�/eKJ�y�A�;����bV ��t���h���[X߿��#X��}�>_��;���tG�ʏ�N�p�|^m5�u�8������b���E��E��d���>D���
��:���t��)��W~e�h��v�Z�?�~Wo0O����������q�!���A�+1g5t""=޿�p������)�$8j�w�#��M�I)�T��m������~	�[�c�١l��,$Lj^�'��(	�x\���_3����:����7�	ф�q�Z�
-f�(��?I�%Sp�N��B&�\�ST�X��5R���R6&�L]���	���v�"��Ta��ʰvTK֠����[(S�@&��}�ƵcQ�)7ƔF]�fBm�%i_	�aQW���[�-Z�ڔ.W*��^���� '+��K	Ly*.��:~Z��u��	Y)$���J.K#�+u!4���/K7( G�W��S�F���?�^�Mg���+�ۮ1Y�3+�д�H3�Ng��+��ę��R��e���4�Һ��p��������c6���;���$���_�rЩ���X����T�Sްp7ܭ� �~9B�6�tG����Y����>	�g�ڥV�1��y�`�@$����ti�{t�wE~<�PD����=G���r��mdؠ]�L�Sz����?/���M�
�� ������E��L�q;!� l��^��o�X��N���. j��P��c�əK��:�^����W�L���mҹHv裙\����5���?�!��M�s�ƅ�Tө�ې�{�(���\�A�'.@V��mM��ƎT�����i ��ŋ��D�JC(�j(��zL���F������wg���]��ӋWwɜ��m�ͧ���ƇtD�r��⓸+Φ@����)<�E��F�C����~�]H�m�vbl�Qad�x�X,d�-7������M�-qO��P}[�z� �R�پ;�8�)Id9�IGBZM�;Q�w��r���ٵ�fwH�%��0}��o���֐L扃4�4� �7�5�C�d^֣�8etS��w!ԸI���f�0
vflk�)����&�]�`�'me�;~�ͅ�j���|��{��I�"+4�Bb��%ѫj�Yl0A�Z�����L��"v�d�����5��%���_�+*����}����E��<�-R9��z(m�O�5� Y��:b2��A� �t��p�Î)߶������ı�bk�.�2j���WjY5���j�	�4�B�a�M�u8�c��8>�(�qS@�j�C���ATcY�M��T�&�a�	Gb(�z�]��NV��/��������T�W8�|#�{�����H�>��k���s�E ?I��%��*��~�ԕ�P��U#?�g:�d_����OA,�cL�����䄨���@~��M�`���z��JW*i�8҂���.���Vi�&m��e��=NV/�~pxl���礚׉݂H
� ���/�����M�����yc.�Q"υUYMejpN�\Brҁ2v�^�D`��WS:ʻ�&����n4�1�t狿��U�y�b��0#9���S<�q�:��f��;�խ��!�ߝݭ�_��זv6 ޏl�0���f�g{���L��M�]�xgZ���K��˩���������؉!+��.��5d�Շ)f�{���eΘG����pX��5��$�J�j�󴫜�b]�Y"S6�aI�0������`ؤ��o��	aXY�����rk�u��=��f �m�����&�f��LX�[̷��'���d��.c�H�1�B6�E�3�eR��^�^��xS7�d-Əp��Fx���t��YRjl��0�%@�UY���F�ED�~��W���-��qIHS���f9��QҖ�|V�q9�=���������s���4����c�ݰXˀ���|>�?�<��@��>���"�t�'+u]z^$�=#/�~�G��F{j!	��￝J��a�&�2�7T�t�KO���\�qJY�Ts��t�c)�@�19�㣷kC`k,� ��퉔9�<,�����)�0۪�f�h���B���ۄ�dB�r��iH=l�~��ʡRXe�H���p.����t�i\yS\'ZyiO�4���IOŚ�V��#��r��M ���To�?S�Z�A*�W��mc"I1v�^���#y��a"�ҧ��\�q��Eqk�6m�&�^P-ʴsd�Ҩj.�]X��y;6�`ܰ1��9���`�w���4���y�h�`���0�� }�O�󟴂1s�bnt^��Y����JTUR��Y=��i�d�׷��g��V��� �&��^l/ڄ�s�a��bc�}��3WZ�����s�LM�-���bIj�H�l�2gS¥�'ACˊ*����]���J�3>�P&�e����9o��	
�qM����q�,��ik�M$����euԐ�d���2��V N���tCfv�$X�6��^�{��sa0�ay�):l�s�XH�`��s.���4�l:VP�u3�|���ԥ�(N�*�Ά�M���~�y���!��8{pP?2ډ+[�o6��L��DL��&0C�u�	�=��������q��l��
>������`��a-���>��ݡ��:�=�PQ�;�Ṃ_eW���P���B���)�ǥ�˫��<����=UMC���zP_��D+A��H��0֌�������{�
������߉g�jt��H��\��E�nH1:�8PlS�Y�w�-�]z�oh�n7n�s	�8�ܕA�����+:_�ށ�	�?���/�rJt�>͏�76<�m���@%u��:��6H��4ɊW����*��*!�P���19!u>(��3��ڂHx�{�v"�`5K�.��~��4��6�e��>' is Z��o�1Ej��N��7%��]џ��t:�
�I��	�h<#�0�绱@ꉌ���3���zgZ�w�e��k×���ێ*롦 �n Wn-�N����b��?��fQV1 ��E�)�KS�����U�f���IY{p�U�)f�çxO�2�bǽ�u�1�w��o�~��}�w%�t��7F��}�y�(ѱO��GG������_	&�J�pi��B�4(��]�	˴�U�q~]��wkj{3o�}�ق�rg̇<���F6�MNRP�xф\�Q(�D4CE�4��^�ǡè��@$�7m��:U�u.�X�Kr����/�Z�3��%��A���#tԇ��^�گS��#�3M���O}k�@����
{n��QhJ�ͻ��|��>�7�ؓ�D��2(y���T4AY���IY�2��ݿVܻL]Gp����y�1�ؼ��H)�S�p�c�7�f�H��|�t�b9Ap�@��/�e��\/dܨ��.o�����h���+���X�m�	r�Q�`|��r�s��@��̇�|�1�]���ˀ��L7t�9�{ۮ�O�0l}�
�'��e�@���m�1�2w;��=�U�.-�Wm�Vg��r�"|�SqԔ�O�-��k#��W/��]���C4�:�� �8��>+��-nFq�B�Mrb�77����l��ϑ�CTq�XKy����,ņ�`�"���!X�����V��v�#9������X($N??�G[�g4�p�.i�h/;U�HeӔ��X�R���K�)�f�6����c����lr�oym��PS�<!���~�@���K�B���dPuQ��W|�Qo'�8����{�yl*_X����O@�8�$m?��+k3ر�hn��je�+�ge������(���`�a��5��چ���:d�}����vք�9��#��od
.\���@������Tr�{u/�Gwm~� </�ࡽo�F~��i;֕��w)2���W��K�+g�E�y��5��\B:fV��Ͱ���^�.Q͂<�T�+,I+B��~ɉu��֖��3A�c�I����9��-�/MP��,�_���4�6�Z���x�0
��j��z�����6��;�K��M��y��-��SR�p�G�(?��@Bí�d��=6���xK��n���P��(��_�)�New��+�܍h-r�&��Z��	��q�WO�����	m���V��Ɂ�APO4ǲ�@Fȯة�}�:�`RN\��6�d�$��nVU�[c�x9z�m
oV��Ef��B��X~�4A)۲\�O�*Z�U�RQ�>���p+�~���')���6�M���I��	��e��f:��`n���i{dw�4�t��شj�уO�Rd����?׬��Lý��-GFB�"{�eQ�Ĕ� 8ŵ�?	�k/�pu8F*b�t�Vg�Nn�������@짮�+m�j̃�m_��7��H���+��w4ő!>��N\�A'i@M���r4�m��45�]�qv���hnT��zk㟇ش�Q�w�դ��砒���T�F~�����`���m;��g�ErI�ZxP�&�B�x�L�p�d����1��}|�>�����.�)	W�"�'%H��H������ɵat���IS$�Џ&^3?z��{\���7�k�y"W嵑`^�g�ru �:l���n$����z�ͭ�=�C���F�����-/���b�^��0�I�O1�WA!������I���TEv>�ᝐ &1�H��Z��������&лB8�U��m����l��8����p�|�^�{�9*�s�m�A�2���z���� ��"�jvω�mp�j]?B1hJtsQ�Di4�k1��[9c"����Q�g�A=�8�F��X�뱥$����|E��OV��ĩ߫Suo�E�A}B��r5û�a����/�˙n�3!gų�`.ei%��	n�8�� C��J�h1}z��<�g�� R)52
ݩ;C�P>����6x�	n�<���nG�j�c/���2�ep�E�`�"��/XT4J��qgGW��0���������ޖ�t[�N�z�$��K{���>,K�FC�bB^Jx�O'���C�h޿m�����e��w��F<�����9��Dv�4p�x�~�7w�ğ!��i�W6<b ���^<f5/�9B.zj�$td��k�W�G795x,fd!�|��K�杰�*��w3��,����%]�m7Ao-S��w�9(��m+�����i޹ɒ2[E���E܇4Z���"�����\"J���f��R��O7��)��D��<�jS�������$���z����5�Y��6AmQ�SN�o�����>�%�8��4��4�[c�n[x���&��bI#`ږ��MHfǠ|]@�(�x]��A,�D��FpRQ�q�
���N��In#�mπ^��������[��6���*�
M/%�|Izn���-QR�M<����Ý�u�(��N�6��C�q�_����E�>l�nt���	��?��O���r��r�c������!��Z��
���������"�`�M�N��N!����ڶ�cfx��b���&[.4
7U@�(�2�~���}w�� ������b*Zd:L��Q6$���K����CD�|�Q*l
�[;�I���-Z`�"���9*�`��kKָ��z]W���5𾸀�v��id�~�k�*$��S�=�W�5�I[�2B�0ƪ��\���e�9��_C\oL�_�Z�o,�ݙl���>�j���Y�!���V��am�����1Y����^��J��̞�]3H#'6�
^�s�a��ᆌn�Gw-���!�|�$Bk��+̽z��v=�ҿ�����W��Y
���%�_�e�(1]�+Q�҂ �jJ�v������ b��#��n��b�|u��� "2+w`�����S��4�U3���աlD���"PT������ȃ$Vv;b}���m��S-�@9�:`8jn�d������⧛y����ٞH�I�2I���T��\����^�(�L���&�B#�5��]h�S��oe.�p~���K�b{`*� ��v�ؤ��r�hx�m䯣�K��X�R�p��~ad~�����_x�>��oI1R,Tw��qXF� ��U�M V�A���kfRMA3���#����������Ӯ6|�OR'�X���'5�^Ma^dy�4\ן%&��r���5Hy��m�D�+j�1��ֽ+���u7���fJ�t�Xnɕ��k�uԨ��|?�.�WѠR��X0��3��׬�g�?��6<�'�
4�h��I������A>z����I���"�.����z�u�2p8��a��f�IhfI"(l�#�E4� �3� >Dr���M�迡뻌��T��Y��Zt�u��=ƕ�&U`����a��ɮ���A�g� �&"]Ăf�z����g1 ���U%u��G���^��pb�w�����I�ț#�9���},
ʩ[�`�DpI��J��ѦV���.�Z_� �ѯ��gCP�%�^���ܱ4Vڜ�%/�4m�u�$�l�`R���S5��]���ƒI����N�nAp>��N[[�#�hC�(I2�y������G�T4�BtSn���#~r)'�4U�v���6h�_�2ZZv`�*a7ͪwR �(�̞o�r����wi����hɾ�י��hZ��/߽� ���9%�c�n���BRw��Qй<t�K(�_�f� ���߂4��HK��؞��hK�JEE�򃸬�ۙ@k�-J=��S���c���Ϗ�Ǭ��S�"����ҍ�����S�^�����-�u215��2�)�~�0�P��''\ʄ`ao�2�T��S^O�;�}�������v`�f\�{���Y�G��]�8�[.��*/f��|ְnc���Ƭ��τ�����rx�v�O�4��� �$Aq
��܁)�z�]&���XF�l�0�l|�"�>�
�֥�5��NЍ�;߃���e���"�p�j6X�}if&�]�K���� ӌucn�7�R_߫��ԙ��!��C�gN�9���������I����V�Z�=	��0{h�5 �X<`,f	��YV[$5^�����X��tB��:<��4��/���V])_T �Ob���ݎ~�*~�(��a,Gezn.���~2��ZS8$A#2�����|$�ܻ�����	@Y����a��%q�$�d�=8 [ZżJ�doj �l*��{���ַ�E"p	�ۓ<é�H�ކ�b��B��},���纅���7��AJ*(� SC@9�� �C��"���f6���@m���)��Zw
�Qă�9�1Ǳ�
ĚM�e���>��CY��S�پ	1��3{�5,D6�_�����]�����?��~���y&Z�yC�ժ�s���[��6��şXU��lH��j4����PI�������T�y }�$}���w��j����[k)���s�?WC?HM~��W��Tv��z����K;ōr��Ͳ���PrD��J�2C-��(�FǢW�\Q��}�M��3!	d�����g����Y+߇�{s���PW[i5�Ȍ��F�l(ar�rA��]�7w�R����R���	\�սu�X�wm�l;�6��V���W/�C����Qǎ�BPS�dX�h,D�bf�%&��?�܌2D�ϐz.w�6(%�4&z�����ۡ�����Y�>�L����y��lu7��x�ٮ8*~ ��54��"<�98�>=��".$��q؇��f�tu�[A�qZ�X�i�X3ju�Eb_2e8ֶ2N�9D�<a�8������`T��g��27H�o R*�9h,4|�;eLwe����	L�xn=�-˳��@���	�<��Ш��̥n�fo���2΁�6��� [�I/L;�ZF��EN�[�(����U��S���	x( ]Q!h���Q�����@;�q���uL����
�I�6�!�a�>o��e�IzAm��[)�������頋��.QZ�$����ٞ?c�m���v�˃j4��XL��L;޻�g�\���ײ�pr֢�Y��z�����������ƍ�5!�jP��#qX
�H�]��?h���XM1�,�Ѷ�n��z��:�徬[B�Ea��oր�M��p�֮S�ԮKo�Y|\�^�&&V�J�slO6.�d�"k��
�'Jŧ����F�`�-��j��1��:	���,N� l0���m�4�xk�������Fxw������G����J�p�1:�DQ��;U�m�b��щ�;�=���l����Z���Aʈu�ύ,�z~
�dO��Y�[<(l��V�_���u����D�Fg�[еj_3��������'��y�!�+.���K	��ct䄴DBT��]�ȕ5��������b.�*�p"#��nB(����D�-i��*c�u]OP�c�e�����)r+~9uG�:r�)"���F ����d���g�v<M"�#�B`jU��I���y����q�\������B�����z�c|���Q�X� dz��"�TiP[�+���4َ�V4��������ʎ�Q+�s�{���gos�Ԇp�܄�X��]�:J,�g�_Hи{Ȣ��c�O��� �3F�\�ol ���/�B��	&�D�jK �~z�{��nrM��� i�Că�y�C.�IUY���n64K���
蒹�P��$��V�����B5Q�u�+�N��p�R؁�N6��+ivR���M�H��1'��,�#�u&yV~�}�a��4nxګ����^�E��*������
mW��WXxS�fEr��r�~��K�f]kj���,���J,Ɏ�����{�3�' �އ�т���09��o�m�8���� �&"�ُ�J����`3B��$?�3LF#�`D�*������.*ht
�E�x�z0�.�%��_��`Y���O�"�{�y�8��G&"Df�<�6ٕ��|��&M$ƿ���A��V����E��u	�
�Z#;����I?h�5 ���p�I�r庆��B#_���6��]
g�/#1N���| �\�>��m�u����pѠ���.������ؖA�IBT��$:�e,'��N��R�=�p:��؀?1z<�7�i ���Y�ړu��]=��}G��,�
�Ȧ�3�_/��A7��F�_��s{=�Q-bx@���C0�����m�OA�&�@
�]t�#ұa5�̹�^�ۺ�j�y$��O��r�i���N��C�hܶ���/����EfG����soB*���?`�Γ\9�O�gXt��7k�3ʢ��r�ԱՀ���6,5-��"�<:,���B+k��#B��,�p�{|ڞX�Ԩ3��2 �9C�@᣺����6 ���c
���Q�[�k���@Է:g�ET���`�i����=��4=��P�G�S����IQ�ڒ �Dp�M~a�f8��tAs�� i�FݰXcs�S��T]r�" ��{� '���͌|S�i�	Ѭ�֙Y�����D�&G�]��[�BQͱ���}�9����j�<Wq��w}������a2-���,�ˌ�
hDX�6U��%�P%'`9k; ��^���G��}K�?X7�p�lI���g�X��C�$FFr��(��J��n��Z�YZ��>u=�yy��.}��`�őQ&�'W �M�����q5iQӰ}9��
����^E��������`ɇ9���8X\p��X�\/	�L�W"��fAR�[4����E쨃�g�I��~8&R�f\HZ�扟�~��R]O��c�h�sʼ���+����݃2{���,���fl�w�v=�V��}��1�F	������-��<%lV�p�n4[�5��vV�M s��/�h�an���\WHU��^W�����@���N���®���Z��sd���6���P�/<�o���G�|WʲVP����2�x4p��DM��ϳI)��Ut&ߵ�2�Kl�}��_g[��� Yk���Y5p���ޏv��H(�J�ݭ�r뤁�YNއ��s����Y�E����p�V�h@�*.2Ea����'���%���\�֯N�'�(�z|ȫt��@�<甓p'dtC�d�)q(���,d��_n6i�a�/���y3��swln�̑�����6T�N����'9�	Y+2�Ym�!�ٳp����#T�JTe���x`8jq\����:�Oo����� }u�e垎"@�������j� D*��o����R��]��Pn���E8:ٕ�*���tڌ�]�FϖN���-%�]�(2�KЗë|����@]a�QD�߂
SI犒)V��቏!Z�	a�"V�q5&ٚ|�h$g��KW�|�K��"J�xD��&l"��B1	JT���+'���=z'<�$�t���Y}��}��5G_:�!e��� �5Ǳ�wPKĊ�"�(KNN�i(�Pˇ'%@�4m���(�@��t@� p���x�W�vV|���U�Xw���Y��7H� a�ޞ�E{b������	���Q���	� �ݞ[�܉��0"��c&���T�H5�����hrc�%�%���;r�ʖ{Y#���M	�������O�����~w�ݗ� �&��|w�Z�Y��DAD@-wg7w�8jǰ|B(�B�/�̔�lf�Mp���}�`���i����u-Tx�=LI���G��H�-���7jCH�7n[��#��߮�O,�@銘�ޏn�eF�p�:o2�+�<A��Q�;Y�g�3����H���iAq���|&/\(�Kd6
aй��q��*�(Yai���@����4]20d����ӐׇR��/Tv�(֔�� D�9���A�	�^�Y�H�ڭ�ȣ`������BG�_wp�+�#�^�G!j�x��`x�d�c��U|<�宂�H[�����'(���9qn��Y^�>[J7��¹�������ǧ@�<B��Kу���a��h,������N*dRqQ}TV�W�{Si� �H�6D��x;�k��fl�h���hp�g2�zI\7�ԩ�1>�����	����v��o��h��Zg/�pM�0T���5�a�4lD}��Lv��k�ru��;�3t�.�p�&!lCVZ��G�b��G�_�\Wh���A�#���3�
��'b�	={>6���i��9~&eY����%��ZqEY�q^���[��P�V��Y�l�}��ĸ�,2I�/^�q�_��^J��f�SS��!.6������G+�.�P��iw�¢�����4������O���,)��xo�J�iʡ=#�0��c���_1s<�l��i�x����>��8�v��2$0���2����w�v��,��\�5�a�,��@�ݽ�%�Q��RW���W>̼�x�aWaC]Y�'�U{e�3F$�}��,IQ��Y _�מl{Z�M�6��꽡�"܇�F�/^�Y��G�U��w�	xx<'��|}q��XpG���gR֮�`�I�=���_���S�}���xY4�̑�s~����CV��JT��<!�9����dv���=�6���b�+b:Z:��mo�o�}T���2CҼ�&Z>������^p��R�%�^�+wky<�9On:�5��PP��~�M!4��tՏ���㒖���KZ���ܐ��Eo��
@�*�ڕڷ�t�r-5I��Q�@ߴ�j����%9/y�D�L�����+��"����s��ҙϨ;���jT,�������.f������1��];o�C�
�οӉ�Q��2�V�1�n%A��b��a<A�<&��� :��Bt'��$��1�j�+�{S܈�O<s�(�r0�,�`�;I��,�q��(�e��Qa%�s��YL�s��6�a.cq%I(����h�_ѽ; �*s���QD�DrVؐ�ҟ�|�H���Jx���K%v�n=�~1��HH᷏vz�z��R���5ť����w�Z �W����+Tp	Xznup�1����F(�ä�^����1�/��JKL�
Y�HS��F�yt�	`u�ïR�1��:ը��ܰ=����i�e�hS|z�Dr�l�k"I�{jl�B�fR7?VtH8�PJ��?I��P�XRm].X��C��ڨj
4SI���Y@�����^v5Y�@-?Nq9y֤�=�����_�"n��>���k��&�xm�h����L���N;m�֪��i\r�%{|�O���#U$�]���~��o��<"e��w)��6��L����"��pt� ��0�JM˾����Lժ�̠q��n��SNO���)�Vw�"9�ѷZ�s��u�������L% -��Ԇ~<�S��he#SO���~�����P���:Jb�4���7D.��/U���wv�eIX��_���9�@��J8^�p̈́��p��#�F��l۱�D{WD0������VN����!~�t�#���k�#]~��WM� 4�g�]�Ӗ��3��\�?n�OWh"������eӔ�����?/7F�QH�;�p���S�d*Evԋa���{d��myD�s��-�2�n�W��R��*���� ����K�@+}�� �9�~����jI*P�B&f���7'ѥ琟���c�$�@���`o�z��v*��4��fԒ��ns�'rGr/V�-F�= ^��<;���F��\��c̉\!n�>��3����iyI��e�T�ޯ��Ph;�xް��h4
}�/��B'�ޕ.�T�&BeyUP�4�ib��"��#�9j���%y�S#�ި ��{vk���Fp5��r�G~�r��;d
�^l���V�S��R��z/,��ԡ5gQ�!O�m���U2p�@�C��Wc|���uط�~��ώ��P�nQ*����:+���������))L9!�� 0���f�������͋'&�Ɣ�d2�F)z�^H�&�� �Sig
���N�B���בEZe��jV���EG/��7�(@Ϲ'���j�i�uaδa��,\Y_2��l�s���#�a���g�.��o��V��W��(W�X�ᆂ�I��e�T��!���jL�	°�v�7�ՍJ'sa�7���&��Tj/2��m$,���R˧�XwM�-��
w�^zI��df=ͼ_뙾��I��ݼ�}�"��>��lV��_��(��y9�@|RߦA�ђ�:���FM7�祀������H�g|"�dgĮ8a��:ʙ����,�$"=��
�H�2	y���	�~�#g���o��ϜL
`�5e�� �jd�'M�|0�~*�y{ov�*�p6K�F8I�Jֵ�`�I�]#�ܺ��Kp[��a�6??9��C{Ue���s�#ʣO��"�L��d�t�N�� ��}ߋC����9�������R��� ��[���ȀS��=�����j<Α�pD-��f˺L��Dz�o �-�VXS�W�ޭ�6dc��FP7� U�EwQ\����]���ȍO��2���n���_�Q��dً4���&�I�F{&�qȡ�O�D������\���p=�O��}�!����x�5y��>�̆g�p�Q���j�B���S�Z��ۑ)@���B�, &óȲK��R�
��u����3����?�Q�庹�f*�j����4=b�8��mM�õt@�8_�"-c��ʫ�"�^�βk����̢-w_Z���촑^�z� ��9/e� L��R+�!���!������v`�>���r�P!��u��#��>!��2����^~�|�]H��P�+X'����o���"��6*b�Uzܘ3����Z��p$1sgˠ< Ix率��݈5�ɛ ���!��+R>���`��5k�3fD��T���R&�F#WE������x��$61��g�RbL@�膌[b[�|������^��wo/��I�b�#�/u	��)!{��@U�%�����?�n�G�	26}�<B3i�bs6ۢ0���;�����5Q��p�7}���V�F1_�: ��M��\)�h���7��e�a�&�7M758�Wsd���+�#�@�Q�w<�H¦��Y+�<�9�T����a�����F�z8��=Қ:U]�V�?�V˭|?M2i�Տ�Nx�%����m���U��Smh1B'�b�R,J�6_b"N�v݇�S�߃���:�8Nr��~.��-?9�:�������^�v��^��gA�Oz������E@�[H ��t`q�4�k�!��c@�OS+���}�%�����W ��J���~U��r���o��Y��o�0�of��W�΍Y���T7�ꩵ���EoQҐ�]@>�u��`�U�IK��d7�9* CRk-�fI��?�=�&-G���f���@f:�B
��1��|#"�?��!�-�%���H��f?F���ǹ�@.�}U�Ղ�hB6xAY=�7��=�"o ��e��m�������h(�ei��Uj�1~�{/$!E<�d�fmV2���:y��3',��ܴ42}|�3����32Jr�}ſ��F��������0ϧ��%�.��na%g7 ����ܚ�j�H)z6�ТP����<>?z#Ä2��ޡ��{�.��%2:�^!�i�>%�W�;��Y�g�9MCsk�U���̿�ޒ����9��7;˼LmKx�����&�������qn���h1��8ǿ����5Q���{�$en�ҖU�|u��8��^��*4+B�E$5�ˀ�F�x�͜��4�c�G�]�1��r��cC+�A�̕�;�L�09/@5x~n�+{j3�S"���j��ԌG���nC1�t��g~2��خWk��x8��Y��޷��g�r�}ף�Zz8^����BۘWAv:��.�׌8��y!B1�^�����M����U� �.�\j�J�kH����OoR�P&C7}���aw�U�'����C���hrh����ΛT���Fv��x�nn��.xYc�v��[~����FD� #p&��&�N��8�|o���Ĉ}���oE���h�*�u�
h^5k�h��O��9vi�-�@�8k�b�~��<�mJ�4B6TZ����=`�<��Ɋ�m��'hg{�CS;7�g�A�q�\) �����:�ؽ�#(?�b�Ƒjpe���iE�0�G="�$�U�5�t���o���5eD,p�ɑ��(�=���<)���yp�g�y5R`�����%����5��)�{�R�8_��B-�{���şd�Ϯ|�tJT� ��Ş��ƈ!&� ��t����B���hN�ّڌ5*����`�z�=0���g��I���3&�4�MKX$�4V��r��-���{��J���G�?�����z�me ��鸗�i@N��n)�D��Y������t��{�0��w�"�C��@S�}}v6m�"�����;U�I�ۃs�`��T�FN�1o���@Xb�Ѓ5�s-A�+SΆ�޷mo/����-�੐�˓�:ш�=Pp|��h9�����;M�EP�T�Vŉ�p=꼛�D[���03����Y����S |0��̶D#�2<.1�:T��H��&�q�{5�,���A���J+�8U�X\� ��9�|oQ/�_>%m����x�_iP�e�6�E���*+�C6A�Ӈ�R1g�08�U�LLn�I^#��6��.4��?[�R75�T��*Ƥ
>����N�6�"ɔl2Ѓ���m9(z]ɢ4z�+�kU�J?�;'�j.��������x�|y�-��K�������V�JB랃��gJ=蚁�>q�2J*9��7������ �����	>ua��8ь�ކ�*�h&/��%Y��QW�Kpj��(	�ȯ��`2�Ԭe��ðv� S��L�(��+�4b�M�V�qA���@��U:��)#�6�N���uX�1de�����獃dZsjj�r�W�}7dwr���1���{5U��h��5��������`����q�#�6F�����i0�����s&��k��������u��������V|��˷	ze��bS=c�:���n�c�Er�o^f57�RM � �b5�o 7i�L�!8�����4?W�V��p�lk:�j]���]ᣉ�N�;�C�a���#V�u%�Bt�p]}�\n�������ͺ��R��ɮ�P��f�&%�����`��i?�]<(�s�`2�ߕ�њ\���0E�c��Ĉ{�c=)2mf�ک�1��\3�.��(Þk�."����,� �.h�*œ��|,���;�\��� �/�E �z>��	 �����\hC
�����)\�հ>��cA��:]�)�ș��:��O�L�#�~��1v�|�M�Z�6l�H��e�����U�Я�c�4@[��\b�e����.��b]:*H��p�{�a�Ϲ�5.	��y�������~��n���cY�~�T��dm$x�R��_���M� S(��[E+��`H�mZ����õ��z���S��>���W0d<'B.T���F z����UdN�V�ܩ"Ҝpq�y^�R8�jA.�J��'�?"
��@�z3(�z��_2�ڠ�9�v���q�f�I��U�;���g�<��2P��ڞ��[dPK���*�L�bT�|��k	Wnﺅ���8<��Tq�Z�oC�vK�~��M\Lp�p�(��ٺ�������{�+594�R�5e	�X(�#X���W�E3m?z)op��R����M�ߟ�i���'�~
�T��C '��Q^O�������N(Ĳ�����)3
.��u^0��y�"n���P>�wl]��w�pO[�x��<��M&�Io)LD@��ꎝ�u�f�%	~��smY+(�q��}W�_���nƫ��҉�� A������i,��Z�X�p7 �g��7o�:�DdPF�m2n�(Ԥ^>�+X~U�&��A����P�r� ���QHk]{��&�w#H�_�nJ5�F'��"7o�Iw��Cp!�>_���N�U��xH�"�XL7DID�x6�k�9��4#��[0����8�E7��G����	ՂTVC�ם�M�K���хM�>���"�}�4�v�{;�s�VA|X@�ps^\�M�� h$��9a.d>_ �j~�+[e�K��'����-��%�fT����&�QS��z�U8�	��58�\�j���ܡm�v>p�|���#��o�FG@��@]f\�h�����r5qe�PQ},���IA������Kt�m��W�l�[�A�j�B����V�z&8�;K�#���Ř4x8
���3�F��g�LU�<1���	���1=Y'T�i�#\�X�[��輤MoN�>�����-��r���ڞ������Ɋ�ô,��j��=��	'�c�@�KCc ���� =�n2�T����F7��B��̲=s^˘1��]uZ0)m�7��R��Ny�1J�V�����hT9� l�<7�FZ6%�Sy +��Ij)K��A�L��f[���@�o;�+�
-Y1M�:����}���c�~<�mg?�.��6&:�L��4G�R�0	��Mv�.�`���R�(4pwm�c<x����w������Sv�	����.�M�Ѧ�
���W	18=���|�F`�[~�-Ԓ'��2��M?����8:��d�DF�ϯ����٘�gR����˟\.�m�z9�����H�N7���B�3u�(�07��B�J2ݤ���+�QԴ5ƺl����Nicm>��M�.E�>�3Zp�<.�X�>�A��Bj^܇T���Yh�Z��c�Y��6��do����;�bZ�F�G�'��U��wd�xF����8-	�G7�~( `�宮̜|3>_ܦ5��3Td_��w���+����[��v�����+�A�N�6����G�蹨���>��_���	�xw�Y�� � ���Z��
_M�G�F�P��,?:b���㻠���1�
��BO��3�8��q��7fͫ��a��ʅ%�Ņ�sk�"~���w�i�O�� �I�Q��,����ah�Z{X>69w�-G���l�����7GyC�>k�U��j��(v���#ߞg�$�n��AO�o�|(�Ě���3
���%��]�!�+��܋c�4�{x��=m��!�98hs�]����a�ߓ��pxNп,���b�j	�?�؈���<���*X�o
��|ޥ�	�)���qYM7��!��b�g�okł�,i���@��'1sc��c�ʀ!m?W��4 R#�?Q��K��ZR`e�����I����BN`ٝy��*N���A�8o=lc�o� D'70cH�Km�H��Ew�G�a)����j���%�g�P�0�J�̈���ˇ�^� ��SC2�p�7b���{�k��L���E�kH��9����R�~�w�^�v��]`,��9��=�Pȋ]ұqxLE�Ms"�Q�.{��{��։A|,pR��{c!-���l ֦r=�N�`�aG߲M��\�c@�ڐ���+�ddN~z�_���fJw��k�9��=��6���b%���)���J\�_�Ѩ�^���[FXl[��D.���^Y;k���86�;���M��I����Ͱˮ�/���[�z�ZVeؤ9%dV���E�"դ�ָ��(Bg�;=C��,����U�n�F]%s�:���r��򁒊���ދbW|�1=���!��>��L�u?9J$Xq`l�Wg*�l���k����!��;�����n����9���@3 3���P���5�.�UE��ft�$A5�1v׸a�"G�lp� b#![n�Ӂ"�U�L܎A�㭓�!��	�q�P��l�#�{�i]�FK�LC�pcn����FK:8�+J�T�󣫻�'8���_�I��Bwd_/��/)�	$w�7�>���ܸ4^��#��ڰΡ���zB��6fM�P�Y ˳s$����MUim�lM�j?��������Z�����c��-�⼤U0";��ɕ�{dzz� UDv��f;K�����O���9��L���s��x?§'�G�� Љ�����:��{�n܉{ij�;7v�O���*/�=��ol�s*���=����Rh����^zN��d?�C��A����n�w��?�:�\F~�R��R��@:�kD���md���l��@�{Q�`�ֻ1� ڭ�aB=h��a��������\�=9`n	�rp[T���NM�[7N�J�!��5P�$|��b�a�¿@����
�7��L��"�u��,��KIF[���e*�uS�w�|�8k2&���	����F���}` ��"4��M�.�Sc&��q�-B��R��E�bLi�7�Z5�ޢp�8��DЧ��C���S�$���B�Hot�O���j>������/[�f��H̽iP�4���Bl~-2�K}�7�0u��h���k��{�l�x�Ff����^�$�dS���&ʤ}yt(#g������؈����'������]���v,��Ւ׺���AL�������t��*^��$H|����9�qU���E���H���sE$�tY-���A�IN�c� �Slf�B��esz�x�!���xo)��kS�r��#��L�n����co����';Q� ��؈�^�'Ck&+v+��e��:�l��_���}\ZҺ3vW���c!$Xו�GFhC�Qt����B��������Ͷ��k��TTOBA�,䜘1Ҽ��q&�2~�q��ټ��-��QM ��J���t�������Q�
	�hx��Z���B��X�7���$,�Lм� f�j:	����4��eM�T� \EoIa����O6N��T͑�I�P>$;a߰��7�t+�B	:T�r��ڊ������ d�&�x
�Q��Î��2}~���1���qG�?V�(	 C=Iô��
�&�VO�n��<[����u����k�5�jXO!yf���[���!6$��l�j��n@������(iײѸ|\��K�W�/h�!Q�}�z��D�'`A�?=}o��ָ�}7{I(k�ul�[����ܯ���g��Uv�W��b����i2���b���"��Ɇ�CI���@⸭Uc�_�ه埨R��/� �b�� A4Mqa���Y)�<�������������/�Ʉ:po��hw�5J0�9����d��F)'��p��p���2���6J�[��{�V���hj��c]��1C�H�����w�Bk]
3?��Gi�1ٚ6�>�-73�&4��	*徉�_�@H��e�W��1���j�Rr����ZKϽB~(	�O���1I[8��\w(����aJ�-7�h;��L��P��8��ٙ�<��'��u��'�&��O㻡��Be���>�;jOO�7����q>�!	2�*,����m�pZ��Y2�
�7���]#�9omY�-����;���7?f����X�g\q�n���,�wM��r����mAMț-A1��vZ�/�����6�-�S�cނ�,Fn���8��Cg):4� �42� U�/����Crf��=���}��1�-����1.������>Ird���&�nt�%]*+\�;����B���΋�+�!W:�v9C���.�UK	�m?��Ղ��4�ol�1��{�b{voߎD��Y�|Yy~���m���_nu�����v�؆[����o�'q[z0��x�,���Rj��%�aMj��9�AN���������} ^�~6e�����=���>k�N���HR�@��L0Y��0��`�(hE�m��I�|=4����{E]!}������bj�VQGK�1�	�2�	����2K��7����l_*ٞ+����lK8�o���;m��Y�g#`���IU���n+Z�vX�{����<���я?�ι;�w�o$u�h�6���F�R�.��@��I��s5��	�!���"a�Hͩ�1	r6v��I����>Hp�������>|�5��ć�F�ȍ�Ѯ��Ĺ���+�aO�/�5��ե���Iܞk�V*����KAџɏ�x��V��zc! ���ے�Q��#)�ӯP�5�'�����F����U�x��R�,%�����{,���Ks&
�%��;����6r�N��C����&ŘTղ����UV'n�XKCy={`��@�~ȗx8-"N�ѡ0�諾ZJ��(��������=�D�K���-'�m��.6�ߍP�_����m9n��`}���O���U�Y�&8#��l^�{�	��;�>��+�D��H1U��+%!�QP���o�g@J�=���x{���\E���M��;��т�@���p���]��
U;|2���FE�5��_P�\�ߖ�w��Ɲ��&��1�˂�)ļ��8�����w��[���ȾU��S�9�Mf>���x$g������G�MK6��b�y�\��H�Ư>�拓@9ԥBGsؾ�^#ea?p�]JF�����)j��W����!��F��f{�h�����	���o�����=��E�
 ^
�D'%vㄞ��{��H	/duFw�G��I�F��+5���Z�#H_����`���#_6��5�BX�Ș����yg��A�Jv�����L.�2Bo�.�����[L��0%Rw���_��$��Gj���Q`��Je�Bũ�="� Ե�c����O�D�"���#���gxfm_ᚾ�[�=��"���i����k���u��,E�8�xI�������2i�&��>��C�� *���y���o��`�
�O �0�̧̟��C�]�dT.B��#yT�2�#�v�|MKh{���˦n���ɵ+1�3��n���]9�����h��5O���<��F���rn��O �����6�;�@��&0�*u�^�q� ��7D��D��)��͆L0��5Y��VTL�9^�4�����t��#>�6��ir%��Vz>�������=4�0����1;�	]���c�d�%���f>-	������g�V�˨���t�˃�s.��%���f�B($�Da�� ;p|���{�L�<�<gB�ހ>����gJT.��ō�� b���`&�Bz�:A�tG���{�]��M�ֿs�YW6 �\��_Cf]��u�x	����2��)Ƒ���_(����J8�1	��w���Nn�z��_ǊZU�e`0z��&����Jq��i;���Y��F[U<�<���H&�L���Rǜ�2�x5]U�o�ܧ�#�� x�DХ�Et�V�BN����k�B���<�4Gg�Z�k��X�y�\^"l.���V�ٱ�@Lt���Q��7�g��YŸH�6_ܺ/���+��=sf���7�I3��wS���f�T�,�=�`����-��t�Sw��:��oG:�Y�q�2�bV�c���9��3J�(��1�Ef��:�"'l=�s���QC��zO_^�%��L�0r{�9�����^y���i>v�y�� �ۃ�6��蚽��S��ݿԵo(n���^c��l� jW\��H�L4���6��S�y���z:�_/h�BvP��)eeN� Ï�����3x��Fn|^�8�3�6ݿ�j.g�Ee���œ��;Vc����=�U��=tǐ�)_�ʧ��r}R�{������#�_O6�o7*x8A粯�"}ٌ+�2k~x����W��7��g�!��8Ұ���14�/}�=�\A�k7z`���}��	 �H�	����ˀ�.��[�A=0��J̱<�
c�Jv�H|6�﹝�=���&�ſ��{����*�Kd��_h@�$��wVМ14��/�
?����:_A��mXb(�Z��<<����*�m��2�3�<A���㪴�e�a�+��(:x�'�!��tt���^>�:[T��4�5���8��
w�j�o�i��w����G1Y�~�`�U����"V8�؍!D���=_%ש����Τe?�%��~*��(�����R��z�����ŏ3h�^�~)�;��_���,����0d{�b�1 �������y�X�	
�����0U7O9�
�o\��_'�;�}ϧ��npQto���Z�8SC�c��ͥ��mYY��y6`󂍹C�L��}zȂ!�,�S�\B�Q�?����ȷeq�E��4��C�;��1M���O9+��d��)�i{\n�j|ޔ�藦_�c+��!D�ٜ^��[�҉�N4���υ8�#$����� ;l93���נcKϘ+¡����i����T�����{ A�|�-'n$gF�GY�"�Ә<	eYM��/�g�Dx��b`ё�9zi�h�٫��T�%\�Rx��l���S��l\U*�� �!��o T�ŜK?�?��ݗ�)�ZZ%_4)��8��޴s�c�g�oӝڊeE����-����H�D7ؘ2��0���Y+�������͉I�렍�w��݀�!�	� �g��h!��_��op�Ů�J��d��2���ֲnpa�B�EQC� =�R�|tϱ����
��?�B,du$mY�'�nK�Pa`YE�#���E�W����[G�Z@#�w�S�k�	hZ�~B3n��߶e6h�}[R����& BVv4�yf!�i�V��7ώhYv���"'���W��N�n$���J·�Mw-�es�O����a���r�I �ӎl�	�4`����mmr� ũ����W�J��x��qx�8�7c��x�S��ik�ؗ���+(�o?΀p�`8;L5���#���"���nGxbe?��L��D���8�a�����Ƴ���+u��-����|�5����,��w4��r��9���dT�!s�O<�F�vQ���O�w����3E;��[���;���܋�+5�FGh��8UI,tָ�7iB6w��c5Q:�f[$��Qb��q�lCw��lV�v7�^��p�7T%����e��gk:K����B��C})a�ze%�1� .�åz<�$��[��e�$+S����P��W�'�W-�{�j6���ߣ����K�*��淣0�s/��ů�Z��D���fd�"��Uu���~ܻ�I����U3@2z���@��r�v8G6J�TDI������s�ݮ��Y��o�E�Ȥ�U2b6�KQN\��?�`��E`.�׏��j���1	��_zy���� ���g3d��G�Y���W�w�fY��#�>==��ϥ����O�;�ťKd���y
����è�jW{����m���]}�3������C[�:��Tf:%���Zrh_G��ߨ+����ߞő
�2G�>����P�~е��[n���VpA����n�=7�C�x���:��9u*���!�k��F{g��T	A[�[��4���Z��R�?��k���i6�;Ȫ�غ�ȑ�_z�1�^pB�r��]�Z����U�C��躪��`vV��rܳ-RE��X�S��nu"�WqKZ�p�q��ݩ���?�sl�=�ԃ�D�Z4D�*Xy���J�T^�0����]�\�����\�Kqݩ
�8oO3>bk�hO75^8(�:֔�[Y@Q��j4����+HT*�N�}��(~�,r��.����b��˴��� v�{;�(h�0B4�d��O��j�c��Ȭ?��璸�e4�:ɏ��$ 3q����7�0��?�*I�Z;1q�c: �.򒘎�#��M��׬w�wӟ�CE��x%,X����5��~�¥�w6Ԁ_��h�RR6��*δoV��������',�`�\/������b��>'�&#(b>�?��u�P�����I/}B����L�H�~�;w��#�7��"���4�8j�.��c ����-&A���w�bR��j����i��O�&�7��.|O������*�0/����z��rcC���S��m~�4�(�\/z_�K�*馃�v_�k���əŴ$`SJ.��U�����>�\q�9�fY�s�1�[V5Ӊv��#4!Bҏ���r��22�q�O�!�j�����^'��/��1�k*�:CFO��aw��PI�@7��1������#l<�Dl+0���	ͼp<�Y��hJ���Ipi���}��y4�[#�(OT�J_1_l���#z��"�[ �r��~j�ƵW6���
"hw���{lrep�<T&o���oez��J���b��OanR�c���Ro�o�G� 2q��X�G�9b�Q`T�>��#Cz���[3����F�\��:jt<��t��E��k���<��,#�A�|�8��eaa;��{�n�/ "����G�]V�����<���UV:z #����+8�H����t!T
E8R�]jD��JF$��o�̅2s����v_�p���`�)���25E��������Q�v��&��8Aǧ �U�p�J�r�.��˾���Jd=�Kf����G�u���;�4��� ����*w�Ilz&543��ra�1;q ��}�H%��1�*��%��(�A�=���y��n�w���Q���Sd�t��c��&F*�b=��\.X��2��^N��{����;6j%��d�=F�=�-O�.��������������.g���0[`ڭ�;��U��T���.+�U��2栠���M��e�J��5�8�Pkq�5\ڂ؈�}qiOE<]KdD�%w��{�s��QN���{��tJ�qAλ���%y3�l���Jib[�o���l�߽��zPBHX�o�&;K4��B��]D��Vp����tr��[�n�2��f>	��=���?�Fp�K�7��o�s�Zz'�C��;x	�|V�A舢4�h�o�-��O���C8#ゃ
�Պ�K"�k���b���f���x��"�4D$٥&�n��Q���~������!I�D��`��S�Є��$�Mh3��Q���=K���y�'�X�%/C�a�jﲨ�l}��� �@���B/��>X�̽��L�]bz\ݕ�Ưw4fM��ԧ!E���fD�Ix�\'���q1X��z��l�	&��!��P�}�٦ؿ���D"�Gn�d4�J$*1�9�Yd4(��"��VQ�߀$�rJ����lf�/7O�鏡�U��#ևK0u�Q���N��U��g�LЉ��8��R������[�o��=�~��<�b�t�Z�S	jl̏����+ST�m)�ѨAO�܏��$��*:�h���8�p&k���ځ�\�.�Zp��e3]o�:jv�4�) ��V�A�jΐY� V��N������k��2�w+Fp~�p`��
�@����{��R�+�1��m���sf<�y�JH�/:��L�jGD��2�ע�\�[��Fuf3��K�h�Ԕ�<�^@�`�=�鲶]=Q�<S���3,/{D����Kv�i�G	ibŐΉ`�Y��U9��N�7� 5T��Z�ͥ��s��\�	�J+0z9�������P�'��c���9 f>���|���z�����iLJe��N�c���[(d�[R�U\��\��ğ��B]����e*��>ʩ�'SH�q޻�0��'��~U�&�������(����YY���&�Ee�Wı�!�z�ԣ�f�!��9�����-O���!��R�~x�\�x@��<�;��JQ�9 +�l+f��d-z:�QJ�S�/����3@�M��Uٸ8e�E�H��X�!�GhIHP�fiU�LO������⃟�a"� <��8%��j.1OΎ��Hn�ϯ���b=?Y��Q.r�h�ס���������&�+-bC��&s�XO/�}���YjRe	�̧��I�_S3��o��X6�j�bM�^�X�(`d���w�}�ԹZ�`�{�E L���YF�=��Yu �e8���.�b��t��ip�r��O�}���1$�>�ڶy�4�;��xbH�;wE��d��HA.��e����'���	��r���/r��Ջ��=�l|y���)0�6?�e�dN�*�����dM1��zQ]��}�-���T�do�"POn��Ƿ�FÌc��x�>���=6B�,��iR�'���}[����h�e8,:)B�$+?��8��X�3�[�����0�e��TP�`?�V�j-�kv�[�����훻�Sù8v�U'*Gp�r��ml����=�{�x�J�ɣ ��s�����H�����S�MjJ	τF�m��p��0�z��ʐ$�4����ˢ����/�UlZ�{�{���Z�ƿ-��fd:"���n<15\��!ka��5�
j�v�ҁ'��K�R���Ѭ���t9i�U���楙
��ܶo�3�k���r���;��7wai_\MU~|�ߓ��1�_���	m]v3$�HBcL	;�w�Y��i��Iy�E�H6����zم1���#g#!�Z.�'�p*5���J���oN����y��&Kj.�TƆ>��~ǉ��ڗŃ;K�:�8���cҀ���oZ"q�O�gX�kx��pc���_���Ѣ�䥀���ɛ�"�]�%`w���P�W��#��b���mwlfx�q�Y9�����{���Ƨ�k��K��)ױZ�.AՌ�޴e���@A��2��%�l�t��*.j� Hq9ֵ^�쫷}�pA����䜗.�]�o�M��c�EG���QAce��x鶸��k��N��Wg�y�)�>�b:��]�3[hg	R�bނE��..̜�f5b$­��^~�"{1�b/�h#�]�͜+�pO���lCHFx	�wۘ�$E�-����W��03���~��^�&��5>�i�1{�J��B �j� ͝H �mC���K���ȷ�.i=�1N	�$l�z���TT���?�p8�\!&�A9a6���m�}0��Lk���2|9h���lj2g��俿X�k'A�-h�i?���(�/jIRy��\�;�hB��8�*&����i�G�t�1��+�y�Lr`>���O\��̄9)���Wh���|(��O�q����i�e���8����\�WAw���l����{~al�y�F�%p��V��+����G��P��,7J�M�����m��gD����g:�����JѮ�-�p���[����R�o�UOgY�"R�����wA�c�'��:�%*	�ĺB�1����l��Ix/_�Fb�t�8؇:9}���#���d��;Ys�b�
����	���n��p0�8w��-u{���P�F
����D�������?����-&N��5�
�=v���Qm�Ū������g�o ��������0��:)�q�O}������sJ���T���,��02TЪls��j{���e9<C1���6۸���\Bk��7��透l:�5�����A_��H�VQf8���r��w�``@��ݠ����u��,c ���-Gڦ�P$��M�88����o)U��3�	I=#^������X��AwJۙQr��d�k=�!T�G�h"n�<�3��`9 _<\�.�
D\
��b�.C���g��y$�Es��'�#Df���?8�d	n��e6D�����l�XP�h�M�q�B�Ij�ĳ���0�Ȗ�tG���M�Ѥ;UA�8}Q��e���+��[Ы��Ѭ8T���p���<��D�Fˌ�%s���1D�Ѝ���L �淬CZ,B�o�`�_��{*�}KڜP�2�̗Zj19��<�Ʉ���P�����0�.��ꛖR���L�"�ȇ�s"��ѐjIR/s��[vT���Ȳ%{�"�K��2d1 ������b�l2p���X`ؔl����`���.�4q��f�Si�ޱ�q蜹�s�h/fZh̯���	]��ܥĠ���&ֽ���6�D���,�#���c��⾉'�HQ�����pz���mX[�	�;�偍���������key\�v2�E�y��@�����a�q� ܛ6��Bȍ�"р^��ɫqj,�8�1��@.Հ��e=�[�O���+��J�"�Q�o[1bS����X�'�֞:Y�7����.΄�C�;���2��Y��EZ�G���{���Uxb'�*`�_�V������_�������� ��Vd��)2a՛�rX'q+��Ly��{C�H�8۲�nZ��~�t�r�J�i��L�������q�I�g���
�\��/�q;1�*Op������>���Xl�/͠ފ�NNM�� cn�����D������P1���~�)ӆ�h��w�%�.2
�s�)����B�\����Ea9���G��>�p�i%�e2���2�����H'!K7���zO�#��B��qPDG�������!̙������/��*J޸�k�4�ǄK�b��9W����j�������r�O��*keЬ�_��_
vD�i�3��)���R|���M��pꑼ^J��t��\����{1g�s,�<w��lcC�S!_q����g�.J6��G�tva��sc�ٲ�-��eKL�S�\�7v��P�A������ɍ�U�8)l
B2}l���-7�D�l��&�n��;,A�����?��𞒒b4����\�`�w��D�@8� GZ�^JP�nNV��uBma�U�R4ˈm�&��UzA8�j� �?DZ,c�^W3
��fW��S�I=Za·C�"�>�#��U��K�r�ܨ����E�)�����Q�4������-��i�QBl��W��4
���QΛ˗�A$�ùM�#�p[������	�#���{�(�n�e\�T}����$�'Uȱ.ˋ�MΕ���i��&*�k����b��B�!z��#�Y����^��۬��dȕjU&�P��F�x��?9�Vb>J��SJv�n�\�R�cp�0P-��&n�>�C�by5!%(�X�7�\�sH�=�	�YsV[6�.�$�Co�6>:x�W���1H���ϐ�j_E�Oz�,F/���[_!/e���)� ,A#���ZB�1N�s�$ޓa�Vh�����/�����&������F�:8��_A4�%"���*^� �o`��U��"u*?�c�g�ͽY_�lH9��O��y0O����q]ϚU��Ci��͟:����.���,��8 k�x���(	�\j� �m�$>u䁳�bf 8M�q��ùu�>$p(F�����Fu�"��01����Z�2������GD��d���(��`�2���a#�1�Q��d59D�yU�џ����l������ Ÿ�����
�e ���'��u6Y�Ъ�8�H��� =�F`�ob��W��jũ�"n�D>:Ͳ��iwK$�z
P�Kv�J��q�% �:����pW$��eIŲ�W*Bq�2^��k������=0Lb[�h�j����4{k�|*�ZWC)�Rg@�~wcw���i�����xPM������U�2e,븓qlV�)8VC�FT�T]rMQ�	�B�$Θ8pS�.E���|����<�HS���8f��.�̔�˖\0�gTAX���)}5Ȓ�J?-G@�E>�/?t�L�k��[��.�Gj+Ą&vkğ��V�y�9b����?K��������(צ�B�i0ʾG�C��Έ��RƛX2� ŕ���ha���%���xh�����;��*�Y�@$R����_eWF|����]��*U����I0c�2��ag����X@_n\��'���x�3�8=C��	m���nEGlT����r�do`r���}'M�N��	wdH�V����"o���IK��$�U�D����FD���
W�n.Nn��������ط�j.s;���V�K(gi%��i|��F�J�F@�Ǆ�4�xM0[^����1�$�("I��S��nuV�����w��;�:��3�=�ؙ�/��T:�%��d���!�.:�s��,��JC�Z�%M���R���T�o'X�����H�F�pWrY*Q�݂M�o`�؏j�mY�=x���3��~_o&=5	�_�<�f
ϋ=�(��ѢK]g�h��e�_4t��C�Ҡ5��#⢲�a�+k6�
�ZO;��þ��>���E�k��`9@���7]�!b�����o��A�Nc�@Y��g��ӿ�/��h��8u��NAn0����H'���J��06� ���4 y}2�F��VF	���1����-*��_���3�U3��xI�.|�,�y����L&e�Va[�
��h����Fo&�r0�$���}�3=�Qx�1�jX�q�B��Ll'�;��� �� F�Tū��W ��c��یN��ϒG���8�	�:�
�`��k���u\|�����U�$xtJn�梩�J=�Q��EL�->I:_�-�N2G�c���gQ���4���+S�D��5��CJ�s�L����8��䶍$���Zh�N���N�O�`ef���"f��#�x�0P⦌�6*�� �H�9�'�9��B�>���&.�F��!ڹ��2(0+�F��CS�6�l�8��ԃ���Wi���N��ns5?_E��{O{� �M�bW�ܬn�-�t�)��pj�h�*�����Lj���r�9�K�kLL�}�G�:��.�9nYg,\�qT|�ݓ�cݝ�~�~77̭�"�yr�;��Ҥi"���y�!�m-=���@�V�V��s
Li�H 1���V�H�auxx�Y288%K��X%a]l�ڡْ0VB�����[5��rJ������c�Mq(���md�j��0�gZ�Q豂�S�/�.���4�x���Y��y���K�;�V�<?]��vH܁|r�/((�T���X]�5��.��~b�������` ��ZSn�B
N���b���2z�'B��=��*����r�'JPa,���0@z�T�'Q�̴)���tt��������9Ɨ�!���^������8/ ��r��9�s����e#&@�ۅ��� kh�Tm��v;�{�f��s'��ʠj;�H'��/MRV��+���J�!����-[�̑�x���i�dz�\�R���$�*!0�֟6.��ӓ����1�,$]/���֋&�D�Fkл����j�:��F���q9B��2U����o���3�Te�i��>��i�7Wڹ��jY%Ņ��׺��@z���[�or��c;��Q�R
x�Y��7~��2������ޱ�ۑ~�T<��Y�,�廮���=�u�`hX��#�嗅��?^0yR�dif���1�bLN�T�Y�:���Nw�BKVq�M
r0[��-Չ�_����},e�[��R���Y$�������2���4]�V�x�3�������6]�Q�xE�5�[��<ʼ�����iK[�ef��YD�f-}3ħߤ��h��Qc�Ꮀ/��b�C���K�SX�]�4�R!u���h����sи3�H�z�'H@�.��D�Jm}ɉ�ۻ ���/W�܊|<,)��?h����T��[��z�'7f�����G�{��	�������d�dzh��[��$�y�$ej�'}d.r���`]�������������¬;��+�a�L����g�.�AW�g4��=��m�E;޶��x0�4SK���BhT^�s�?��(����H�+4q컑�, K��1�r��ߎ���T��F�-���1C��D�[&h��BM16 ��-��p��nr�����G'$,R���jSw���té�&!�/�S���%f�Yu�b����gn���2:}�u��t�P&0tCBx1�[��hN�v���-F*t���J�!�m�K�j�x��z����V�u��EX��9lU�c��}�������wDo��*.麉�
~w��u"����~_�	��x�c��{�� ����ba�Р�=��i��4�ˀ��8�GS�,�(ʹ3P&e�ʮ*&k���ZX�x�	��ٟߑ�h�9F0A~C�����Mʶ�P�"l'~#y���L�u"���p�ּ�moK�
�;!55���I��'P��3A���WF;��Sx�f���H����(7Y%u�T���֟v���8t�١��"@�ѝ-@�PgVtԄ�&ʔ�zb)�	W�1���0͞`�A����w��'z��	)8Fyw90��'6�6?����cf{�$o$��:�u����z�@}ީ��چ�����9'���~؉>�#�������8��I��/൩p����x��Ŧ�!؂=��JJ�I�ws�^����l\�Ϟ`�-}�g[��/i���W{u��?<g��4�T�ϋ��� ��4K&}!��Øt���W����W}~���]���o=���❛wl���~*u���Qd�e�(
7D�]�f�T�C����d�����A���k ����Y�dHi\6�^T��02�6�s9^�_@F�4��܅h76�fט�\L��n^����
>!n��Z����>2�7��X�+'￣t�7�,���Σf�4֜"�zW�:�,�@,����?�>�?e�<��ͻ�1��LM�*�|�$�&zM��H�"{��F$\J�1kK�z�
|HZ�����:1�w��I���{|l��o�����v�,���N����m�L[R$�i��Y�<#�5�$Bʑ�isEN%��GѶ�d\�h`����b槇�q&3�ii�2U��I�.�8�)j������iHD�� �t���J.��7�G,�[f�x�	~��Qת��s�Sͳ�E&�N��C�F����x�H2%T)1��萹���z5]����P�=�a���.Y��6]�.���ӹ%�Z�*��9��q׽d�'�7Z�s�"��Ffv���%��լ 8�� �X�$�ͯ����Y�������^T�v��/Q��1�'���8
}&�Xb��z9s{� �����
���AG��MB̈́��ml�z2GI�`�r$��98<���N�L�<�wu����W�d(�+��2��(�H�c��x����i��e���"Ҽ���n�2~�l2���YM���;%�#���8Y�x�s~��#9�
��S�jY��ݖ� l�{2�0��3��w�hމ׏�	��	��^F[��9`��˅��D�����Fc��l�J��$��=�]@0�q/t�af�^�)(4�V�� �O���8�����j1ߋ��(ro��?s�T�;x�j$��
\32���P�XG�E��M��Gqol��y�l�c�MBrF[�w����P%3�tO��1X(RGm��#��B^I��Ƭ~���^Er����3��"���Q�������y�[Q�o#��[�V�`x��0p�j�Tto�\d�N�k�����ά{�Ţge��":J�z��6S�~Y�%��U�Gh�(�����e軹=Zwi����
b�yj��|�0�+/�,Q�F+��bv�w�	�(k�nc�-���Hf�:!a�j���Wz1Sg=S�=G	!�p�ӆ��|K��Z�o (�bp��Vu�6���0����7X� 
�)�P�K{�GRd��6Z(��v��A��a��jd��D__�ͻ�9�-'��ƌ;s��9F{��$�I�����K
V��1�v���Ԉx���(;?�A��rqO������Q9��H� t�����	�����׎�(Q��2��g$�'�i���0n�l�zã�f�� ��dLף���� <UiUq+�����4B� Oh�a�X$뗘0iK�za�,�w���c�5K��P1p<�BXa����q8M�1II�x��/�[�M���ZYO�U�H��{���zfvM��b���wU͘Є��9nZŖ��#fAs4�D%��̷��4(�ʍ�d��u���������{lQ���6�ˆ�'��Ψ��u"���(6�%ٔ;R"��Q�C|0{񏴤+50���<��]&h�gV-�c=��s{2��O�io%.�hhh^�0x�t��GV�����,�7�ܗ㐋 �L�YH��Iɺ�ԁ (v�Z��jQ0F�E&�;5Z�(�`�!�i͠s���^�3���~|��@胸0�ѩ�!=z�i��Z�pb�|'�Ǡ�B@��V:7����"n��ϝ�X=������W&��3�`M��ŨTr��z��g���\|�^E�U���~ޚ�Ɖt�blB��D"�K�Y#��\P�P����p�_�K-oIԿ�|�%t�� �����vvթ�v���/�e�O����-�ѧ�<�?6˟J�GV��e�!�L7�S��X�(%�V�"K�UJ�ϱӥYx@w�B��~�V��������� ،*x�Q��.ÿu�B��S9�b���
Sg�#qf�BB��wY��T3a�7M���T��J�}��:h
I
q�,z�;�a�ʛ�1�O6����G��!j�\��(�[0���h�;$�4HK��>����e���1'vv#�1�Ӹ�T�^���pF�}�y��v�(2U꟟]c�}I?1�o�p�7)��8�U1<��49a�|[K�uNgS<��+n~ֵ����_���Ʋ�\��R�koLB��le�4ě�-&KV��&|���[�@���p��\�����;�%�rHY�f��mC�A���zAP2H�u X>����4�����J���g7�:��BP�c�-�<d�sA����o-E����V��Da��ͻWе$�v�R12(&װ��hH��Ay`���t.r�	���W��FjJ,�	R;��1��������&3M/R"Y0qKח����l|ط���r�M
ݬ8����
?�a�|3ԏX�o�b���g?B�@$���o`���v���	�xNx}�z�l�ua��|�r����D垺rìa��N��5ق����B�(�J������00�XlU�C$�6o��j�lp��z����o<�1��@sP�D#�>{+�fjf����_�	< �M=�=��]���+?�*5�i��s��R�c�]�xQ)�^��u�@֥'��0wcK ���S�7.�8�Dv+�|[1����=ϸZ!�R\�&����d{יc�����V�Mol1��q��)�Ā��YH�f��ӐE��G��D��R/@{Q�3t�~�C�f�>_!�vT&�"*KB���_��Ӳ\�&� |�3�ʏ#�=Em/�c�g�0:W�����d�����[�>�NQ����Q6�y�Q��\�']�J)H��!o��/u���'8���7������Ǭ�-�w ůJQ��R!S[��z�e/�d)O}�a�'Ӈ��hm��������+z,r���&�p�پ�k�R�%|%�isBWk�R��Bf)��C���	�V��7��Łp��a�Q��HO�P�������n�\@rFk���fr�*��z@s<M�_M��0�����Ӻ�� �	�Gp�^#�rOER�r�^
��;��E����^�	~<>����Q>�X�.�z� l?�4i�܅f͒!�U:L��� Q�+��$�2��!Ts��ㄭ�_!X�8����!�l}`ؼ���l�~�} [_k�c?S�r?H��}��p�Ʈ0��x��Q����vb�7����χh������l}6���{��(	�W̖ҏ�D�6��|�[�y��dީD;L'O�M8H(.G�K<A�F��8�C��h�Wm�ZC��&0��а��X��;^���y��ո=����~{y+��4������ʹ�k��Wa ��#,�<_�$x��x�=`���=�s�3���1�{�Y��#��ό��#��H��F?s�i>���z���W�H���p�-�C�{t��eű\���GZv���f��L���}�H2�RC�z�6	lә��s�C�λйf��9I&�E�ҕ�,n�pS���o$���J���v���'�����*��w�d��2�+��DA�SgI�C������K�|��)�����3�$��HC}_����ED�����ňU����"�N�?�#؇R������w�0Do�����^���'7�w�LA7p�;����ܚ�G�� 
{�gI����1ak�������S��cj�x3'LѬ?�~qo'��6��#!d�#�:�	����(D_;8�R8%�0��W%����DT^�î�N}�t���l�z+��q��9$��]܆�e�Q�#�4�:P��!�8`P��r�</�w"A	���PC&v�]]����4%w �R(�Y?��A�݇k�n4�!+ ��M��d� �5R�?��.��.�_"F��)��x�<1(���XĬ�2AS���#V!cZ > 	��g'"Y��  b�7�qF<.�C �'���z�-"����6�������\�N���]�a@.䠈�Wf��E���!! ��Ѝk~��yD�h��˱�H^ՠ��΄�m�_��&=T���`�۾��J*�*��.x�1)0�r��|gS<����%r�2K\��0:7��
�l�5�fn��;V�}���&����.�[6J��>�)W��=��mt������blxS��&���b���k�UqZ�8�
�?[��۬т�D�=���$�&�낕S;�h��AN4~0Ą�y�"�95r\��i;�Y�������gF}O� ֦wa�; !�-s>0]�)Dl�K3R�U�;)5�&���^� NTޤJ)=B�<I��۵.���o�ׯMlb�2��/���D�p���q��X�P�){ڧ���7��y���?&�.��5�M���g���Tc����\F%��Zv�9�h�=������N�cw�A�BJ�B���G���\OV���
4k� 1�O���$r�����1��H0�G��+�	p֏��_��g��9�~�q��6�)r��(�U(�>
���>tMl��A�K�N²�Qtڶ��ea����'�R�����'A�NO_��Ut��XQ������ɒw�h6ޟF��A�(��8�:-�����'>w��ĺ(�q��T�Π%W���G]����r��QX�` ��jo<,2��ib�Ԁ	*�ؙY�<ۮI��J��G�������m��
�\LKȤ3��߆mc���@mX���C�ǂ$�Hc������c�wc��[#m�.�9�����4�u����	�E`��<�3�`��P�:?� �:68@����4o�W!�'�zO����8�on��%2�%);dK�[T-�w���N�s|��}�[���[� �/s�K�:��ж�o/W?����s��~Ӻ���ooz��uR@/3OI���͡��ڵ��Ӑ��$4��0��b.�߅�_��EdT�m�u�ܸY���~0}�p�e!BTN�C�X�[�F��G0�%^��1�7;��C"���>��_�:��@Q��jIq��+�y�mH��.��v��E�,;����0�\pc}ƥ��[;8^��Ih��*��`6J�io��o���wi�6��0�Mм?!J����?E�/����qy���	W�k�z���$Z\��?�Jw�㩦aU�`�	D_�:�8�8^�+ �d->����=�)�okh�Z�4����D���Q[�~�1����1}�,���q�x����g�ܧ3�
�p������� hҶY�G����-t�qf �D�R5=9��ِ���[ �t@T%�a�?*ʰr,���[J̿�0\��s��[���M���Ը���K�\�|u4����pY䂌jX�J.UȒ=ߗ���u�f��@""�3M�3hˮ�O]|�����{�&c��Ϙ%?ٺh�5C�r�;��]e���� ?
�΀ub��h�&R��mO��a0�S�z3��ތ�\�c�� <�ҧ����Mc[h�?���e�X�M#!a�,�]���Ο�$�����C�m�c�H����d��$Ӥ�- <%��8�m�<o�q2'pj<��Q�dz�W��DR������ f&����X��d���
1�1�~�t�{���}s�
��C�:e0fA.U��2�
�%q�cɨ�곜��?��`�mT �ⲻ�*�&�d�f!rӼ�<�hK@�Sk
� ̣��N�lYx�hN�b=lf����e���`�����z�
���}����Nc����������*���j�t}5�j׼ذ漱G~D(�Z��0Ts�}b#4��Y(��ݾK
����|12�#{~�RG5<�(���&9�ʓ��D���.}-6!�,�Ze����
�{)�)r��ui�-���K�%�����-dҔY�1��8t�`��M}*�/�}�s<�����xx�N?���e�xg��9��+[f��G������N"r��=q�Z�����dAN=�]Q�.Gi��-�v��+y�v?򠧐ζ��M�`2Ic2��>b��uрeiX���Ͳ��`���b�Go%yQ|@�wF޽f� ���_S����B�d�7�)pk������(��s���ҏj�8�� �u��0����������{v,gb���鲙N/FjJPm�0�k>/�	�Ρ�xε���U��.㟩'G3�cc ����Q�W�X� @z��#��0�:�.E���)NZ��!�n�%��E2|c��g���84���Ƿ�
v��7��̖��$&\{əRrCw�[|ȵ7�G���Tvڭ�:c��1w%�&��IZ�)���&�ϴ�K�E����5#��&�5&Wd�4gp��^��y	�c�U�M� q�fnr�����;L����B�Pˡh��;�O�.��#��^��b����$�V���G<��׹�M8?���<H��\���.V,�nYh�=?�|^�����Ч<�[��O>n��#w��yl�V�5	t�ue@c��.��zE���Xr孅�_;�����P�0��h *�M@�����ⴥA���� �����C�/�Ϧz'�v�"F��u�{F�bf{e[f���֖�e7�(����W&�����N��u���������"��!��끈�MhC�>�:� &IX��:�d�|TU#��:���G��H�s��szƧg �Z��`
"��c�i��|s��#I��F�9�w����tDա~G�!Cs�ev(M��&�TKD���<��VT!�]��'�c��s
�@߸!ls/�{@bIxJ�S��`%��k��?0H�Iƕ�!�3mt��>��u�ȃW��W����c�m�7�p���ma����銼�+l`�"O��^p���+�{-E_^~rYj̚�C�֣D��ͻ��Q�u�]0�C&c4_f��;������4�n<�H�@�@5H��)],ĭV�V)�g雜���Q��,+���O����ǭ�nξ�E]S<.Qh�@�:?�p�P�Z<~ۧ�u,3�sI�2 �ZiB�k;�叆ہ��&�t�'�&���Iw��l�\�l��Y�C�/�)i��
c�v���t>�N\�b�SV ��҉�P��
��_
�b�,ػ=>������ޜ,��2�Gׁ�z�2Y��Q׸��S!��qr)�(�i:P�HF����g�\��*i8N�v)N᫘Ff��u4r����X�crtS9�`x�M���aQ��0Mf�hAS�$��������e����`��a���OEQ�}=@'{f���؍��lEY����>�_����ݝtT���������L���'u��iÇ�����<���
N'KE��)cI��U�#dݘLs@3�6 Rfy;'l���5J?<(
nl4	|Y<e�4���L�[��HZ¢$S� ��	�|c3�k)��#�U7�Vf1dp�G0�S���V�r�g���V��I m% �mܖ0N�,�r��wDBH��D1e�;(���)�������1����b!bb?�p�M��3�.�gs�ݎ�nR��A}�~WH��W���R�᜻�����z�Ci�+�^vs��Ђq2	�R1^1;�S೹�hY(@�0�|�.�!%��R�
3��'��D�r�Q)���_	Eu�T��O�d����QLTğQ�P�|ӽ%���+z�p����W�ޡ"m#���x��]�Ǌ�71����d�)��� ����d5aҼ)ڽ��n.�>���d��!zUj ��u�k���;J�S�GB�o2�Ռ�� M7H$I������	(j#SϺ���3����ou�$�����#Oo�ʰ~��N���psB�҈��ǃGȾ��1^V�R�w�q�κ������}⤰F=�g|+��]m�����B^��u���LutZ�.&F;��������u�%ݔ�_)W�Q�򽁒���K:�NK[^�l'��!;z2�!�0�"�	(|� ��ߏ��=���,����U�!Jڍz��W�oX�h���e�D��B0!�G岁�ß�}�,.�lZ����r�T��2u J��C_�4�|���K�����C_j������)x������>V��"$�,B[��M�',��H�����<¢����r�^��4ef�!P����}��J+t�i�u�"[�gn�ڱ�
wsS�v��s٪�2[�~���}ʈ"�PUf��O��j<b��V�۹�6�-�L�JF�qXt���7��\Ā�M�n��P�Y5�� aD�3��ߡT%qk�Wn(]3u:���i�'ٰz��z�{z�@��(�S�3�&6EE�_�˜����;��*lZ�,�I�N��$�珋��$��	����׌Ǳ�vF��������]R�xX�D��:���Uu�HS� !��q 
�o#����;0��\2B.�����1{���[����X|�M�ߦ�RU�%0H=����Б���)ѭ�.��w*�-�(��O����<��jz+_b�}.p�|-�X�'�M�q�SM��Pf �5M$��4.C�QG����B�Z��0c�8#� �j��Q�
�M�� }���KrNz�ey�.4�)p 8�įb1
^�����K�y1��S�;�je�Ŕ.�#S>��̼▣6.t3��Ń���DW�'���wj�K�<9��3k�W�t@|Y�E5��x9��}Ạ��4�� ���\X��ŕy�v��ߩxT�9{NU�:n����g�h����̓�s�c��ym%�]'5����8vc(v`fZ
O �"�rYp�I+�U�^PZ���A1Fsu9�X�H4�c�b��Y�ql0����?o9b"U��T���w�{Ur{�Q����-�0Ѻ����n�+�4U�]���0sȒ�#�v�Y@C�2^�h'��f���某�Lcx"1�W���ѹ@o'Z �Q�Z.��<���`DZ*#X B��F���W�+�$+�.�!\m���~~!!�Q�/`�Q5?�?�M�w�j�� ]ו�^�H�$Д�\ �C}�O̧5���2̤�>��6�a��5Y�(�
�����L��wI/��� ½���%z��j�9y�`�x�������?m�s>hfH�z��z�E)��[���kUk�g�I-8u�yü��) &+n3�:V����pL9�D շ�������Ia�&��d���F��P<�P�9�x����|�M"�p��m1�#�����v�\�v���1�A��b!�/��w$t`.ZWTb�k6��xB[U�j�:$���I��T$�DॽZ���~��0W�K��LC�ć�*���C��t�
2�S����A$�ij�E�;5�ђ�߉	A|�T���<�`[��D�VFС3+�LK���	�{�'��ty'Lk����%�Hqޫ j�#��[q�a�d��EU����zM5x�iso:����<wW���L�u?)�9�hb}� >�t��B�Mɭ^��j7-R����S�8_���������P}_6%��P�&��d�M�#�?����?�['�-�+�N��\,�2�����|�k�Ш0����;jo_���ܹ�5��	�{�F%Q�P8������������9A�,��^E^X�_�9���!$�.��
F8����R��m�:䃢PRS��*T��� }~Y������)����N���:�G>���Y�U;�]W���ɷ�z��{��%�g���iNR�1�������l���Q�aqjĲ3�R��_��ʳ+��`�4��H{��[lBYδQm��I��b{K��@�bSߴ)ƴ)I�[�8DE��Y�0��̇�b����\�[E?��USa�� 3I�	Ec;#t����tp��4��	�<K�2ӄ�5��#Rd�� 1��ǂ�7�\|&��:�/A ���3�?-,`Z ��H8�O	�2n�K��aӻ�S��O���`W:�����/�KOc���,;X�a�l��'S�a�&�v� ��oq��u�s�qvI36ۭ��s��j1"��h�-����s-���	ozX�y���])=���Ln9u����w�9���0|�fd�ހn��tIa2m<�u�=b%B�\wJ�JO9���g�h-��p0��!)����	?Z���&�����o�z�p� �L��"/�ћ N2���oȞf)�]i��c�Kw��I������<��d�i5g�e��r�6$��ģ�\����]JС�n�Ȣ�p�sa�x���0i�#R��>�g��e���	T�;�B�ZA{��m	w�����;i��cOX�8�$۝vb?��૮y'ug�7Z��k�����M2�HB�S��
A�9��u�����o��P�<U�3��}�v�L,y�'�=�ďu�	h�I��%a�CKHe+n����z�����vǨ��M{���ӅAL|Q�19�TMHp��_ �0��Z�!2�l�~9��ڨ�y�p"��ׁ�f��[��Q̙;�<���t�dn��8����L,�#��}o��}��f�no��M��FG�_��).��c��	J7"���M�x���U��)�Fp9��D��Z��@�};;���7k��M��UqJ��_>��r��><��6���E0��ֵ+��!)ү����G�?9,�߿���z.2�P���unz�d������%�Ӹ8��*ix2�Z���<�J��;/�b��_�Y�C?�^�hؕ9Tnl��3��T�f��!�v���(�L�\U�d3�ͪH7�n)@�ٔ,~#8@�M��C�����Y�C��S�h�ރT[�2g%����6C����zqOj3������O��M���ÀppY]Y�#��L��E�4�'AZ�F|x�3��ˣ��s��?&;KY���@��7,������x���Nϳ��O1u��Bv�<~�� 5�},re���_���iu���Nli�4��H�z��&f�˷�E�7���Z���m^K͝�8���{Jn�6�D�_8u�/� ���Z���MEW��M�>��5��˽��3<ގ{G��K./HkpKU����;���Qt[�fV����9��=f��1	�xO��{��H��gַ��rus~0�v�l:�N����"�Ol��Ί�܋���x���[Q��υ��*w���M}��C ����D!�ky�/�l
�W��?����څ�g�HM�(���El��b�T=&7Ş� J�%t�ő���B���޷�An�	 ���*-ҫ�!Bd�d2������'r�S��]ޭX��T��7�����,U
��[c_��p���u}���q�¨s�όpN�d7�	��wd>�n}=����I�+���U��U\����UV1 +YqAg�0.�ǩD�e�?12p���(
pa��U��\���1�-&2i�U���K7'<�p1�ϑ��դ��&��CPK\e{Ď�LY1�#㯍P0X =�%����ЗA�g��p#�n&�OE���b�ƼT��+pg�ZGi�/�:���]KW4Hѭ�gԠ=e�9��S���
��3�j>;��O�v�=[Ԡ
���Ч���=�O��h�7~����,�M�w�l!T�$�[�KQ�Yd��6м|��R�xj̋SKj�A��	j��D	K
f��;*W��bH�,H�����*w�H�7k�ob��qR�VsX Ȁ������7�"�~ƻh�a����ӵd�ſ��ƼK���޾��4W��/����Y��Ť����\(\	Ve()'1;�<k�TА�����؃���Jn���W��c�z	�E&̯��j��9�l�Ѫ6_Z���r�ϩ��6�353�7���=^�M<[YD��Y_lN4�l]�G���I��o�i8�l�4MG���A���FZhR9@�F��M�Z��i��(���֑5_�?��	G� Q����h=��d��z*a$�	��m���+k�^H������ Փ�z�f>��z%ǚ0�fvU:KRa^��)ar^S�Q�P5+���p�^�{���b\��m�����K������2%��������(�K.#KG3�����0(}�na���m�>�j�hy3��+��3ɱ�䮹�J�3�����k�n��A�uvAcI�P�|� (�҃����,'H���;)�gӇ�;� ƑL^��͔�h ���:���6���ܗǃ9��]W�X#�Z�
���%���`[���UIT���P����s�l�H�zR|X�T`Pm%�2u[����A����V�+O�50�Vۧ^N�KG0��/��VA�;<�ᨻ���R����1�>��N-ڀe&�)�(��jD!�*���=i�λ���.������ VA��7L҉/�.�<��_.B����ٝ �/�h�1� $��ߞ2U�ų��!$'`e�:�����a�Vܫ0-^��]X%�*�v!�<�MK�m��]pw��Ᏽ����t�w̅�et�E�V'����Mb�L��.���oUĦ9�I60îD�����E+Vj%L2���]���lt��Sڴ��Oa��4g�)��j�bM׺���m��t'9s�S�'Z~��L��W��A��쁮�p���(׼Is�����T(ߖ!�
�0���nsM=�o��[cD�Y�o@���f��E�k,Dm�9��^�`����X��C���P+�Q񪀴���T��l���K�-xAe�7A�o8S�X���-|2x~��9�}׹����$�s��I��}��?����v�\��ɞ3暥?�v�qe!?$D��q��ĉ
W���g7Q�g!�lγ�-�iX� ��P 	"܋�Q�A%vfݐ�=����D{�0s͹$�9�+�NhusZPD���ciW��&':�p�%�GyA1��$���P�ʤ��$c�	Q���=l!���(�(&1�����x�&2Ѕ?2�َ=-��|y7�H�`I�S�ϸ�K���pҫ;����
��W���ݦB�5E�oz��Q�W������Mޡ����B�P�A~G�,���Ѷɢi娬�Žz��U_)�n��q#K��$�;$\�bÁ��5(���������@�g� ?`��ZX�3���D㼪����\��ֶ�[��m	n���_mokN��
�"���"���j�!o!uI��#	��!���\��;Їc�Bݾ�2^5=�J�G`�:c����^U�^$$؍��|���Ģ$H}xm��)�A��M��'aٰ���D뗶���!Ph�+�>�M��~}���i��]�;WZ���l,����re�o]�F�$S���ޢ�n^k�~�x���"I_�莸���$�z%,;����Ǐ�+꺣"��)�x��3��9@ke�����1�4s#��3A��ڪ9-z�OO�L������7���=ئ��	��ԘWq5L������T��E�~`��������L��TܙW@<�*=�#����*�C�����Ȃ���W�]|�1;�wv��V�d~�f $��.�d�I6ڢD�������`Sz��7z�AN>��� �&F��D���5���Z|����\C�^�Fߥv�Z6K��Oo����oK�/��ft,���p4����{ L�
�%��J�1rjqE��w��8�~x�Oo:*�᎛��qr=ďc�Gu����j���\�j!@�G��#	����Nulz}�0��P�i�\��E���2Dr�.a� �t�� ��r��������%���fW} ����"��Tn<�Ɠ�"�92纂A\���@�!��:��SJz�'�)�+�e_us�<�ufAC��M݄������+]���!����PL^���䉆�[G���s�q&����e5���A����i@�e�7��z�=Ʀ\�Y����c���-1���^ҀG��|�(5�D,z8f�c̉�cs�.��b���\ϯ��\"ǣ{-�����C�� ���ו��X����)� o��Ӎk׻X��p�jÌ��&��1%���G&8η�&T�.��KJ�w;5\�u7tzaV�����!RX�P������b?�(j��T�P�R�S	�$6���r��9]N_ ��z+tۓ�;� GZ�H2viY���G� ,;�ʠ��b�,Q�	��n�������䧡�D%&�%5p��@'�z���%H�\������{K ��2�P>�幎U��f{ܺ�|�#�0�e���+��Ds[��<�j���/x�i)���H���8J�g�~�@odT�bT<��Ƣ���k�HK]#�$��f{G�/��I�p����p�q��#*�J{jm =�D��,�I��I���+����np�1;�o�f`A���"4���wJQ�Q�c�%��DGx�Y��F������z�8�R�9X 	��ʜ�tN�X3���Sp3"�O� �MgV�;�����2�����/�=��pxU�1�&� ���Чӂ�@}Pjt�? ��
���zǭ�f�haNJ�Ȟ)���+����F���p��>�!ܖ60凁<���fL�����������,-��� ���OˈRS����iyy�{��b���{�-ŝ�{�o��w�R`E�\)�˸#538At�3���܎V���@�z�I���a~yr��HShy�w��*dB��O�Nt7�6;<�M�-<K��͕�����Q���%ڞ�F�cW!��Il?���	���0{}�Ad��7+�+�mؤTnT.8f��3>��a>o�]� Eߩ����&��wi�Z���x����J�'� ��!a�6}G��MPY�_}O䳐�B_���
,ߏ�������_�|�H�}�Ζ��T �G����r=Y�W�:��0:ǁ��;]�w҈�bM)�]�P(e�����j���( �}��r=f*Lbk���_������
ќ8��_���i5k�)��☟<��[0���[H�"3�>�O�rO�^�5��u���A@�_4f��&FA����*��D٧�
��{��kS�(�j�����ib��/DL)��"ZZ@�?��cy	Ǫ�X.��1�@|��ܫ+�j8�$٩��b�z�U$�M\+���ͧi��/��{tN��4�Y���l���NFJ:������~�`w[G�MY�zٚ���ڶ��U�
�0I�Ӛ:ր�t�X���62�r;�3c8~>��=#�����RQr���x�|8v���X�rJ�!O r9���E�eS�����u��X���,��Q�b�H��^d��wZ�O��������ds�vZ ��w�]+����k�G�p���?��<�m>&̝/Acna�پs6 �o�����y��[Ƭ^�����]�V���@��$�y�n�٣�:�1�6Gв ���j���t�u�k9Y�"�H��Gg������4��f|�v+$ �=<��➧g9�ճ_�S�v�ߒȏj���~	)���R���X�d':5�b�����eoG.�!Ԉ�G���
[��[p��r~��*t?S��I��L.�}հ�C�+$�_OE�����������r���M����p2k��FȎ
�B3�
���h�=�}�b�}�)��J��bo��_�x �ec�R%���Ln�32�a�D�.�|+`ai��X�R��m�]��ߵL�m��G�KQ*M�:�·̜9�o��cK:J�&�3t>)����(`���\������%E%��;��������jaҐ���G���!���Y����ʌ�Q�q�E���N#R��%m���$)H���ݎa($O��;<��Ɏ�f�jq�h-�l�����ԩ�2^߷�u��Ǜ��ʏ�qW�c����1OB�R� �� �(s˰�n�/"^�i��m^��.͛�6�";:�3�I���w����.����:}Y=�=ٜ���2��ގ���Vh�;y��L1�bC�[�j�O��;r58�x�4�v�����	��6�o�';	J�?h��Ą�ĄA�i9G	HQ%:��� ��I�c ��ϰ�q}d����Ϩ���V���}X
��3&�ҸYZ&:(��������g�u=���I�?��(X@+�x�~�J�~Í<4�W��z6NO���Bit���>/ź�)zq��X�,���8}� �h*�4|��^?�����1J};l�,��<�����m���Uxw�JNEr%�����>��:!J k�9鋮��ݢ�����G�9�ЍF2��: |�UԤn?�މ_�̄OS�2��$���&U��K�'9�7���"��Ƽ�-q�����i�HG��qi5�=dB�Q��nR��d݀V����72%�q+�\�(�^���L��$�5L¹f��ثN�0��*�S��l�0�EX�_�X�#[�G���#�:T� �
B���v�8|,���K�F�z�nO�w	�~�5w��Q%F��,�7а[N��ӔMcx����h�p��X+e��,ݠh�f�B�nP�p]栔��h��-VT�A�IqA+?�P��+@I�=�0�P�t��)̦�Br�ńG�tC=D5x-��az��kΒ�Q)�{J��vu�cMG��&`He%�l/K�Ρ+J$�f�#Q�k�ܢ���8����s�m��˹gP*20��Լ��äB�ṾM!��E�1r���Q%M-��س�Q������ɄQ" gu4���;~, �Ӑ��_���H�C�r		e��V���s$�a��|��d��/�qU������ ��g����y�k�lz5L����Ǉ��hg�4<�/��C���G�&Ξ@��1����3��ߤ�z����쟇y_9Z��kZ>�[�N.)����_#�f���wQ��f�?�p�c$T�ě�\1L�^ss�GB�馺��!p�Zu�ېX���<���Y8!3!nE��6���	���,70Zh���9����4��;��H�<Ap컶��W�0���ؓ�E�����ԐB+j@׭�-	U����3IO�s�5+
�\��G���"�e����N~u2jF�qJxqE��ƀȧ�U"XS���9���0s��j�^�4� �A����M���Z��%��9�3o@�V�Gq���>K)�ʪkSe(�s��w�.�J�Gf�ɶ*gfI����3�t+_a.���1nMO0�	�XM��6~���Y�Ӵ����h�l�U�����Zuul�l��.�ƇO�B����:*���qR��R��$^�·>ǃ�J��C�|E$�k��E�Ku�߁��oh��c�h���j5�<4���y%�kc������E��y+�ޯ<�^�ܻ}�v���1ڱ��fȌ��p�����C)�8ͩ�ū����ŀ����fD~����s�S��,�J:���-ޡ�UK�X�S	�uݵ�"k�^t,��{RV?a�8_�V�U+�R��5q����-wݲ�iG��+���<"�t���'�*3�ۗ`"�}s�p�CZ�O�A��ٿ�Oղ)\����^3/�!<R�dv�P�1GXG�p���t��oLqU��5SZ'f��;�y�͏�Yۜ@O�{PY��^Ӎr��~���"���`���8%�֭gD�~�D�rY;p	=����'{���̕�}�+i��Ժ����6<M6h
Ԇ���
����Qt�>���1�L��������Y^b�2�/�������&���ՙ^���0.K#^��xU^>�Q"�'��ˍGUI��1-���6�f-����$�9C�Io��$HY��j3�N�˭��o5S;��0�V�l
 �O��Z���f�W��:q�\m��ɵ���E�k������?>�"5��;a`�ݝF��|�0�qo_���q�]�V��H��h�?zA?u3��c�}���adC,l�O��\��i�����
)8�_�����/�)��AA&���`�O|q���j,�֎3`l�GMe��֝�����jm����+�~ED�7(��db��QI����J�7�DGw�-N��_r�z�BH
�/�.�ң��V�
��,A&�[���pƱj�H.u�37˃������<(���W+�i�f���M&/*�1Z���7�9���^^j8�x�B��	r�����|���/NW<Cv����z�
!�
��D[�k�����塻gQ�N�V1�8������W�{s��<�����+ڀ�ޅ	I}Oh��9B���yawۜM�h�a�~y�s�Ԙ��"�� �,��{]+��x��Q(�-<i�Df�!0EX|E����k��nx����C�����ç�΋R&�d�0Y<ϰ6�p���?7�U��Nqr�%<�
�����]������e��NҠ�y͘J\ᡍ�:4��CF7���3$�l��yᄷ���J���A�=�K���q�p��<�������"1��-��5H�B.ǻnF��s��ҟ�~w�w+q��Q��ي��-F�iL<���7��o4�>4��6���:i�f�Ys�8������gI�]�-�oDb��)NUrXW"c��?��#b�jӯd���h��$a������e7�kS�#���#��9��t���4���G��0���p��4�ڻ�Y�k���}�w�_Vz�3KjH�*��@�c��G���+r�N]Y� 4��`#��-w�
�-{r�(�Mw䪵\z�J�qn�朣|?���~�L;������j��A>`�&�c�����Vi��5�6a���?��y�(0|9���M�%���Aؙ/�S���E	��/�"6�pR!���`0�ZTB�9P�;�׵�w�u��l��n2�-'j2"JǗ���(8�"�w�(����p����>}� t̝f*.q�%������Y�Z�I91��O���ߜ�C�%�y��=<��L;6�����
�o�RE��`�-����D��
���h�ٰ�pp����Z����2܅}k��p�-g��X&0dw/��B�|�즓ǱX,�-�D�B�-���D�d����\¯��-.�4t��������J�����MK�|�׶�K�+��-���L�+q�u-FX���{1�W=_�6�\v�sq`���J�9܇�_m�r���Z��z���ʛۇ��zž���N;��`U�Ң���fN��"� &l�#��(t�����Yn�_M�x��?fH�me���ܥv�ү9Uln'-vy��W��gR��Nj�Z��o�2g�k�st��=2at �uo�QN4(-k��c0�_�񤘡^�����Ɉ���M|O��n����D�EViv��o/jPϢs�z��|���H�� ;#�wt�N+�yn���&j��I#,d@�@�����V?>R��#0���WX#րH�叒���>��06 �r,N"�u�������#V�s�����c�ˌ4$|�%�s�x]0�e
bJ�A�֪� �����U7�	��5��q�u�����t��̐"�|">�#1^�0I�o8J�?2bl�CR���GW�ِx���k����G�	��O�D��������R+�
^'N��9&�}�G�:�]Xf��6�O�t��I;*=MV��F��Z��4�!?[x�%�����ά��1
�7�S�B&��{SQ��BH��T�ny�8��<�:U�����[8k�O���
[��(��I0��W�|16(��� M���H�2r_hY�[�C��$~��65�}�f����p����K�`H婠��U4@����2	;���v�f����A�9��}��޾틚m<�g�#�N�^;�VP1�%RGz�C��>YZ�g�y�������W�쉰��c�(k�T��3��Bx�A�"0��cd8��Per�3�+���Q��^-�xj�4<3˸S���2�}9������"-���pDwe�lۭ�����󝐋knЇM����)��q�d�V�*�E)����K��N�J�6��~��$��y��
$���(��c�;In�yp�"�[g�Y-�[� -��+�p������G��ךE�V�U%�/�n��	m�O�k�VY��u�k��d���n�p�U�@副rC.^O؊�$	�l�1�W^�J�J�:�~J��z��H�1���J;Ҧ�C��>�������Qꀤ-��2>6M�o�H�W�Ƚa5Q�����j�G�?�� <T4Kd����!`�����k6.���B&���4t^��̧H����4m4���#;�0;�"�)�e�g��9ŧ��Q��?)>��*���l�JD�� O��RY���r�I��E:b�$�"�?��1Xt[d�*�9a�l����mo�5,˔o��?�[oQ�~T$@��Z�S�
Wͅ�ת���x�&|*?7 l4+�j9�XBڑ�j8�jR��R�#*cm�^���(5�O��P�/��Af��K�u�HVO�z0n
t��Y���rN����4��:S��:�F�i�Ѐa�6�Us��.�I���Iх�!��=�''��T�����p��4�H�F�ҳt�I�ͥ��R%�����y��� `XmG]@����pw�x|��Y�۾^ �f�+�$U3�G��+f�?��X<9(����ތ�p%7$c�4t>в�`vb$y�`�%��W�|D�v�8xn���p[7�����3K@ff���x']*=0
��0��jf*6���J&c/{�=��#��R��G�=N��� b�L�3�ʂf���P���c ژ�tbv �p�/��g�e�,ښ��p�HZ ������7hC�H���ځ�{Y�!ђ���5�8��ɇ�t�hw���O��� +�۔����nY����44H�w���u�o�b�:V�(Ico�
/��GSӂkF���V����C��g��`Mz������g]��g�g[�3�n cק8�Ú�q��B*-],��$8�N���|wv�{I��^&� ��F߸��L�D��SM *�n�J;��_�O��UK�N�<^ŭw�Av�����q�i����A�n�V�P�4�8Zռ���:�l�>��O0
�+�����+�@�qg|�J�(�v��QjF(��ZO���@d�����
�__����*�����}Thh�-����||��O-���0C�T�u?5�3e�n����o"���݀���y�� � _�yn���ە�63��w��T�3�Oq�Nl w������Ejd=�c�3�A�P�NG3E7��{�����o2��Y5��:d
bX�jH��wP�����������gz�g����v�R���V(V*�ɑg�)���EL��i�IR�L�.���e�����x� �	.�O/.0p8�]q$��O�Z��׀:�<ە�o~%���` ���1��|��BMُ���޺/W-�&S����h�m��̨�Ό����+.zZC@�P��&m�Y��p��V���JYp[c�u��E�j�\V��E,e�ˣ�i�87�KH�9w�tPe�|�����h�|���׃�Ә��0v��#¤�w����]��Rlrep�@��I��g�o��Aڇ�'&�
��xg�*.�&oM�	����O�|'���V�7��q+���5`�굄�My�r*��uV�;�[�g����]�� m
~O}>��:�2���C}9$Z��(�y��s�DsC�?�k�����ё�S+�BE���pڳ�誢H��>O���ዪ=� �_8�(}���-�Lvm�'$Ϳ��`�o�>蘏(f)��rA6<�4"��FZ*h(��8Sw���#�;j �\��ӝ��c�m�V��������+� ���Y���J@:���$o����-a�H��GN[}�8p+�\�GΣ �br�s�p�H~��-	����J�Ȁ�ɑ`��~� c`�D����j�]�A��3�osNL��>}�W����Ov�r���,�p�$��~�Q{ϼVτb� n�8�>⮿��-Pe��G86�I�w����&�4�գX�M��i�=�"�c�%����Zg83����Иy�W�,��yg3�����*�E��am�]��[{�>T�� �C'2���\�~u��x�(����/����팄�'T3���������b���8⑫Pt�Zq9D����p����P��nf��oOe�@�]2��t��ۦ0}iv4�|M�P�1�G�gx�'&M|p	9����(,���>~23������m>�>���ٌ�eVH������6<�:��
�L�I�z��A��{�r������a�>���r����϶#,"�x��101���k��?�3�:Foۥ0;�m"�A�296�3���D��<��J����6����P2]����g�Ē��UU�&1�{�/���������q�{ѿ�3��IX�ڪ6=�xI�{�� .����(�J������;)�:�*~��e��ص�׍��h�Xr�&��df=��s��
~ ��Aʕ�]�Nq@�ޣ���h�:�Ʒ<�hq��v	h5�^��0 ��恦~��=GPj�>I%%"xe��ݯ�d�� D^�%�lw|b�[Zi���t��kGB��5Z4q?����KZ�	)YM�K~��
�3D��U>�mQ����A�p8(��M�rAs/Q;d��~-c��4��Sx�iV�Ҫeݢ��i��$m�oa�s�C�܊�F�X��\�	�-49�ݨhEDAC��:��Ώ���i�\�>2��hn�gʿ��c�m���J鯭������9�}�j	��2K���^��y���d�q5ymV��m'{�=�!�2�<x)w��`��������CZ��G�N�M�x89q7~��+���e�x��XtHV�Z���D��s%
k�D�s�:S��K��3���x�U�G.�����~6W}>����̶2�ygb1�y��k	���#�twĺ�3�#e� I���-� %������|<+vR�����K�'A[]
;�lu<�/��)�Bf�eNMhgp�g�|7�f#��)�_
6?�<��5�in.�8�|�]�(N�{����R����	r{{�ҮU�&'�r�]�~����t��
8������ �uj\W}���ݧ��Y��	��|�s�|�R�VN˖�����+����~g�h,L�h���f���nJQȧPoD��@q��31��)���ȉa�id) ۇ6E~Ǐ{F8�����dC���m"�(=�3#8P 4�g��c�
s/Re��dg|��~]�?a��<��YE}o*nn�v$�[�+E��pb�_�u���C�b�4g�M�շl�^����ꕞ�,���9� Y/�Z��+�9j�}���(5_: $j�!E� �[~�I�+X`3fxD�G�QUiX�+bS?E�w��u��a��~�8�O�f���C��)v�L3�֚�9�WǓ�� *����5{�d�'��HP�Jk�����c�0;I�j��Hy,�~6�f_�<�T��'�\[�`�ǌS��)���~Nt�uBK>�^"z�w��z'�W�����JA�vyUÿ۳Ty�Ɋ4�'6�1>{(r8�J�K}�|Y�=@�<0 z���1��&0�����Ժ�x�:1^��*�L�<�����D�9u����� ����af�W�����
�|}�����
����L���Ɔ�=��N�� e��b��2x���f!����5���<��<>b�̃��;sw?�O���e�x�]T��Y}}��&��p�zԣ����0�\*WL֦ȷp�-��wXyRͼ�q���!�����_vϋ~���F���J(S�ޠ�4���ˎ��jy�ɖ������1�Ѐ������R�T7b~;:9ku��(�a�Kx\�iw�O�/=��?s��$[5�՞��S#�O?�����e��Q�b�ji��S��L��!�e���a���Y9{�k\e|����]��,���d�|�W6��J�D[��f��gƀ�4�?���N�ϧx�o`q�c�̊�b~(��� Y�πsy^,N�@}�T���j�6(G���7��z�T��-{"/��'���bS(~Y��z#��h�f�9��s���JkF���a�^��H:��g.�ԩYKqe@G�|���������H�U�ߢ͓�c'9�=�k�V�~��b]���6`3��بx(��k�5�(��b��Ɍ�v隧�R$?lޘG��M��ɍ�i�ꕠ�����\/p�ۂ(�xE�8V�Ý�y����*�ݗ�M�(W:�3��`]��>�	�����P������Vȉl�	f����g��)�����.�5@�s�zlԑ+�V=�ńJ��G��G�����Dk���9�)ҕ���;O��뤓E��u����q$�{� ~)��<�|y'>OK�Y4��NZ|��"+���v�m��'2��F) : ��Ӓ�v� �1�an�Y�n��;��Tmc�����$D'U���PF�c�r���u�6���J���vߝr_�BN=۔j<w��٦�������Gq�6ġ�� :�Q�����6*��^��=�#W�S��� ��uQ,����� >�/V�Q��_�F����`�{�T�D�/�rY긪]��
]��n�0
6�Z[|�U_�����nR�:�;kH��S��U� Q�+\-��������je�ʷ0SJˉS#l�9%K�L��A%I��	�X���LE�ʻW�A��b��<�J�Rr1�A�͊�����הmhq�T	ކ�{�*��z��zA7H�w�
>l��H%t��f��b�b�Sa6Qf�z}�=N��4Տe�=�BY���\N��{�.�ڵ���	�M����a����vOQ!��{w6yi��ַ�wa�r���_xP��h1Q�g���wN�P���}�],���,��}��SJ��-�=Ԛ�D�®�\j�n��Z���K��e�!?�q{�5+�=h9���$9]�f6��a/����/y��a�Gg�d�Y�^��g�Kwb��D�_��"�O�Ǔj}�����'S}B��C��}=����k�]I	�A�n� ,ڟ����y]��=��u#�q������_(��fr���roca$-*�	��Y���%#2�S�\�Z�!�W`��V�V�F��b�{���{�*	:]�����f9hX� E��I�7�}�	����-/�n�B���o���0Ľw��UŸt�G�:��@v��"���!�wV�5:p��dg�x����j�����(��R���-8Q熊Y_��M�&`Q����Ύm��=5AV��
mF;A��<�Na�|�m:���ܖNd�=(r�V �(؜N=v{�#�,R�z�k�?��\ET�҇r�Ο���/���=�ر���W��;�WC^w�f|�oɅ6"W��~��
K���!�	ED$��~�-ƾp�C�yT���\_~C��a�=�3bܽ�\W�O�P�� �{̡�zy���ok�p]B�0-4A�f����Rq�> v�d���c��	3����b
)� �=�\1��r�6T�#������������/vL��K�K%"�Vij�y�W9/by���Pmp�������m\A׊.&ހ���}kV���tf�,7�\'���o��1l��_��V]Hf3�Dђ�LW$}���|�W����#{2�{�`P���k�+@�?L��?�^j�Y؋�E-hd��-L[r�:��p/8�;6(a[,w6�v(�i0�뚭�ۍE��+�<p��=��_j��H(�X��4[�Q �� ՂI'�-M6�� ಟRa>��O����M��=��x|��T��\f�c��O)s���mih#���$��(T��K��a�`����\�y9���+�j���jm�ױ� �S�q��|n���R���X�Z��k�=[v��@��[�(k0*f����=��͓^|
�q�ӫ�;0=�`�>�� Z��ʐC"\I���+���|-�y*���乾���~.�`[e�� *N�v�n~�zI&k�E�sU'nM��?�z����hᰄ!i=�N��+�v}�o�}�Y��7d_��6~����M�B�7��� ��b��c3W`(4_u��q��ɼ!��0<gi�J�W !	�R�B��
�ݚ����:�?��ߧ��-c�pi���n�i���i6'�>����w�䘓(�Y���U6�A�������!����K�;���<�g��"� k�Q�����W����J��'�A��d+���{�CcF�ЂZ���yڰ��`ҏ����x¹��J�~��m|j����z����(��i&W|Y�IV�u�M{m>L8P�2�(��N�CgH��lN�$Oi�)������Bo�	����E�9��!"�)h@����:Ώ��'������IjZ�8A����u8��).*T�ɂ�TU 8;���dTr��dRr��$����FY{�Agq����L)ˊ6��<K8�����~Tt�纺V�ey8	"@J�7$4���bt�&!���P HdTi�SU�f*=b��	3���	�I>Gy��fV�\J&� 宥w�Y�׫_t���~Xf%O�jZ��}�������R��lʢS��ܩi�g��zՔH<m2�[���zX�T�u����]��G�\}}��Y���.-���b��8xe?m�H�R]b���k� ��Q��H�$"����U�'�jv�D������V�4 �T����clg9��������t���BxK����?v�۔O��-�!'H�i�ʞ����؞WO�A.��w�m?�K�,:�Y[w��+�\b�*�����{d�+�� ���ܤ��p��R���Z.J� �W5C蕃хA�s��K� 1�2�-��SD�v�oF�����lǷ� Þ��5�������h�/���"(&��%o�0��[���J����B DR�J�v�f��i^�A����#��P~�Q�5wq{RѼ�x�?xѨ��Y�ZI���5�v<�ʒp=�zЈ��t=��&�����"��Y�Q�S�EKf݅}��|
Y|C6����"V���[U!���a�NΛ�aMyȲ�)?�<�2F����O.V���&��\�j
��cV��;�HAq��g�λ���0�3�z��ow�1��٧�F�����Dh+�ЈDl����Z�wI����O
Cu��1c��EU� �	�	�)�oX�H{����-��Y�as������HF��G�b:��w(;���)Fn��H2��:�0h�
!E�̞���K�|<aX����eF;��w�9��f<��[C)�|�S�Қ,�����:^F"�ƞ��*�w���1��"H�2!i�p�<
_OT��p��9z�>�?=���#Gq/����U����c�1�ἵ@��7�8��.wQ��B�t+攝ЄI}1`[�f�����)������w���e����O�e_���m\�Յ�&�"y��<��+x��cA0�/r��0�O�)�WH�W�%Oԡ�][G�~ou��n���!�:��١O��Yl��`z�$9����i�.�
c��m�B�GH8���˚x��％h����������h�Y>���Tԇ3�=��Xo��Gg B%�;E����/���׊~]o�^���{�Hn���5����a�\��ϽlB�^�'�/f��x�Ж!���+�	j˩�r'�ZW�z"��8\o	P�I���>�! ��u�Ө�*�Kq�YW$�6oV�[�Z��&Fp�#z�E��56�'�^P��`���{�$A�
B%@K��&Ɛ��V��2y��mWw5�����G$��1/����c�x)�/mu͟��&��	�y��Q��e;��Mq
����Z�/��?	���	c�Ќ��;,�DϢn!7�*�vx\���&�GGRq"7�b@�i��q8�o&i�0Ѣ�q�M�@;�@��y�Sd���`�x^�K�Z���4�E�Y5�j"�u���"R t�@�P	*��|Q��n��iQ;�P���4޷
G����,OgR(���)s}1 ���=�������XoI:�U�<\��s�q����y $�/%Д�.�����z	��և��#B�snX���U�<1�i*��q-@\���T��E$ !�QVE#��^�7c#ǘ��$���r!�Ay@[��K�����
�'�A����2O5T�Y'D\�[��4c�'a�OSf�<����h]��l�P�5�'&�� <�����̌h���]�7NiI1��f��if����Ϻ�kd��.��K�٠��E��>��-۰6�9���@A>K���CN�q��B�ej��2��y����zY�xR���s�[3An�q2F���#�������8���4����jx
�[���>)���:��eX:�%�q�s�bY�G�ӆ.A��t�(�/�M~ܹݽV��N��Y�79	geM%9"=eX���@�#�=d�7#8a�-%>�Z�N��8x�1۵xb5�bZ�K[�����,�L��<u�Z�7�C�+�G&(�������TÌ���jS���{�熮����<N���:`e%4��Faha �G�h���U��{$X�4K<�o-�|�C�v,0[a41f6����跕w�@�C��'k��7g�1{Dw�d߳��vI�k�\r�n�˥3��{	Mw(�s�zjfVz9u�:ng���2*�t��J�r�)w���`K��hE�Ϫ��#��2j�ȋ�k,ӣ��Er�-*_9W����7� ��fO� �M}�&D
��~�'�D`v���[���0<��Ն�YN6��ɱ�(@Y�~��T.��'�Z�?���~@�����h� �&��AIE�+^P�՘�t�����X2����9��Z���,D5�V�m��C�l���q'N��jr��A���9^ʶ�qn�M�C�����q���7d4�D?�-Ċ��jL"CX���h����J����[$
�d�Yf�@bs[����/	�M�NU(�p�ib��ݜ3�>�7���҃B=!�A�d�_TVH[i@��dFI������n�B�b����k�M� ���l�Ə� �h�e�&d!�A"F�`�QBW
v�*l{:��ɚ3dF�x��b�`������}�U�����E�}�Q{G��?|� <��G�?��|�)O t� ��m�&& ��l�(b<+X�d>�����=���JH�|\m8��U�������@½�_3��K��3�i��|՟jǷ��U�?ڴ-�3�6�@36?k�t�"<�'����4��0.	���G���7�ƕ�3�Xb�\3�p�� :��N��X2<�z�F��?���`rw�"{���%�#�N�	�7���&��o����6���ґy�����k�*���}�o�[.a���ٝ9�I�+�,�{��K�����6>}�P��D ���������U��-,wD��5�ћo�"���A3bx�Q�l��_�L��Ս����6�-[{VAO�$��s��2Z�\����Z�enВU/W$c-[iV�˽9kY��!	�U#�-B�HM,��i�G�S����x\8y�?��� �<A���,u�f�0�?���3Gʃ�6�c���3�8��F�c�鞇�����Y�	��1-�P0{ ��퀍�c��\�҂J����B������fX����[LX��Ǒ�v:Ur|����IF�����p����i̟�`��c!��I� ��<iZ�T�`�m&��<w��/α6
�->5X�u��i���/��DQyo$U&W=��+0c:�:�4���7�㙯\�%�|�B�	�|`���Z��1-��:��3T~���:�Q2bc���,�C����^�:<W���Ğ��4��C��/pm��0�ݹ�?s���h��~H��Z�`�J����tݗ��)�m�ϭZ�/Je㉷��"'3��fU��4.-�-IWħ	��&�7�{��8�
}ʃ���`�I�r�4L,dW��q�&�B��m/aH!�)w���f�(��_��̹�~h/�Zp��G��d���!���*�W17�h8�R=�Tj�z��j����@p*���Y�F�9'S?c.]�D<�
���X˯)Q77��3�}g?4�(���-t��~H�Q*(y�Ǐ�ӫ�7ǖ�_������6����S>SUͯ��--���s��=n�Z���j��AcT޵؉lX��q 㿠.�_��ڸ�/1�4M�h�"�׶���B���L� \���9˳�v�X!��ZM��&R�)��
�<�?�ZF!�5cr9�b=��k��g�v"�l�۟#b�b|!-�͔�䬤�D�B}8��ɩ*�.ئIV+ÄH����
����[i׽�0��s��C�XA>J6Xʀ�[�/"�+ʼ�������L��\���W�ըj`)�m B#�4q�� �8�3Y��wF�rU�oc{?���ޣ���C�ɠ��dwU��� �[�
u��F먭I$�U����^��'���.%�+b�X��Y�߼���]8�#�S>6Ҩو��#P�fU~&q#��q{p�Dn����ɘ���t�eM����c��U�.�05H��YzUl��-�X�6C��˛V�pn$LI� ܵI���_�Ĩ`���QEE	�Iy9N{��(Dۙ��w��$���W#uVs�jF���Q���j��ֵ ��݂�[��j=4�U����-�(�mEj��Ho2��sSib(��p��硥��ڽrh�O�cobq���Ϭ�dls!�$����yy@��U��~MG��eu=x��E���'8�7�����uk�)	V����"��ٌ���t��҇=`h/p�\O�+�N�Ge���<r��*�}4T��5or�����*�G�[����Y�d�{�{��RTS�q�Q,���e{_���3Lp�g�ȟʸ��&<r�\-��%l?���Y(Pg6�t	������F�[�2i%Y��F'�]�L��5\�����❹X�xY�������ٍ���膫�A6@8�K���#'�ź��gz0`G��IE�f����~}ؐ�%�r���e8�����!;��Jw_��B��"U"����Z�~�gC�	�Ul����;���(qZM�j���Q)_�h��sH�z�͈`c�۩��IhQ�P*�5g���"�|�^Φ���ַ
���+�r g
�"�8�������Ak�/��������֚E�_Z��\���>hvUJ���E$s?e\s>0���( U�7�����8^E���8��^u� �)K�\�S������;@"��4"��]�d*7+��M9�߿me�)�$�P���K~wr�T��GOU	�K�����a�Ã���^�rg4��P�9F8u�����d��V�hi�����q���y_�<��!9:��>un��^*����9�� �ꆶ��|NE�>$�HŅCv���D6�ޘ=���K��%����B�^|�?dr��u������B���!�PXC��9�y���1Z���>�[Y(U{E��S\����~��j��	����5�֠�2��0Wq:9����%��k1��
b���:ĒI�L��T��6��g\n�HI��L\n�bq��$Y;?&X�E��B��$�M4���;����7���E,�g�M����ݷ>b�S���aJ9ѐ;bQ��6�&��ܻ#�8�)���O�I��{̜R��,PوDl#F�3�����
����v��R��ڵ�M�w��Yh0�,.����o|q���f��"�������U����)i�]��/{�H��%��F_XHj׋�/���bok����Qd��k�^��a��pcT ���%��?%R��DSvB��p�������d�ۗ4S��bZ�\���0R/�'�j��*��㢴w8�W4��sS7��'��1>�ЉT3��Q�HÚw�T�ٰ��D��J�A�۱]�҅�%��ژ'5�Fu�`>��
�݌�1�y��c��(yEƺ���mCqM�(�
�
�l���������Z#��ϋ_ҕ��lU+�(P�g�@�dz�7���6x�]3.��%K��G�c���6�f�8�B����FJv-�Bx��$����g�S���N'������I}h�8e���5%�`�����`���9��w'7L��p�_C�k�R����d~8��
]97��0V���8��P_���b^նT����W�#~nE�֨��pD �> ԗ�{iU~J�=�^ҠqB�q�uNS��V��9n>1��Q]��<�#�^�ǖ� '��6?ua{�P.�yc~��)7h�Q�2��H�T�/�����`v��h�~�*���}���:]=Q�%^J�%���Z�x��7/5���O. }`��_���g��BX��W��WUB�!P�޵���S��Ğ�kN����.�T�!�����ZV��R���6^5d�`�=2+'[���/h�������mODP��/%t��ỹ�Ʃ���_�+唷p{!3�ꕪk�c`�a��-Q���v�9�|���X��yE��b%�cv?�W��%���)ѧ`���I=���Y<��W8��FjZ�^��$�"4Y���H!��P	a���G*�~��'0��+�5�Zҁ{D�����~	[���z��e�^5�\��`�q�b�>�*7�ous�|i��p�������Mjn��3�.��c�o���U�g�c *pIu�I?g�¹�v�!�:/Z|��*�a�aH��B���.�z�5�i[p��?�A��ٖ5N�xu:�$�]b�a;��Zр�S+��̀9?c��DB�u�8���&P FU�o	/i�`d��̑��B���R����U���I�ϟQ+�S���=r7����u
\]�fI����X>U�_f�=m��f� U:e�@�肑c��Q� �	��bfۿ�m28x�QU�}��P�gVt�8�����3�Q�q�A�ˬ�x�)��y�c`���$Dà��l�g��ը��I�M|��kX`�Cp����ιu�1�����LK��8Jo��_��>-&(Ӭ��Y�6���N!��ٻ&�r^��D�c4�B�mT��oO�
�&���/���߷$'��YU	����S]~��xǽ���/�Rep�Ca}fs�ǵ��fN&��9Z(��P�:��j��;��^��+��m`}]FQĘ���j��B;P��?đ�.ȓuU���OW���	� V?�_�r�G�E���@��ɜ:h�q�v���]�I���/˔n��˸�)<�3�{�N��y:���@�l�զ���G�p7!��jlU�˝�?bo�]�������Rװ���o�4&��d�ɻ��oFޏ�>�8ݟk����y�_�Ii�$u�(z�i��*q��1-�+��'�S��ڔ��n�����Qrϯ��'��
8C��:~�e�̓�Qō�|L݂ �vsLb�	C�,���f]k �vm��ѓ�<��d+�/:؈-�y�M�Q�!tG�L;?#��{ ڹ���7�*΁�;#�PO�8�nl�3���PaR��[V4�����e�B��4l;fk%�O��2|2L��}�z~���T[�9��9V�-��/���t���(F�`Q��6f=� �[��d%s~�g
�,���I���,����u������:`��@����۶�A_�l*u#�Y�nEn���P������ۜ�ȅ�u]�i�U�x!�r���rr�f������4�6_U�Զ��ඓ`{r�U��¡��Q&$(ǽIQ�X�2֋/�
�������=�bq'Ê������3�����s��������� �ޫC����%�zm�Ʈ�����Җ�=�{=�V;��08[�0�d�s*��@ao��ZO-�2F7R��}I�di�pv��LMü�i�)#>�p��� ,{��2D�8�#�"���(g7Rq[�G �S��$���q�N`��JT85��c��K�\o�p��ii����y8m�e8\�+��g[%��M��!�]VQ�2��>�u���1ߣ��0�8b%Wk�S�T_���p8 �]Yo�Fce����*M�1��>����	���~]�Ό��$D� �ή�R���GH$	wC�_�d���s��)˄���%�<2�a����0����*�qY��"������j��~
�6�fe��0�׬F�EI�K��nM=�N�)t���G���X�
ԃȟձ%8+�+�|z]�3�H���L�B�H��å�C��#�G@�nr���t�-6d0�T}`UesY�� U���׻ٵ��*6�O��6T�G���쿄/�)�n�ʁo�}D�)1�M��6J��v��%ަ;Um�@2Y�Ɵ"+k֐u=5��Il���;�Ѯ��xV/��9�Ӧ������`e��S�A�7�Tr'ۚ�Ø?`�/0
@ |,�!���]朮/���t
�7Tmrs��K��k|4Y��pi��b��N�]���r�ёS{�'xCN�s����G>����h�ߨ�����s@�E�Z%���1����d�6�Y��c����/�zB�ߑlXy���܀p�-M�M���~�Q�:�aբ��3d�<AQ�k�R�6?JՅ�`є��%�����d�և�;���C��[L�?���cXrn���:�R�e�<���i;���$Wˡn���H(�?���*v�b��wR�C��n��3�9t\�-7��Vc��?ku��UvIBPE>��eE�yT���#�i����P�_lir�>��
	����E�'::����W!�ϳA�>ͱ:�De�~���P
�_�1��bT��=,�ŕ%aP}Z�
y��th���X~#w�AA�]�}VtH:Ps�Z������:_R3��-\[*��7�',������&a}�Έ0Y�°˘U_(�������PS �B�߻��2�qS����
�W���(�x�s�R�C_x(��ݛ|Z����N�V�
�a���E������y�
:��Q�|ճT�vN��	�������r�$�D�o����`�*ڻ��xV(-@B�g"���*Y�+z��l9�Ř��		�Vn�t~���>��z�l.�Z�J8*]��%y��[�6��ґ9&��T� ��g�L�( �-c�Q�
I��(���޻�E1-��;�C폟
���
�Ԣ�"��%Q�wN4:��g}�S����ȿ�~���SH'�k�Kv�͌��(�S�u,������2{�#�ءuZzIn��x�_�%9`ЗA�<�~)d�骙q�Vy�u�P߯���A���S�B�	��x^x��_��Z!w�w�p[��>�l�=��A#������Q@\��/�+'�<�H@�B.��䏌U���y"�7�
SQm������M�I�R�:�O�탌8p�׍&���� 0)�Y����\��r�S�����N�_�j�T�m^���J�:���O�C!�����~|�Ul�պ�ވ��XN���'Rb����J{�?D�]�Is�����4��b���5*���q఩x�]t:6�?2��-%�E0�	��܂��#���mXN� Z<Z�@���?A��v©X��v�CGtm�ϡ�[K��^Ѐs���K��`�����ךM5���b�aFVY1�>�������2O��{�n����	 ]�������^�Ѐ���˸� sh�c"�h�s]��o��ӏ*$����x,��!omY�~O/M�Ʈ��S��|>����3��݋O!W=�퓂H���T=(��8�O]�U>���x;N��P	{)���t7	5�j�V'�%8
��F� GV�bW�oz(H�M����
!���|�&�L�=�6a��f0EqP�o�Gk�Xt#����/��$ܱ=��c0��������cO\7l�:N�h*6�X�|�P����2�"��&W�t�|n"Y�7;��:�ڦI��R��k�C?T�(�ze�!������h�{�(A�
�~H�*��B�7g�Յ�BK72��I����A������D�Þݛ�;�=�H(Q�_ ���q�(�F��b��H\���1���!"��$���]rs�}8�C��_Y���<��L5Ҏ�t?w�Թn�SR�U.S�*�kP��v �Q�iEߤs^Q�1
+Mw��?�Hv�ߋ�w�
�E��4��c�q� w�0�T�3>�)+�e����|d-I�4�R�$��Pz活�'х��z���|@»����Θ�e��I��vp�0;�hi۩��ܗ�|�""����ڥI������A߃Y�:,Q�K��Jx�+�1��&j;v-1a]h0�<cF>�j�!(�0�_J���S��F9j���+Ir���$>�XF�ژ�wYs0�����	�w4���R�ɘ*��0d��	ݺ���R���:u�:��M���a�m���l/s���'867��"=���{;�K�7��=V�:f�%�k�߫������~cQ&���?���q��Uo٠U�>uN�^]�r��&ܮ`o��2W�Z��z�<�sW��)��"Рw�b���O͊-�[nZ˨"J�؛�?ڴKnuϗz�0�)ƣ�m^z�6��|� �wk$]�\W��L���#Ӣq���B(t&X���z�Il�=E%��X���@��#��b� ��M��P~���2�Zk
9�#�	�-���]oΑ�_��xfy�.�/��a�b8�������#�ZC�l�=��s|�V(��I����<t#q��<@�B��G���G�9��UCo�E(�[����r)_l��!����
�!ۛ]�qw8��q��߈? ��o�݃&�Ռj�EP��Bj���I�f�^�xA�~��w�a��~]
 a���Xq�>����\p�wI�v���*Jv����t-�蒶�9l�zRF�A��2��67�������:���Z5e���mRp��S��awf\S>x�Z�^�	�+i蠤���
B$VR3[�����2���$`�v�Ѽ���[3�������>�\-@��N��.�*�{���/�&	�B{U�������-��'9(_��<^��ɴ�Ɔ�^#�쩤׳lXV>x��^T�m���".�% ����^�3:mH+��]Aw�%�T��N������H�%��׬y��$��&����c�8u���a:!i/Tq@bՀy��ԍ>x�4�]Vtt�쥛�ѕ��+{h�MF�q,�F.'FTca-�T��ۍK���5UJp����$�q�Q��4q�y S������G���HQ�)r'������$���N���H���aś!d��__4`j���<� !:������'�!�p�dv��~��D�\���ۃJ�Y;z�g��0 <���3I�j�r�8\=^͌d@/�R�F�Y��Db��yݴ�7�\$�d�������G��Z��&�FD�̆�
_`�u��,|	>}U���1�&�}f�c���!ˉЙ.���i��u�͏�q_�1�E� %|w������}�Z��0��&��4� |�[.݁�;����Yۿ�����IT ���^�7�O4�G��id��H�8]:���|����[�\��D�L���)Y%R`o��zC�*jh��~�"5�uD,yx	t��@G���N��#֛��6�ѤrQ�f5n��C�suy4��Ԑ9��l�5����eC��G׎�Z�~����SE���c�כw�������\?��!�?�ۑ�E���]�m=[�w����.���<��(�`u�ի��9��Ⱥ�=�h����c�=��$�H�%B�[bԤ�u��"�s�u���,��3���6��l�;�k0�(d�Tz�����9zNb}��8���g��ϼv���R�B~�XW� �|	ZQ(,*���,��v�h���ݭ�U����s�ma�f��l�$v�C���$SG뎧uz�I��V��1s1ΐ��x�,�Ff@�����0�I�F���$O�g �tCH�"_*�"�ckڡ��[��x�0��&�o���+O���8(s�/`�m����V٢6s
יJ?�a�y�ۡ�^�77+��Կ�����"`�lY�+���4����/�y��y��ZN�w�uɢ*����ط���r4�?��2���k�#�v��.ǩ7ԥ�4Q���p���FH}��7�X(StTJ� |���b؋De[/|���a�_��N���	��,o�V�YQ�P_I�2�č�%�9<m�Z�����d[O%_��<����y�*���m�|�i�N�N�=�GS�S�*� ��vNKe�	.�[���	�x�!��@?� n6�T'��Y��F!h��h��J���ks���g�����>��G2B��z������j6�u0�[�d�(]��P��SC̤�	����E��L���8_�O�J���i:�_���'I��V����	������W>�g�Kt��+N%V��s��A��Hzՠ�1Hs�g�:���o��5�`9�Ѱ=R�F_�&����Xv @��ޱ3�����婇�Q�:r�&��Q1���G���.��#���|������x����W!|ѭ���,K��G����9k�%�P_$㑵���yj��A8ܫ��D��̐�4c���'I3��ĄN[�޺�6.0r������j"|����뽐Y@&�lZM퀉�-�O�W-�F?i��;t��EA:є ��^��yG�vn\�-G��M&���`���3,�H�B*cK9��4�[���^��F���x������jT]q�Hs��,[��C�?��x	�+��q�.��=m�����]�[ERR��Lĭ5���;[}P�ç��8;�O�Q��z���aƄ�{z.�_��-_!+{�w)1�qY�+��G�-��s��� �D �Nr��k�<�����yx���4��~6+��(�!��BqPKDr@�"���ԝ��<�#�8�Z?.:�+�Vi�|F�%l��A���W���=������H.��"��#t�;HC��1m�=�-��lԺ9�PM��,����!�-���36�u��	e���"�k�y͹M7E'
:������jw_���'Q�n��8��+�b �������|�tĭ�L1T5�O?R[]��~�^l��\��(��pgu8�g�,m�(�S�E��%r0�^:�g��=dY�$� ��W��3�Ɣ@��q�[J@����&�Әk����ʧ���Ftl��B
5��3$6H�"ׁ|*��g�3�+�t����,[��ɸ�v�W��aW����I׿w�8�t\(�D�*ٵ���Uiɬ��U]�!���s���[��b(�I�Fպh���߽$*��[k����:O��[� �qs;�DԀ4d�ЯT��_���d�2e.(�]Z_���'~4�Nl���(���1��[-P��K�B��ɲ>P��yŕu�K���6���u�֤A�&2q�Z��|e�51�k(�� r�w�?��J����x�i�V;ұ��
�,�*P͝�5�$�6\���C�mi�9��ǎ�a�HB`��P�d�:$/=�7�XqIC�X8hN53_qJ!I@?;��:`�0��;ص���K�|�b��i ��?�u�/�@"�&���gw5��I�J�`� �{�1n-�y�}k�R�d6�C1�"��J`B�h�Vi���Z�kS��$(6�SFA��J��Q���t	1p!�� `�U��N{s@������B�&���p"G6&��S%�U��&��O�3��4O��a`��4��$��va��jy��`A0�'���2�>���b�Շ�Rs�EVʄ��@�~}�β�ʰ�s��3l��	a�Jfi̍����|crɪYN�$͐R�.��ބA��놢d��&���15��������`�M�\�4�o3�'
#����K�S��U��qۥ�2Cא
�$����íA�F=��[�����;DQ*y��� n?$���?"���g ��7?`y�W�Fm�hW�H���7u8��EΥG/����>,ٌ����P���!�{Z���I
?�@����B����a���~�;� Q�͗M���$.]V.����f]8B���"�p}t"�9c��XAT�>��eD6ƒ��]��e���W�q#[;�6SQ�	�z\�+-�9i*��*�����g��,�> ����_���׸�f �����6!��Xv��N�/����p���K@ITLk ���i�.Ω�<H����2��bJ�������WDP_0���)��h�WNƷV߾,)UG��g��������C6�D܎(!�=R���[��������b�l~V���x֣��m�0|���4ȗ�J�uqw��ǘ�V;��@e��|���m�L�r۸zka� iぶ��9 ḓ���Y����H�9��������K�)��_�/v��������ꋭZ%(�D�k�(���&�e��d���j�~=���ץ2��k�4 ���f��U�]��^� Շ��W>�U��B��jx�)��LR7���Eh�*�F��FD%�L/c^0��E�;�*���1%E��+�\�c7,)꺴�u�wZvH�e^��b�U�j��i�9��"��t��R�����&�"ЈD�[w�t�P�c<�"[Zg�( V_�ZȖ�Żh<5BS��0�)��堬Ȭ�J祮��A:�Xk +~���9ގu�\j	�xH�W�Z�8D�Gr)����A�����0�����Ԕ��֠*����<�Ч�������L�n���V�j5֟�]2R�ۿ���|#kH�����ئv&�)��_z�g_�R��Q�*��{��+��gd�"�}�[&��lj�Y�N!�4�n�Nx3�����`EtO�yg÷�3���St�F#��r �����덙K]��Eb��c_�S���ѡ�j�n¡��}�@���uɐ#��f��w-���%%�Uki%��j�����.�x9�Ӝ���jrc#��8��	�r⣳n��*W��f����I����	6v��pj��_��TN?ׄ0;}cc.�X���7.҄�� ě��5 |��O���u��򓚔Ҧ̉]�����$�OX�*ڌ�c�ީs��X2�G�n�J��'%��yc�a�=�]T;V P� H�:���x��X����"����l���[fS�H�n�rNPN���@+ő0�ן<q\��$�����i<f}��y� �B�d���*�N��0S�exo�Ŵ�ȺadSv�o����(7xD�0�Y��M���I1�=e�V�u�� ����J���m�WȽ{kE@F���sM�Xx�>�N�S� ���L�r�t��4�_��_���q���M�.�B�ְER�b�B�9m�ƀ����,�+��H��a�\�1��e�>�
�*�Q�3v�{MD/��=	G�{�Ԋ��/d��3|��D�����ə�-/+���0�L��I1������$`�zu�
y��z)����<h���\��Ȕ�"�����W��R�UA������|����4������7*e�|V	8�t�_����4�ز��r~)�ε���VDz��@��Y(@��� T�~b]����a��7D��-��Nψ���J{���R�0�e������������DƑ}z�"�m=^�=���M^�T3�x��b�����Яb3�K>�>�����s;>�s8���ck(�?z�*���p�y���kK��ȴih]i&M	�ˊ�ʖr�>��gj�z�2�G[��kf���٘Жh��Ҕ�o�Zvu��Z�P�����v":rOh� �@�U�N���z��vX�A�5��s��5�0�'��-�4re-��Ӓ���O{����.�k�r�����<N ���t��CT^i��b����n�»՚b��r���fm��%��}]�@z�a�q��@����O�˭�n�pCk�ί ���]2*��[ie}�\ڊ3��p��_;QQ�K~%��	
^��!qe����~�m��0s;�cb�g^�+c���\(�Zט�D"л/�чt��#�PW���0�]I�P�i҆�������	�)�h����l��uҊҜ}�ny�*����e�r�4.��0�a�� É&�>��~�d�A�67����= &�a֠�?��'�T�{G�,u"���,X�z �'~hPEP�{���H�. 5C��Ig��5�� 	��!��d��T��Y�}��w�Z9�{�0a�+�C5�%�ģ���¬xޗ#���qP�B�'��?^Ǩi��%��r�G�ʩ
�6�.�����(+x&Jb6F�ٷ"|�B9�D������͠�"�w �4Z+�3G9����;h6Ƈa�E��I>�c��W�$���C�Ġ�39U#�/wc%S	&%�a:)E�m����#�ɣ��L|=��E�j� '��V�c��^r]�� įˋ����ӄ�&K|6��J����гu�&=���g��݀y5�+�w�! ު�uP7=K=��b��؏z�(\�jF�B��Z�18N��vB�Bo�y��T�f��?T��9��H2�-נ���gޙ<�#�ݗR�F��o�!��f3�+]�5�yb��%�6͸�.�̠S�}gȻ)*y�:
S#�6KPb� �G��H�/���%���ѽ�K(�?-�ׇ�1몲񘔓%sE�fK~C�t��[�2����'�['K�8҂�L�,��(a�]P♇�� �G���D�p�<���u^��U�ʥAF�}�%�k���HD0���l��ҵ����C�7-�R�`�GUN��+���T/R��G�J��L���[�j?��ђ�%�v��xg��j�'�:sz�F�R�s�ۄ:���a3���J�����ߙ��tt�/�ٓb�=�d�y�y�20~z�E-�l�2��팾����}��q�J Wݪ���c���4%ǰr�v��l�&���+�ʷ�pL���X��n�&t̼���E�5␉f���9�s �z*��֮wx6�����y���ZS�EϦ���mɫ��?LGш)�KZ�J�I5K }m�̒F�M7>���|��h!,Gi�4Ǳ�{�"ʠ�ۈ�R����"��1��C�??��6D���xML��|��6G@�F��{m�)�ٟY��.��>%a�v����G^ e�m*�ǐ�Nݬ�p1�0ѲŔ��)mˇ�KC�m��Ll��}�s	�_kǶm�Z�$�B	DdC_E�>n~��ٯ11T��V�elbW�c�#J̣@���Qn��<���?�H� ��T�&z�\�}:�V2j�;6�
�W8�w)�^'pJw��9nY�Z�m� h��A�dhz<tB�S)��BYMM?�w��ш����z��Su��F��Ϩƀp"��y�E?A��0�yΊ�Pd���\/���5��r���x�q���NЂ:��;��7�����ʋ�:��g1���9���`U:u|��Ύ�{�'��.>�9�_����Cgш��V����gj��];"���!��~y̤k�7� ���7X,RbFf7���r�����w��*��c$�|?�D��k�י��r�}�N��IU�:��#=m��$����NS.��z���>k��$�:�gL~�y6��b�!Z)�K^٘[K�ܹƝט_~n�^�H� ϋ�0K�t��A�B��^9D���#�Xo<���$�>���"���^`9*��q�����8�8t��b?]?�,.��B��)�_1L6��(V�	�`O�}�)$!�M �����I[��+t�pu<xd;о�GN3ʾ�#0Ԃ�l0�/EΠ6^�8%�A\���׭iR�/(v�>A�ݡi%��T\E���k�ث��o	:m4Xt�e�\�g	����%��,��G���vn��p�Ԣ���N��L}�*��AԐrw#@��Hu��(�Tcxd��Ʈ�G���gy���f�e3d#���T����WhY3B[�L�ÒICX�S��m��#�K�I//�l��4�+b�q\M��\X�,�Qx�"^H��yӸ����M���A�J�țA� j}2�
Ʊ��Ə�R� $�3��9uC?D�6�#D��C�P�3v�:���Rs�ʫ�@��6��\xH1�C��J[C���O�ۀ�'��=�p��W�ljBh�Aiy�%�)�I	�8Nq[	�P�@+~N ����^�ѦB߭}�h}0��QH(L�VA�C�W{w��Y�����so�0&�Tj��S��cV�~S�e$�0A�b4A!BK2�N����8Қ���fp	dm.��~�׸����KvLpC���7!�O�UY��)��7�pU�Y���A\�����L�K�L�=� �)4 �;�ޕ(>$�GTEc�1⸦w��{h!=@� \qSER�a~�l�:�3�ީq���׆�i�3t���S��ϸ��[�B|?�:���8ߧ�t���lk���O	�D�N~nr�d�͞����+�O$�A�K�e$�c}l'�˯K��2�:�+~(��������Q�x��:��o�5"	��~aD`������K�x��5�i<{#L ��S�5P��AZ�E�van��e,p����n��{R�g��E+�"��|t��c.<\��K�!Qԑ2�J�Hi�yq#��'�xޯ��ؑ��.ܙ}����y��`�:Va}!/�%��1y�t��w��@V�a3zI8��mBY~>T��|T���<�2�4*&hr|��%:�0�u�B5�l������!�z���CP\=]��O���|�؃���z��S�lp�D��k��ۭt���ȏ��D"h�[g��6��9�Ia����  ��i"�J��}M�8\<8|g��<�X(�B���8�5}0���*�Kv�6�qHiW�.B���z_�\v��!oA4x;��U���U"�l�E��d'Â���h�l��j��L�)p��	Z۹�w��.{��u��[�,��<Z>��C\�1�L��,�!ᕳ7��kg�.]��.�s�9r�RX�1��b"������|!��aTL���t�C�IQ��6���"�'}X)���9�Ԏ2A`�Mn�Qu~\�떉~������R����z鱩�J�˭�qTp��*����H���SӔoM�#�3C�Y?��G��b�f���6:EA��((:ZQ��!���SJU�����`K@�*m����#��C7hښz$��7�3�u���AQ6s?���4|��Aݷ�I���L})ag�M�j#��
B�k�D�N@aS���2{5��އ�,d\"���n۩������7��g1�,?�,�%ʈ����Ȕ0H��d)حåWtP�`dM*�<RH���±�����PqO�|נ{q�9��|��aF��>)�e�3��Z�G}�k���`��ϳC�M	ʺ�@�)A�
}��%��A��O�4ᗠ/8�ړ�ʫ5(�9}y�V���N������l31�i�5���arև�R[��r�}$��01�[^�3�G<0t�%��ȵ�������MUMFZ��X#�?��&�8`�?��t�%��!U���R%ƛ��|�y[�M�{Z<�������	��X;�k��A �Ïf�=f+�q��s>.�[��A.e���(Y�"E ��'P0��+����6NPDʒ�x��&|gO�R������ʤ��%���u^lo�LE�@��*:�6�U��PO����`���7���-���E����D�:C�i7Y�F�����mP"P)���ȕ���rr9MS��glt6g���;ԙm��WF�^��֌�CUN�h�
ԃ�[�F*��O����v5b�7�/���oCQ�+�Α��1�"E�4����a�Q�ڦJ4Ց�fal3��?0�_��g�%�=�Vw���~ �Hw
�r���_?�?��@���+r7s�����G&N�_و�tr�LM�W(bR�U)�5�2��˫��/y��ݰl�p^ã�͜���@���P��f*�R=�ǉ���W�ME4B�m�GQ�L��Y|�U��z5��.裉�"�8�EI �3n�cI�"ؚ�+���x� �a7�О�Hh��&Γ�aץ=t��kY�n�i�%Pf�&Fo����Tֵ	�
��]鳾��eD(�H�Pu;3�U}���
�łc����zt��,v6�� Q*�W��K;��΅EBܧ�%�������=�iJ�jүX�C��A#ҟ}_�46�Qw�����=��q�n�738���wϘ5<�y`j��}gR[+Yi�Lz�c<F(cHS�{�6?˄�ߏ�(�h�ڤxn��>�D����'��LMo,O�ӿ��Ob�������k�
F���R��s�b�A��֣� �\�%^�I]��>�����H�$�Ku��oB���'5�[��.!������M)dN�@�'!I����H�'SL��k�'�&�YVMx0�#{ˡ�i7KeL��x{g���m��X����ǆ�"�௯��)�Ʉ�͈c�1*(�:��o�0���i�O�6����W�ɝ��Dc�BM�r43({� 뼙�щ�ͱ��B�a��FE�$|K��x6�&G�T�nh�HiL����ѩ��Ε�{�����q��!8�L�Hgvթ�΄c/1,�E=M럽M˹�Vù�F:n\�.��yX��#�׈Ha���f:7�U_�tq�9�1�n�C �K?kQRH 0_8� ��������w�m�`Ϙ�-g�' $�{ڰy��R����dɅ����WV�b�S:�\�K ��K�����䝆��)o�d+���u��6�Nwh�Op��R/��W���3�ɚ��/庺��6�klj'x�E�Τ�Q{��{5��Ȟ��n[N�m���莦��`�������q�e�*_y��瞪����"�C\��I��Q@t���a���r���i/�(	�2;�X5��κ�!S����:�7n���@��]�bMׇ�ؕ| oa����;0����A����K��s�o�<X��w�ݔ���Q��$���5r����V�BO!�[Y<P'��0UQ<&�9���\2�i1�S�Y$�ͮ��)u�9e����q��.��=�+�Ϡ�M�`1;f���_����_�����T��1R^��r�p�����Q�~5e�8{�z�а�U���Ǆ�Z��+�A)�y��40��㵃!��,[���T'y��m6wM��HR(�����r�8�!_�j�,/��#�_>aJ��n����#U,��LԲ	��&�va�����<
��|�r9��Ӫ�zQ��w��ak����foy���'d�v9t��5T|�PR�'����~�~�G��V*3B��J��2s����9IaZ���&B���	��W�`�{D	(��u�8.~�����ŵ�XX?B��tB~%`�K�Ћ-�O��p"�ZF��sך��S�L7�_����N�XNY����S�[�|����N|{@�_V��q��Z���Z,IXe򝹦lD;�>u�%Nx���sJBoO_$4U�P��v.vƦ�y���l��N6s�]�-��.^���*'�-�E���
L�h](�I[7�^��4]>r���LW����${�>����=(�˅=`O��,��58��1B9Bһ�����;�l�o�E���&�%�)�'���}�U7$E�}:(�d�� vX���=�(N7�xf	�aBm�`ڎjVj�)Y��kE��W�D��O�;�b�����-���y���ຯ� ���@l�$��M(�k��Nq��6�������M�X���K�+ip�
Nd�\)J5�C��!��(��� �Y���ۀ,H.��g�VLR��6Hê7`�'n'Daj�T�n�?
A�_g�Kt����2dev'}?����s��_��=��o|�]W�
a�s��U�B��L���#{1�p�!�MN���$:�vS��Ś�n>|�t4ʢ~�-{���o�SϨ�[����@"%S�i[=����_���DKMI�ImgꈠH���%�)��W�q�+��x9�^H
��$��T9#�g HT�g��q�=U���'��m_o�?W;a$O�l�#� ��m%s9���Ok@�$,�q�cD0��&��,�:���yK�LrEn*P�"��/A�c&�M��q�L�2A7���F�x����t����L�f�ο����}��o�
�t��>��-n��CgD���[a;�<�s�>����C�l��V�=;���Ғ@}P\4}�9'6������g�����V6��:Z���f��OL:�5���L�M��$�6�ǵ	w�#��]!��"3���H�ǣ����4�i��~�ɼWS7�a��?���8���J�-��+��o4���@�g/,)�9E����
��]��M�3��X]�$P�����r��[q����l��I�[rP
X[�a��*z�t�xu^ge���H�l|4g�{ج��4,N���w�T����-ͧ{����b���>ِ�~�E!��#F�(���2�1�Uo�3o�0�m�>4�;�ꆛ�H���8�P���p�\��w��,�gY�V:!9j��9�O�>���Ofal����v��<�tf�4��L�$#��c*�4�K���?,�lH�(�}�M�|�J�1�u��~�.��K@�	P�t�cr,a��L9`d,T��5�����a,w��'h���n�?k+�I�0ʍ��I�C��AKH�0��ݫذa�Oc¯���I�]oD�/����zff��g���G)D��̆���e�d!��}>��Z�]��`�򺔩�~N�담Ҷ��&����-Mq��YY�^��u�Fi�}[�ę(�6����,`�?ـѭ��rjȬ�����֔�x�:	�I�{ h �L#X�\Z	��]߂���?J\�;�3JۍP�^�{����r'9-?�U���r����a�;�T�cҍ|���/�4%d Y<C"�;�q���zb)��$�$h)��Rw��p�W�6�>���#u�>�Q��%���O>���膬��E�{�d��Ƹ�+|�HN�@ؑ�y�^X�sV�Lp9�����YyH��N��;�3,:dV���+�i��畏`,zE=�/�fe�L�������\���(����0����k�&xg�-�RƼ!p@���.I��f`���l�d�T��D3������9������÷4��{�@��G�S��^V�T+8���D �tv
�E�D� �GQ3\��4m'�S� <1>�E
*�����6������Ym�ا �_�N3M8"կ�܃2;�ria�H�M�~nRɆ�!6ҿ���0�H��H!UV�Ãw7P(�oR�=�zV:�o��<e��L��H�o��Ѩ-ǈ�lG*�������~N��e��A8�ߢ�����`v\/%�r��O1�����d���M%���]���%�<Y]����ܶ+8��E��ٛGz���۝{�iPf)��w\���ɦH��d��E��l�wXy9���CpZ��*�3�eb�ܰ���|2\�	��x�Ș8�Ph]��n����ͮ�Rff��W83�Ƞ^�^�"�77J�M���H�w?���ҐU�X��o#2��)\c�!��1�Nj�

*�`��D}�^���(��= ��xs,��j=ڪ�8�Ѝ��+e�T�����^>a�#s�(v8�4(�Y��e�B����ׂG�|Z�^�巁���]�#.1Z?���.$>��p$�����6�|�7�L������0%[�	��nˌ^��F,T�^)��YG��q�L�-��t�0�ƍ*��-Z�
�����x�g����.�NPBQ�ҫg��U��n��'��M�6���J9���պc����47S1����)�Б��C1�{���}m�����̛a�`��ZA��,r9�v��o�����1éM�9:���q���n�v��I�	��tU"~-�
��K��9�E�U�vD'P�8y� SC"�ۜW˥}���͘p��z�w�4���>Z�w.w�Q*\(���$���rZZ@o�7�j�|;cu�<�t/g�s5s����_/���=�eZ�1Z�h}�Ah���ˏ���K^%��!�_V���c�N�`9�����j�� ���1��b��l��9Z�`�;2f�Jܽ	����o�\y�E�����R�2v�/"^��-���y�$b֢#3�m���@��Q#VnY�'�x~Z��<C�p�"�Ǥ�[�߯%Kcp�T7>�F<��9�~@3����%'{�:F.�/:2�b�*Xۮ�K�%�C@饀��?%����M�%�T�v1sA��!�������O����������>�fТy��'xw%@�M�_����)��q8Ւw��e���E�z���1�F��L��u�W��vT�E˘���BI��g/��>h,�B,�0��m�d�$t)���Qȅ3���Gg�Z_JmC1�9����8�~�RqE�x~��*-6����C3�����RvJ�V���堅����p�a	�9' ���=*�U��sP���ćp�cH`d,�����ȿ78b	�eY�ub����/	B6�X��0�.|���>����M����r�zU,1w�5z�@���g�Np���V�X2��%�:Sg�͊�'��K����o{J�yD4z�좇��$���*��n���'��g�@
���-�'=���J� ���`P���fRv�9(|��g4�с��!7&��s�%2]��`�%,0��H���ēG!��sZ<] �X[����fB���f�8����ҡ傀�Z��)A����Y�O�ϻ���s��>X�gA� Bʓ9S�I2df��8��!�o��
0I��+ڇ�{��.`D䂷�"q4�-�8����kx/�������U�٫��=�M����I)�3���D)PF�Ս�2��H�y^X0��c�p��a�5�;?�&]Ë(��:�@�VDήJ�`���%��SY�	^"�n�}�HoyZƽ����sHP�o�ћ�(A��69�8�W�,S�bqi��� �a����;��@*eH��ԫ����m�����o�O����2i��l�ܱw�I���/�7�H��ˇ���:o��b��(G�lV	��y`�R�M����lq:K���~p�{�/�9,�}��l)����}"�������ѝZ��r(~���;��ha�w�o(���Re����n֗���w4Rt�Yg�{���OV�g�ָ[$����8A��-F%�:��;g77+8��^���irRS9�S��P(�똸4��F@��h��������ͮԮ�rK�9�~�]�M��5�@%��|��IHg���"o�X!��ڥ�s3: 
gc�G������:�&~�S����0� m*�%t��; ��.���t�cg�a�Oo��x���s�;��y�c�K �[4��������� ��%`� �KO����f	���}Z*�^��U-k�N8����)��P{��qvm>^#�o�������e���" �.�O��߿a��[�r�sQ	@����/կp�~��N����/��[r&�Q���Pqp>\M�,u�ڢ}��]�{�N����#��玝�
!�܎�m����N�_�� ̊xNV=:�X*�0�M3LȐ���]��6ʢc������)3]��#�����>u;�D%2VBc���Yz!a�rv�V)]��D�чTMa�z(��,Y��E񙓤H:�E���繡�F8	��B{_w��4���G�E�Ѷ�,��#P��>�z�v����"�Ш����1p�Pك3����x�sK�kW�Ja�[��L���}�%�3��Qdi|�%���Eu�_�KR������t�cz;*x��_	u�K�9'ة>��x>���m�n���+t���ޅ����	�\�l^y2<��V&I�s6w���n(���߿ӖiXČ�WX�U���e�ve�Z�z^3�	�_��%̈��+��S1S�I�d��,8��F��4ۏ� � k��|]����:	�)���#h/�]y؈�^&�����oR���Ĕ;k�)W�C��UG���Kw�5�'#�kKG��R8��X@#�F �@�d(C��t�	q4Y�ҧ%+����]��)�^]�1���½L-��Uղۚ��TQ�v�CQw|9��%��NO�u��?�u�q}��@�T���>a�
̨���yOI̳隫<�E�z.��>��h��W��,���J�2��qN�N��Yo�o���{��L��r��C��V�[H��x�X�_��v4��7)?Н�u����h	�q'$�j_���a�	�H� �P��=��
�ѳ������� �n�}��EF�d�p���΄�<��_i5���w�<ل4�z�7�H:�wg�ID��� ��%>Y+Ŏ�O0���{#|�N������g���궀�/Ә��v�X��:��g��o�j��8���Ҭ`�o�~>iݨ��4&���^cv��0��!�`(p�	X����-�- �
�M�}:Z��q��	3�mF�v�OK8�i�tKA�9���>$�v�|8J�qR�D��
'<�+QC�C��* �bnbF�c�`�LEB�7�S(�V���OHG��8P��.{U+�_���n7�-Z��.W���W{�2��9�*��[��'�T�^��|k�����s��|d銟&�2�-��a	�T_��٢w��(T�J�霽�V7��G�%'֚�Sg�(6����QX�6�hf��d�Y#���SG�_��T� RـO+?���(_��\&�<y���?2Y��D"_�է]��� �.eG��)�{ �+J�6�:Cu>ە���k�Gc�yZƺ���Ք���G��	���n.��4�p�u��=���0�'("]Ŵ�y�F�<����o��@�,�.hk~|�T��k8$����' .\<_��%�N孨�8�>k�ᆯj���àV���xF��
l\@����hp�Ltz�_A���:;8���7�OS�@-���J�@%��.cV��a1�W3^����\ yK�M9M��"�Z�?Q�rC:�
 �Ja��AJA>R��������.Ҩy�#|�s��Ӻ�z�~V�C��<'̽�P !�Q�����&�����?�%���	�	{�A��`�ǨZ������H ����H�&�*���N'��U��4M1#&`��y��g~�Ώf�g�G��=��W�צ�No]�o��l�|ɧ*�����<9��q��-��h�ΗFMK|�^9���fF_���m�uJo�v=���kv*c����2�rC:����23f�����>����rD�q��h��D��*˼c" �e!�.��pq���h��������o�;�$"�dk�������vo�LG�����KZ�'��mt������l��V�N���\8�e�ܜ� �>2���[G���YbT�⚿����kU������N����P1���I�Lú!���+y?��Q`[eXt�+����*z�E�$�N�> 4�|�u��48Trρ��q,s���� �=Hj\7�]�_t}]u4�����s�':�]�I�4p�����c�	e��|���gu���э�F2���v�A�nN���H�,8�\].V��?��t��E;B����4�ɋ�P��Tu����P����~�è8�ת_�Cމ��KE8N��޲AG'(��+�A�}�7� Z��'���ѸMQXxl=HD����hKT���J�M�w�]����\K�;Ӕ��vaCOb�������p�g�fjE�>m���|�ةG$�=�M�Ëm���f��N"�ܸ =c���܋eҠD$���6δom�C��$h����{Y�5C��,�Z�����I�S��Xaۈ�N��5X>��U}�TX�f�i��D��cH��O��W-#貐���Q#$2���4�-���D�!�؟\�Ys��vL?
En��a�8jA�%ML-�A]CwG=Z�G�q�Y�k�K��"�US�3�	�CE���A�M��<c�f;(IM O͓/@���+�J�#f�m:�,k*t2[�]���C��SH��i�����6�pɊOx�����*�����o����3����	a2l��Lf3CR�1�[T�ܬ���U��cE�c�Z�^�Y#Q���(���1�Yqm
��܇ۿ���3y],_k/����"�����\�3�-��h��2Ԗ�!_�~D{D��M��h�({7�r����#�PSF���ݮ~&A@��7��0	m㾁�� �l"�}�w�U|�ߓ6�tO';�k,����6��?�+[�6d�S��rC�T�(v� û�w_���O���aY�!�EL�u��~�pl�9�!/˶®��=s������^����}�.�>%)F�����ld�nF>Ma"4��1D�s�1x��*��� �oH�IԸM�e=pqy{�jI`�#��Y���Yֈ19g���B�m�صY�#�%����Ŋ)��|��{J4���#FʎS�1m._�Fd�(Xx.
x��
!�c�"�:��|��3�ͳ�&�/o�|�^�`�+��T����oH���$��e�_:�|�+%�bY)��»����E��"{��igP�(�0t�g�j�o\���1��&�K���:����"�S]PђM�_�0`���?�&�����r\f�����o��ED;_٬N�ۣ�?��-Z��w*� 2q��ꩂ+��ȉļ�r�0B�a��1k�b�U�]Lq0��v�	�t�z!g�ȁ���댵�,KZ~�6��K٥�II���A�kF?}�]U��Os?hޣ�TpeA���a����r��\�K���#��V��;��ܤ
�gz���96��=YW��kǓ� Y����� 2�e2��D8}~K�dO�1�b���1������:qP>TF�%�f.�L�����T\�oG�|ᅻ� Lqieڂ��HTr��ĩR��y{����S�{��dǣ�s��i��U�*a>v͒5�\��	ý�-7/�JH��O&���w�Wa�h�f/����o;S{��\�g��O TKgq1�(3��,2��Pm�.�$���.8L����G�V5�Y@s�0U�-v��;�7-��BnX��W��FJ�2��KXES7�Z�o��M.2��u�� ~�C���TUr��]1*�!&����計�_P��[��4��]���/���=.��"J���=��n&��Y�DP�щ�z����	-��}�@�Pusƅ
�a$�� 揣vq)ԓ�!R�R�{fW>\Q��؄nq�m7��[�:-]eO�k+n? �&n|���c^��2�\���ҡp��#M�H�@~�U�iy��0y�c)�NA*���
����������U�l��~3���T�Q3���ѕ�1�۽`|�(����}~��`�)����"&e�;H/_Н��(���_��1��@���7&����[��4��8_�]+kI��ѭ��}%�Q�l������ʘ��q��Pķ�6������l�ҍy��I�2�
��� ���F����5dR��l;Zo`�)��2ʙ�KB���qY�L�ȏz�G��1V�s�e��0;�R����B	d��D�b�RY��Zړ�?g#l�SI�|Z0��v��n��!)����f�����8��A~N�ܞ�z��Fd�4)�����7(K-����h� P����z����ՙ�X]�Wpn\Ӗ$?P�c ��:�6��).Bi���(wEG��\�O�Xk���~�������N;6X��=��m>s����戴���Fl�$vC)�ԆP��>t���=�Ȥ�&G{ }�H4��c��t�BΕJ�`�A�54 ��F�E���%�b�h����:C��\��<�+����R�~.��@Q�c*M�_)�6y\�r�`�P�E �N�5?�OUgn����Q��>�%�q�c�5�P�˳�bV���,`��NI�BK0� �opp�ѝ�/�~;`0;F6��1X�r�h�9��=U^ I��~��z!��~����ɀcQ�~M���w���q�L��j�\�S�m����H��+��Cg�GK��M_Fw�_qx��cI����AI-)!J�E��5p"�w�2�'q�C7��=>�1����r��J�/�&6zU]����a������}}/�i�=����Ey�'���V����1w�={�,�N�i�4H�Rp�` Gݙ��81�|h���p�g����Aӱm|�9�KT&�1�Z�2蕞�H����(F
��NWڐ�M�fbQ	���1R��E3$=I9��<�mf.�����}���u(�}H1�7���V�O�z�Pt�F�$�;���83My��mK��,��ujCO6�{C���&z�?��;���9��}*8c�Ձ�>ӸJ��1���"�� ��W%�e#_V4�ed�Ŕ��~�T��	0r����N38������s����7W��B�m�,�Eg�'[Lnr�h����@��Bi��-�ڼ"��m�ڤ��*��ҷY�}-�%D!��t����֌�d��� ���#�(�|x���N83GNs�\˙�!�!��v/6�?^���J�;i�|� 	�?	�۲���3�{K�	T-DV+Rom�9��V+�H1޵�i��mtE��6�ޗ��
�'>��DE��s�d4�����؆�Y@�%�3�kPݝ�|�+:� $���N���gY�:���c���I��᛹s)�&y��@��D������z�:�>��.	�"Z-P#�UJ���� ��b|�۪���ۆ�x���m$��d���_�����+BY��LX�<�ɯ�8>'�#�>����0���G��
��ۣe� ��}���^7��{�g�����g���f,:|��L)9�)r�˓?�<l��{F����8M��ξ�_�`.;��n�^��}�_�x~a1��~+2�Lp|O���������MP��G����ș��ZW���� 'T�iN1聰�����L����ñ�B����S���.�t�93ln#��a�7���s�F��2d�'����ﳡTR����A�},��,X²�C ������a�
�l�YcI{�����W�>�#�HP��({�S�6�}����l̓dI�Zt�(^�qoF������&zm��Y7<Wm�B�sf���J��ӫ���ȭ�֥��_�+<��b���Blv��j �/���`���.��Nx�>r8T]�^�[�F.Ʌ��)h
F��,��nĥX�dD���|ڂ>��ڎ����hq$�=�o߯�n�np+A=˖��ƩL��c'!%��%o�,��C��q�
MV٫�Ӝ��-������#i(z��/,�ɐU�~&Ol��y'�t�Vp]�m�fn"u��Ͳ��YPqP�ޤI�ąj3{�&�� 7}�p�x�7�Lp��"`kO�$�!vt �Ĥ�T�^�1��^"��=Jw��>��Q��l,wϙ�<J!����AO3��~$�i����j�w\��H$C�5�S����܋Tˠ'�4��"�/���� 	���<�~�2+g�D�CpȻ˘K�D�f�)%�������	O��/�ӏ��V�9���q��n�����4�Z�w��,���+`��z}9Z��� �s���N����ǁ�Y�J#"=�-H.ߠw	�*�(XIvҾ��G��1���N>�G�V�A[�S~[��t`k��H��V����jw5�|�4e<������;;ͪ�h�H������F`_�&}�#�ܝ~���*~�z�x�+ԍ�H$�)
,�vf�fx�ִ�V�����#kL�2��Q��FTeW���(x�d��-�$·�c\&[1T���[:���Bv�D��)W�P��U�.���;)��ލ��`�
�ԗ��%����C�r�Hn���۶n�a�״#�`U�����t�Ş=�4Ɠ"Lď48d()k(�C;!��3���*��Da����FEZ���EP䯱�Ft�+�S#6�q�Ɠ����5��\_���8�uO� y
6:u�<wq�So6�Q�	v��l�آ��Ȩ��:N9��J�Dp��t�Q��:�ԅg��j�I��cpM�X�vW3�k�)ɞ�ƶU�s���H���>1}B�s�KK�m��Ӱ8D̏��]���(v2y#�É��w��#q����}���˧WL�(=CU��"�i~7���.�4��A��Z��#<
�d���=D�s6��V(��I�`q<��<���o�='���-�\vkI�l��봪�$.��?�`>qlB��hG.�&sR4h, ��=m"��Y"�\ÎJ��q�Ѩ�P��he�29�n�cJ%�.ZުME�\��:*�O��s��-���U�2�fa4X˲a�F�1]SK�B�-	bz��Du�/��jT�!;�����I�β�O��Q\��ANu0�ǄEl�	�҃A�V�د���b�����7-��ؗ{W�O�f�Ƨu��o��xt߸�Yv�)���>w��t-^��0&�'ȿ7����� J�F^���lۃ�P��_.�PF�V6U���+	�Յ�05O1h�Є��eh,�oq��byvL��H���g��6�$#	��/�ĝ�萹p} ��j���jy�
�&��Dq�]����S$ٞ�b�"�䂐����ʏ��j^�9/6�rq��(ߦ\��(9�fXb[��O�%��CD��7����^.\Y��o��cLF	:�"��P 7����%�R2���?�@+�y�lxv� ��0����}�$Aѿz%\P$	��D�&�4[�S�A�2x��nYW|��N�<	�gG%���y�����AGLW�A����z�d�Ś�C櫿�n��-hl�k�0S}v�=��D[ib{�]Q�=���)��;*�Y)��L�T�w�F7�)BM\�Y�Hv\�U����A�Q�c0N�"������!��#h�:�Q������4���Q��j�xSiUS�jj�z4
��������ʹE�n��:���q�c�c����+_����[f>"g��}���� ��7�*�]�^��R�֜+�iu ���Z��8 �L�NC^����0�?B[���A�Pk��|4տ9o�!�Y�d���h��l��Vp�� �yv��j\������<k���Qdy��3����=���G��(�Lu��Y��,� �#K����Ω�F�ӫ�Z\��iئ�G.��o1_ˢ�1���R#^t>��0>�̓�4��ct���2���Ȁ ����7�$dIˀC��!�**��B���c/aa�8.��1�¤L�_^���Ma�t;��:���%�b����.�8
7z�$�|E98�u4hэ��ӎ�l��݄Ƿ�D�ޓ��oz�(��4V���S�=$>e��=���z��� ���2���;���\w�E
�Ҵ����7�&`��r���*�M��6��D�K����]��|60�ķԿE��YM:<���m-C0��x���3��
�!�m���˩�����]�����t����MQ��9� ��qȔ�a�W׬Ra�^ԖNhAF�{6cȀ�Ń6��~����>>�;�h,	�_�:��˶��"��Ϋ�eTN�.P���͖EyU�]���;Q<#�/��|�夠�wno��Ŋ�"��x�� �!l�f���B:c~;Y������}��A�i��'�&@ҋP��A�	Gi�i�����8r��i�B縶9B������P��$i[����ꊨuS�o C�/�c��kuM=�/'��%�gAÆ{�+���`�>j����=����� n��a�ϼ�#�؜x<#X��e�vQ,V�G�1�G������r���/O����!��2Z�j J��k&g�]��=���L��∳��D�?ޮ�큄,,��Z[T���ni�(��p2��8�ew2�+���ʓ�E#X=��4�uFo��1qk�ˠ ��oe��AjW:��k��* ||Y_I_���?B;���/�0�}!�H�T/P�q�;]�M���\�֜,���:��h�Z��c�6���
vbd�<�ءHJ:��"T�<�8jc���������_Fĵ'7$΋ӟ#pD� ��[�䐦]��ȗڳ���X��Z��p�9�B��P _T�1���s2q�޴���y@L�T��Z�4��q�l�4.%�©\$���&�4[MQ�?��u~x�̀�=?\l�M��6��@[LL��bt�����C�|�G�s�z�v�޾�k\jsP�X俪< �`��F��u�>��<���&�:���q���R����QD�n�\��"��I>gU���N�8G�x}���ރ�ti�p�>e��HY��J�1���){i�.7Ϭ���n��ڹҏVOIBr` Tk{��Z�
o�g">�vP6��u�������D�����s���;D@�������a}z�X����F>�ѓ7(����Sq	�X�֡�v�a�(Pc�Rq?�Mw�W"����w�Ҿ�y�����P6뢯π[��'�G���w��
A(|���� @�����ԕ�,$ml�)Z�u�H���j��M/�v�?̝%�U�0��<N�f����4�Q߶qoobֿ�Z��P���`(}j�G4nD0�h&�'�-�S
�bI)u�^U-��<X¸�	�-�Қ; �A`�<��c#dޣ_9�#1�:d0D���~�/;�R�C�r�Q�?X4��zB�����m�!=Հr�2�h��Nrg׃��A�T{�(����Z+g�r��T�J�$�����#�5�$�JE��k�r��knV�D��}Z!�>�V��V,Jѓ������jb�
3q��t�;a�nbB�%N C�4��/ ��P�t�[]n�@�	��xȡq�9Fʪ}V>@�]�_���'�W� �r��xc<}�V\�Y� F���OLkF��{1B�?[m�Q��	��X�
��x4�S(`��:+sAZѣ����������篂�� �=r��-�OX5k�{D G�8}g�� �Aw�ɽ���/� ջ�Nl1[��+8�,tF�xOd=�u��$/T�Q�$N7���}V u���o	6��r�� �:F���(9�&��5��=ߕ����}��:w�)�1�O�/��}�������Qs�>�&1(�|B�6���z#�Z�W�clvV�x�j0���{��U�r���ڡ��,!��<�q�{�U�xff �����`��
Sϼ� :7�M5�A&��B���\����Ì��ՏVO�'��0���w�l��Q�KdH[�Ez����=-����f2��=��S���%k숛�E�d�^���e]��UĞ��4<�c¼ޣ�����Y캤]��5�ha�E(����ԓ�N�	��I�_���Bw���O�I�$�\=�5�;a��רR��n+F���3�T&V�	��0=��W��'�|lNzQf=J����ĵ����:���v,8S�?���>9^mIW�f�̛�9��y����e%I�//�+\+h��{�����K���=@��,,R���h%��^���؟����J��Wr��d�����?<�	�8���l�� !_���g��^S�J˚�:�m���-h'�?[d�<E�+U�{a��ˋ����}z���#�==����#k�O���`%��HSu�S_2�p]�0U��ᏗSS�v�[{�*e�8��GH��*��x�r^���yN��@+!e���m|��rYe �Q?J�襀���$��39��	��`��d�Y������3�`�%�L�
�~]�e����Jز{�5k�8h�c9���oo֑,1��x��Q��
"9�l�,�`���-���l`(��l� Q������b>�_z�p �C��UUbx� +*���@�ٟ�;��g����
)�ؑ��D����+��p`���T�0.���X�?�oX[��aˢ7Q\��Q��&CA6���,��F�Y�^����1bVP���h
�����z,�_���h�=��j��~!���g:��Z�.]<���:t�>Jħ����]��`�e��H�W3���nP�m:\0+Κy<|��Xٟ���w�[��/%���k�tL!�����*<.ˁ�Ix�zx���w��oh��O�	�kE�]T;&��^�������*Ҋ!�㫘�j0��P�J@����Ɩ2�2��C�sC����d���'#Ƅ�C�<W9K�n״�){T�6�	�~�<B0��,O���sp��Ǥ��O�ܛ'�������Cy??Bj�_�甆�f.���27V�	��e����,��O�ͬ%�5����C�(��#�;ā.ۻ7:uLA�M��i��χ�'nh�Y��5�u����Y��G7�:�ė��=��/7��@�^�N�R���cv{�H���$8�Tuq���?N�Uw£�c���e�!`�SP���*`
��t��>��H�E�x%��\O�gf��5�/��awt)�fc��n�=�(&BÎ�Gƾ/���hۻ.Xp��Ԥ^�i����d��K3Y�X<	���DhɁ��[<LQ����-����E3*�
G�s�鉿Ҳ�����:PwF�Ś'���ю��rl�x�2�k�;G ��y��~.$��sk�5�GN��F��%�v����/�`������Z���	�$=�g�a �_��Ż�4����l��yeB��G��S�A�����{S�6�C�[�FJs��NA�[d�ͭ(���1Ɓ"�^mߑ�}=j���kޜ�8ہ�짛�B��Y��Ҷ����|$:/G�a>�+�`b���6��cS�:L|��@����J�+Y�z��l�����SK�f/��/5��B�3I�!4e������&p;��g[mGZ����c�7Ezk����3��)�:�jcN��׿J�o�r{`\S�Jt���V����V#�jc-���HƵ���,��5�O{��٦��Y=�.LN{��f�+]d�<��x�ڤ�C4Tbר�?
	�����n�@�0K��0�yմ��!y�n
�u�ϗa�%}�F��f���)�H�t��0�1�d�T�[��U�V��N�_N���df�ui���U�QWy�(����9
I��V䫫�LuR�$f�~y
Y�kַ�z�W���a�Ԃ�1���5ƛ�֡ɦ˳7�q��:$�#׋7����X_�T��]/bN��3f�r��i1巏#ى�_%�1��]��C)d�tۇ�<ꁔ��Œ��k�8Z��r\�^k%Q����.�-7�B��.���K���-:�0�ˁ��ث?xHG�DЩ]0�90������^�4�2#��1k*��]w<�X8�S��ɺ6�辩Md]���<��9°/��(W��h-��Z� Ly�� g=��O��Jh;/Rl�D�U]�8�����G8 j�#�Ω��3.~qf�@�츕�S���-��[u̡8��$)�&�o#?X�l��;N�EXG>8m3I`�	[z���x���+Y�4?t�����|Zz����@�����E�u��l���C�Q�n�^��`���̓�Y��&��W@Bf�n��J���*�$���iV�Z������4�B�zV�޿i�!vlu�Z�AM{b�P�0��(b���q��^��8[G<�Z�v�S0��NC����*U�L�v�ab�@��$ѿ�2$ u'�*�X��(�2Mh�tdq�^��3+0��~�-x��W��Q��A$��d�Wz�^׎KHf�!�]��/7�Kf#'���]�q*�^mWP�VR����I#�0hk��x��H�ݡ��l�(%+�P��v~!٥��_q�\ɺ܃�k��&g�ͨD��f���\ӃgD���l\$�S��Mf8�`���l�@	>�݈�4ۼ�u�c�R<���_��0X����V�����^񿟷��_����6�y~S}_cBV�Z�lMȟ�4��7���zrtcЙԥ-)�I�vTb�Q>?(K�����o��&��=�w&���[����B��رG�7���7<U���s���Lt��S����N�l��u��>�R �y5�t���rB�n�)�a��2o�}]�/�S1���-8��jX�zp�����Q)�W:~��8� �`��U(�$��CX,ǂL)����D��e�����d٫Y���R�m�^�]��d:�zz����VF�q{�-���zot���������)$ge�*:���!��#x�	��fs�XO7K�� �+���/[�ZҼ�$Oѷ�]��^���Fwnմi�l�<���S�ب�GhP:��ds���3�05�*n]{ ���?cט�B���i�4P�ȴ�1��N��h��V2r�|�Z]��bg��Դ��0d�;i#���Xz��c�ޑ���|�[��^5�^�ɕ��ݧ�6�Z��e-�
��Q�Y7^�Jxl��ZZ��_)
q�'&����b8�h���F��!,U盛q����]m���3Άd�#(�n�9��%�Up�ކy����,�^�nА�v��!e	����Ki��<�$j�e�9S͏BmF�;�c�.r^gߕ�b�9�=^�Z�bV/��r<���u6�|����&A�� ��P�0�̻��=b�:~�(����4)QڰK��g�փ�c
���'�	:� #u!��nDz�5EE`�Ӻ�Y�aX�/�b�Ɠ�dz���pc�rI�=N���B^u�^y_~9] �`�4Ѳt�i�����+̣f��Nj�$� ����5�")�&��#u�u������8uhI	��k�/����,����u��H_ġ>#4�g��F$�K7(�q��y�TV��I�4e�ٙ�:M��a�9׵�%��n�,*�~����}��e�h%sA��>����[�E���p^E��|�,/ۺ �.q/��Q1�����YL6X�,[��d�i,:U�K�M&�4}��xT��*���������[�T밝�"��,��Y��>
aV�h��nsGX�'�d��~䊨F[��+�P��aM�\�|ˬzqm�cn� ��y����B��N	���e�ݤ���APA��;7�b��ʶ���뇍�Y���S"�h�RC<U�üX�#H�6el`\�{7B��盆��?oLow(巬��资z/A��j���@%���[@��ݫ3��dC�\��)7��ƾ�n/�X�U�0�#�_-���0	A^B���`�?�4��H�0���������Xmo�X:ɆI�?����.[	+�e�?�q�$[SJ*^+���ҘMm�)�����<���ڇ��L���0}VdB��8�鸩ZXnW]'�Mn����ő�n�R? R�@����i����Q;mڵ�Lɤ#p��E\��NMS��/J�����T3����<����TfǑ��Ȧ-�z6���=B�뇾�:�������`�&����.p輨��+՚E���w��T.#��`oҺT�I�>ci���?��c�+B���,b���3�];G;�n"^b0S.�p
�ί����>cӣ�E�c���4�Z� �|�M�Z����[D�2�����Bl�Z��Y��BA�?J{�v�	��P�6��qd����*\d��������A��fj���(6kݨG�����B�}��و9o�h*g$6�V���hne�[�b�6[n�l��"p����*o��r0�v��^�N1���7��1q��YL�����W��.=+��ȸ[|9V�1���V��4o�`L�VW��n.��v��Q�iO�_�ͫ��	G{Ɂ�
����+�ǭnV��{��Q[�خ��ټY:�|��?��0���H�Db5��nD��ߖ�Z6����_LӡP�X��歪\V�]?���Ȫ -46�0�tJH/�L�`��Y�2'��UF��{�x��r��U�e�����ug(����i��ʷG�]�ɍ�.}s�a��LL���`R���p�sR���m+澸8qV��~,���s�������p)e��� �{���}/��g�G����y���{hh�"o��ju�||x��#�b��C���{C�D�ʈ TN���Bo 1���=����M+�oK���/��=�7w<V���d�/�	�
�IR�A<�H��N�1C��7�0'�{*��zKi\8R�;K��yW�@��oy8�|l_7Dy�뉙�'�j3�gڝ��B�J}��������\�H~�v�NOO(�y���퓞���QМ{���PI�o;	7�y�:�#��	-�)$C�JJ	$�<#��Y�R�T��ɺICݟk�-8�_s��f�uJ���5� Yǥ��k��s6\�=������	�7�	
���-N"�3h�Y"�/��F�Y68l�����k�}��G�fi_��Y��~'�mVUU�N�\��5O(�?�&���-c�!R$���ۻS���x�5��J�1�Պ��sW�	���f���q�2�I�4���A�=�5\�b�
/��:FJ�#d��]���L	z�2۬LQ���=�1�[u�30�`���1S�idL(�J7�6ꃁ��7�ԛ��~��􅎭�Eoa�J'�EZ	�m`�)e��jߒ����3�������p�T�컬�%�9���Puy0�@'��9Y͆��cn[Új5�Zj~@O��Ȅ|�i����H5��W�(��XT�Z^����)���2a���Ha�9�L徏���I��%|�fu׺1W����WX����ͬs�nU��*S4�s�g[L)�`L�IM��Niy���*Ӱ�?p�\|�����})���C�������r��0ުla+.��M>V�.@���Sb���M��@v��t���������Ǌ��~{[�"�e��E�� ]�����	l#eT\�f[�d]z]]F&�K��Q4ǐf6P��G��a���HW��U��W(Kֈ�'���>j��SՅ)w��SՎm���
}��̇i���Mï$�0�j,�g=����FGS��:HEo��9�r�tH��Ƹ.\/{0�w�g��u&�c��KZ y�|�H=��Ke8{�"o��s([��('�����;Y��b�����zm��2`��O#j�Ш��{��J�q!ZaJ����P���ȧ�;��J�n��G�x�����϶� X��ճE.�$����H�pa� [YQ�����2��TL������lGaaS:������\�c HP�}�Ӭ!��x�rh�֚�x�6u<m�H�p�q�'��YA:p^1���d�L�¦dl�9j�9�8v��𡧬��y���( %�}���s���[ٰ��	+�����)�#��/Nh�Q�=����Bs��8>=�;�u5�<�mdPe:��镶L-�[4=�$��
��9㗑3o4�����h�3�fs�b*K���	�`�O�X�:�%z�U�lTMޟfd���e]�7P�FE�������d�f-ii�tSE&���+����	ƑU��T���#������e����=��U�@�h@�KD��I�#�$��aN�?��3ۂ��������S��R%��
�g�s�}#^�p�A?�w�WP�q4�o�tw�#p�~o`�;��:���(�4�r�GscU��R3�q�y����/7�k�b('���2��4%#?"�~knv��>�+`oB�ۦ����ch�U���%(p0�, 5G��hz�	?��G�3�N��m��Ͻu�=��"'�(X,JY��?������]E��Gtn�Y�H>�����_�_����&�Zn��_�B����/&��ɺ"p����,��<�#qa��X����{
JEZ�4��s|Ԥ�t��V��61�P|�R=�ֳ�Qe��>��m?�ɛ�b4"�U�.LOE"���:>魙
Q����=���=��l��t�t��A�PU3"t�k�t�vbv)wڅV�O��ED���{2�^.i�|�O&6;��^�w䊦s�(c���������{��P5�)�:�D��k�-E�X�0���쩎KJ���M��6��zլ��~<d`��=�-��� �ъ>N��ˈNaq�|Q�e�z	�s򖴃mS},��`ś�����[\ݚ
���r�j:t�仇8���"4E���,T7O��4��������>�&�:�_��;�I_��'X>d�-�-|��l����,U�:za�����N�m�c�7��*ࠂ><�e%��W�ѭ� Y1Q���\3Q���U3�{ʡk���k-R+8�ٶ�:[*z�c]��������x(��; ^Ĥ��ȁ(�|��38'�\���}׊�P�m��\i�1�FJK��dZ<�h�WJ��T�``�-1�h*��7I$#�\Ν:5�"߭��;�}���+;�͊����n~x�I�_�]�~��?�+$ ؖi���	w�n��Ύ��Պ����C#�!k|�бm�Qs��(	��l @ũlo�̔��<s4�Xy��뙒��:iuF������1�+j�[��~'�[zS[.IT�X$��S�]��E��;h<xdڄ<S6��x;��՟Ƀ�jר�O���Q�(����`d���7�R;�9{̆�FvK�fF}"-b8&1�v�q���s��7�Sj�W���b���Y�O��g*sp!����c�訣���������[<����r�����@�	�w���H����߃n�ضe��݅M����Q�`+\|��"��	v3#���b���ڲ�^��-e߮�s��j����^@�y��o�D���+�@F"�z��j{��V�Z��.,.��.��q����X���"���U�XE!�9wx�Ɠ��@2@7�0/��P�S����^��?���(ĥW��BA_�~��:"�*ebWɀu�C%�͝�i̒�ji>TA|��x����5�)[&�P+������Lt�ݚ}#����!��H�{��´0���Wθ��X��|��Ա�֙���ͅ˙t"^��Sd�ƇkK�q��n��k�?g������b?Ǧ�rK�+j��!WW�$ L��<E��.�9`3@u�8b�b���l���d�z�}Hn�"2�U͇
��d��2��&�
�+�b:�lA���EP&�A.�Xs�	�&Pl��8p�|(�$_X^Ƽ#e�"��5�#��F�m@)���'����ʩ�*ݛ�h.y�~��3Y�<��Xm�H B� a�d�$p�P?��+��x���}57�m���.��f�Fj�n�W�]8{hR��h�D�:�vW�]4XF��+_d�v�=�~ �R&~K[͌�_D)�}a��x�����^�t�9�s�V���iګ�>���
�VUaY���w����:��ͽ����]�)7���)׎dT��q�c�_�@�a���"�3R:-h�O�z@�6�B��q�OG��Glz=�4����~�6	�%#�o	8��{�E���ø�;/^�N���,��>�A�ICay(��d-KI��+��fd@��j���!(�Za>��hO�l5�� �Zq�܏���J�5��e�x~�v�~xa>��q�S	}����Ӵv��~�>�����o���������B�'� d`��F�0�;|��F8��Ȗ�Wh�9�0G�Ė�˩.D������!�4�l���n_��S�{?3���+>U0��9��\�G����(	�`0�OX��!''�(�xtY�M8K��ڴ�J;�'fg����c����d.� W�)���ˋ�L�2��A"�UD���	S8��mt��I��r��f��<�m��ǳlJ���R�^�)��\�}~]�p+\eؙ
������ւ�F[�Q�8XJ�R�yV�c�08Oĉ�"E��@R}��?�����Y��f�0�}Y�:��ZsL�C6jd���)����^=�tX>�mE����P.su+�)�9�	�\��.@+��/�D'V�b8F3�dw�~�>b�y�1��
M= �b;1��,�!"��b�6a�ZiW�E��	j܁��Z Z�0�e�#n���W
N*))�g��t~��
�Z2=z�SBe�E�$Bn�r��NY`e��j���;.̙R��yǛ#Ĥ�F/x�$O�w�ۑ�;e�:	��p(MYvy�"��
�u�5ھ�M��~#7�:���Γ�%��A���-��M��.#s��r:�{�
�3oG#���[W�t�q�kղ	�ڡGe��\����II�O�Nf ��yA�8���i=�56ޖ~�}(L��!�Q���Wo����N��+�_0���{��m0˭vIb��@T��E�����:'���y��D�#�h���1u��C�F�$Q�m��� #�_B6��lr_Yc9��G�'*�~������A��Lʊ���[r5�s���D���v��x�6��!�O� �!P��$-�������u�> �$��/S�b{��V	^̴�X6�F�[9��B;(��'t� ;AoO�>M��	〒p�0�'�1��c�T
s�7��c8�^���:h��P*S�P��@�@�0�NL̋$!��fVrw�w�<נ/gWk�+l��J�Qk�������ϓ�Z�g�&h����1K�/(���)��恠���?XQ���I,���ҫ�� �W�@���#���Q�{������������!6�p�\@ۂt����Z��T7Uj}�h��"�
B���Spm��1�.b�rץ5Y��+�S>�s��L�	��WCFjS��*J��jCX��$�m�ru唪Ԅ�a��ƆC��4r��	[H@����+w����;�<=�*�aB��ƯeW���o���Z�Q���(��46���0�C:����I}�Z������/�^z�܈n2�����# J���u�ɜ+���dn��Z��c��QMD}x"{7�[b� ��&D���~�C(�)oN��6��,i�,3��J���ȍ��e^w�ޮ7�N��	�ƈ%��C���csf���h�9�1�lV/��h��2zM�����s�I�����|�nd�Yz����u�o6:��O��M(}1q�j���Q��dQmj6��G�}K5�[(/����1����1��*چ�Q��gb����d{�5
d�P�,K�RT�&w�����4v.K�i0������v8_����6�e��hJf"c���.A1*C��|�'���}��0[ɵZP��� ��e�ѳ_Z+��!8To �M����K[�*�)�vd{��>A��?����6�s�f�|�⸵������yy��y���N��۹S��Z1?"A/���x����\I~@b���)��F�Ģ����A�)zw��������Q������d�b����U�;���4��٢��d�� +y|��j5<��kO��=�?���,���}岵����EW�^~-���I�l����Y������)/�J�iet��v[m�@_k����t�s'9�x�~�C���
�#vn��.�U�Ce� ՏF˾� �+�9Pj�����3B���^����Rgx�A��>����kP,b^e��Y5�	�/q�o�(Eӗ�=�9�`�����t[�K�Ob-�\�:�i��]�p�k��M2�mg&e~�o�:iM�*��R#^_y#/`�j���F�t�/5�K�i��b�땴.�H��1�ڷu!����}#V,�"�n��nv8�1|�5A�Γ���'+���^��U^��d;�����rv�����i��s�ek�/T��V�^G$�%��c.�$:1I��X~��~�-���Q���1�!b�E[�A<ܨ���k�a��>\���8�p���ۄ4kv=���0�����`݋�[��������×`~[h�y]�M�3�y�C��##��+"��u$�~.X�MY����[�F�q��{�q�j��_� ?� �_�P*�n����~�fY���e�p!�DΠN�آ���W�#-�`<c�b�~�8��0��w�@��l@y"�WQBW�B�i_d�#���]�4K��~_���l�}#�1:����T	 �x*@��m��=�J������[�5���"W��m��h���}x�U�ae��Bb/D��]+���YmY/#A�%m�8�
�&��<5_��ː`� c���9�Y�R��ձ�E����ph��l\�s�!],�6�9��a#��+�N^ɵfAJ�麚�p�⹥��.�J�q@i���^]!Z�r���k���D}�H��N�����h��2:�CP��D��&��vu$^��S���`���\!��fͳo'E옗���R�7Ю97�3�+�.!�g������q�$�I���ؐNG`hռ�������z{����M����������`��@v�"o�`ws�Kg7`z��P��]�By�߾�"4�ꔬ�P���v��O�0ҜN� �%�K������G`�z�zGh�l4�>��֣��p��� ��NNl��R��TnX��=?^���],��V�4N�/�h���F�jy�,�U��"���� ~^wj=��S�'_��u��(�ZP�fO/.�;ژI��*�Na=�����C���}�W ���-�eg!�ܡ�>\%�t�@j~n�B����M0�jH���T��T6Oz&1B�<��wM�N��B�D��z��״@:ks0@L���i�e�-Rq�͐ Ÿ������CMW���v��c*D˱��DV���6����L]N�]����~���U���9tþ3�����3��"����,�@�x�,��cH�kbrT��Y��x��K����G���~�j��\E�ìِ0=����$�h�l�d���R���?�y�����ϜCxK�e~��;�~����sJ����.��L}�vO��i��*}0�QI�8򜗉���F��e���̷η�7�Hy��E(]T�gF#�K�NPԩ�H��r@�O�`�؞ ?�cs����8�["k.���*�<g�+��%&�#|eM�Id���$�@5��:�ɀF#w֗yZe���i��q��3;�O@3r�9I����P�d[�)AƙȨ#�����a�IL���@z���A�a��=��n2�-"��s�P8r:z�}��8�ݍ3�p�'�ۈ��a�H���ap1����W,��MS��t_���:�iSCecq��@��`���z���5s�.SǕ�����N�j�=���W��S��[WMG���@/�(v��$6��6P��$��I�)���* ��OU�ʤ6ʚJ�p�[�m��L�帺(�w�+��TT	YH�g��.p�	�1�L��i�0P���J��^�d�c��.ua�/}S),l�{�^$
�&P�3a.�^vr��O�z��(I���Mv�GNr��s$@�n�˟Ҟ�)� �@�:D��	{�Rb{�ؾ;r�Q�Z�j��ݳ	IIs�~=�T�����U��^ �A��/�e�9����Ѩ���Tm�j�#�1`�9�w��.u�����y)���M����E�in��~;-\��,mH���IӐ#K�eh��s��'z{����KVݦ����s"C�r�LQ���"{4ף,���e��@�6y�u�Ͻ�Չm��S������C��m�bx�Yc1y��G��V�3T<1*��G����jyxUH�(��:��R���e'�F�d\\�.ݴ8�O�K��Q��W�?$;7&�I�3qz2�6~��$t,

!��
��8�!�4`L�r�Ot�YR[Ui�Ǔ�1A�UxL���@k6^f�dqEbʐ���y���2�����}�0��7Z�1�	���t�<��_o�	Lr�e��4�Y*��ԯZA��47���~[ȠD%v%�(��iJ�2���u6TKZ�S���)��^��r��K���ns3i(�0r�ghb�by�Q���-���ܝZ<~c�wW��@q<o&���hM�����$�N+
�N��ʦt+̤&/��E�@d����=l���M�N}0�7cH|�o��r�X���Yeא�	�IX �ԓ����?��?�	E9yf���-0����ٶ#E��s�#cS��3�R��k�0�w[�8k�?�����i�Pk�b:��j�ehY���Ǐ b�v��X����b*e��پ�bC_�F��,єLOa���.��<��(�U�h�>W+u�lk`d�
lmy,����B�ow_�::T��$���pg��G��A�x�d�)����|�9�����:{������4-��تQ�0�[����4�۳�
�/���;-
cv��VT,�t�Ai���^6(�Ԭ�W!���j��v���}U$�'�����K� ���n2`����$IQ�:� v4K,�Y2�Ό|�k��Ԭ��K9 :����f,���=���%����H�O�?R��ލ���8����%.���W���'T\���R�_2l���T�{�ٓ��g�К�u��\ӧ\Q߉ɶ-��u1S������;����u�y/ʑ�p����ٽ�E6��b+O�3ӻ�ڱS�u�7��ە�$D�n�B���u�4���W[�;�/�잀��[����*wB��8XN��!��$��g��J��;ڳ����"ʄ�����t�1y+����}�2���ؠ舛�4�4H�hF2�2�ȸr�}�y�xv�ckЗ����g�5���ﯵ���ǡi/�cTq���x�k���n.e�����;B� �V�9��d��],�I��$8��s��81%=��5`���}Ռ��Ow%,JD_L��
@��U��2nB��{�­��]%+&��E� ^r�NY�'΃9�f�l��ێ��7QNU����{#@�@ A[�{ش����*��8�0�,�';�ɜ��-�Q�L�+$�_E�/�Hc�x�Ѣ��?�u�N��?�0�ޜ1�;e�5M�����ӽp,�P.�:�N'@��p��Jв:��3Rʏ���3o>�
��΀�K���,-�	?���~gx8#��2���8u�t��L�:�t���)��ֵյ�K�@��R��5�$�6�����8,>�D��.O�ˈ�~>�f��uB��3� 	5�QN�·ݚ�"J����x�@�K���#B�d���k��S��nK�L��v#wv�iFa���T���]2���)^v�E��:�7$ڑ�ߠ<�F�I�D��Pv�F���ׇ�J��_��ƨ�|L���@>�>������x�Xwvx��EO��t�oGѱm����A:���_�҇��!���32��s�1�vK�A1<!��u����S��y}��D@ F��u�a����N���Y�{�`��c�Nq�T<�j��C�9ZЏ���&j��c!&�l_�3a=@�?�Y�� ����$�z )ߘlL��o��LG���D����h(�C�<"׮=d��֤�ͭm������.z�����rC��B�o!�f<�/��@8^����g^����֜9,c^�������~�I�1j]�7�c���-D�D�Ո�1z��2'ܵ��S�+���<Y���ҲS/%��l{P�&�W�$����,��-μ�9%�z�@��t��gu�Zl>�Θ[�C���)����iud��j�۫2�(�$) 0����*|@0�Kr�U]ڜd��Em2�e.<�R���l}o���f��|PZ4���Zި�D��.�Ǐ��D�'<�W^
ыS?�7��\]FASo�X�zn��2��0(3��v9 �lO"1>����i� ��w>(�a\`�z���6�ug�޶.�&�"|��2F�� ���$��	���|��������a.�F�y�&�2b��oI��*�M9Ͽ�)O�4ը~'���nh<a�X==���ĠK����ݛ���N(��yΗ�P��o��0�y��M��O!e9y�.D�?�گ����QW���Uк�x�VMC�R���r�9�v��s꒕�"��� h���@vq(�ڜ	�o�����~��{ƦR��i�.\������-y��š���9��M���n�/��ԯ�?NY��3�mu�COo8�tX ��^N�d��FFu1����^�`eoٛ
�pҧV���o�s��C�ߩW�k��Ak����vH{�X�<��q＆.��j�zu�A�=���<���t����l��g���B�f\��F�^�TTA}�m���I�1s��}VL�=3ʉa��g�S݂ɮ�/#!������;�ZUA������o1hPnA�t�A?�%G>_��w���F��|�`�h�L��=![�v�B>$�S�"X�b�C����Fo��a-��I�4z+�}R��N��>��+�i����VCI�$ږ�g��
��
�n�!rI�;{kZ���,����f�#��Xa��3��k�v�Rp>�ΡoaG�H�H6�3��5���R8���>w�دߵ�
.�皙��J`P�5�΢ܯ=��=~�g�hz8�_�s��L�r��P>r��M�j�>���~\�%1Z���G�#&G���h�f��k���"����U_ _adv�Y�@Td:Q|��A|ٓ�,xk���;7�!�~nԖ�Gw1�n��8���e!���ͦc���l��9[�u��Z�$�@lX����K��vg��66��}~��Ob�)~��~�Y��MV�Y�:�91�J��}N�]�	 D�i����S�)*dR�G<�>Np�F�jz�<SN�a���d��~�q3�v��4��2��������{0|��U��v��jD �9�`�����lQF�njH��X��NHy��+(��:aj �z���f�̳�%��Sh�$0��X�_g�%��Ta���f�`�j~J7��^ۻV�)��6�u`�������4x$�튎j'����h��7!�AH����\��c@���P()H�~�^�m�wr69?��ĉ��l`K�5�G|a-;�������*��ێ��B幷�[�־y����!8ă�\�q&˴�A�m�>`�jZ/ �zF��[jv1�#��J��4��)���)�6!�0?�p �="G��BpDX�:��q��A�d=��K�_f�⍫�L�~���3�A	�����^]�[=B���%�C!��{m�bH=L��B��n��g
3\8_o7���
�j��Q5��	�3�jvA(�}c,�jC�-%�p����Lʍ;p���bf�	j�r��Y�g Jw4%橰Q���N�f�>i�dvѦ5O�{�v�u��d�����3@2Ɂ�+�	B�]�=�_���#�9<��R��ؚ��c\�k�.b*��{9�Qv~�b���;�����C�]㍰�lk�S8��W�`b$�D�pGؼC�q���f�gj1��^�)j��w�/!���XT��KOZ*X���u)���L��*e�3�*2~ɬ6U L�^��E��J\��G�-,F�i2�^���PS~h1WU	,�*��OW���c4�5����Ϫ�Z}���(�ovo��!�:����A��O���BS�W:��U����,�P\�-9���z��j�(�����a�Ǒؒ0�Q���`�Z���q�LT��Z�����%A���8f��[N�S)�M��(�ʡ��X�<�t��R���=fvT( �J����:�-#����Ƽ�;�}y�4�BHk�g�]I�2r�Dl�:��`@�Ժ�p� !l��b�����\e=
�Uo{���/�����g?�ͧ ��4�f4X��+z@d$&��(��s����'Z	ǣbR{�>��٣�Y���a�R�G���q����>@5����X)=(�Z�ɔ1>d����v�rԕ����̀=�쀠��/�ê���/��o��T�9&M�,�~�X�>Bt��Z�r����<E(l������F�`-��gdJ���,Iٵ�'�6�1a�P�*Qy�>-���Y[���{m���'��Y<�|S���<�?����5��@v�{ݺ�([�Nv�Љ+�ʂ���%T����y;Rc:���F�����l]�0��o��8X�O,!��dzH8���0��5��pJz�Yr����w!rII.�[������LQ�]ȷD�Q�����Hj�Q<0K��?��
_֦`�#��U��Hw>ld��ΥJ|	n��[`��9���1��i/��gEc�t����t&�G��k�1E=�M�C�ꦯa7l�-^w�6% I�c}1^|ˇZ6#�����U������9�9&��D�$�\���Z�/�n���#��uF��~>���GT�HtV����,�ͪ.WМ�+�
Z�E:�k��:�rǓ%9O�h�ˣ����e�|E�"z^��b2Q
�w�����@Ѕ��(�:?�dHH?`�q
.q!%3 kd�N b��t%�B9�`�凌@�VҮ&%�߁��D���H��R��X�������m��Qx��}����=~3E��iv�
�<�lcYA>����]�F���g&�.��c9��,��qԛ��dy��S� �2�2W��
���E��"|�U�+�īR�ϳ�L,*��č�LN��n����S˃ҕ���	��b4��_h.��rW���m)3I�\c�9_j���0�bk���j�W�vj�#��x�:c�zS�ꠥQ��0��ag:G�
\K� �sB>.�1н��?�rC4|.f�Im�x]j�ސʣYpz��щ�m������ ��� �^�=��j9�ܖ���+�
r^[:w�br��NkHVF �� �X{��e7�[�j��w(�������z'������Y�1) �ƣ��m�����)	��ߞ��Z�LYK��:9K6W�Y��Cpvk2��z��ے�W�KXSum�ˉ��@Q)WW/BdV�f�nM���Ɂ~��Uv���*�D�j-�Ir)<5��VF?�#�T6fs����U�6sr�Ŕ^K�|45D2��qv뜧=�K	��Fg��D����>i��� D�B�P��X�z-�m|��OS�Ρl��.q���d�	r�0Z�n�08:8���n�{+Ji���߽�YZ
I0&:
�%��:��:���~�}���("ztT�]I���y�ⰖE���l`\7IzU�� V|�H��o5KAn�ʢ��\L�����h>�)���@���M�2# 6S�q��C�Jp�8���>��Y�K��L�����[E�T�����s�L;R	�JF�etb���ٹ�0�������
��S%�~2cx�P�똾Q����BT#wzF��-�W�E`
by�b������1 ��=�dG�BZ�g��yp(��X�蔉%���oV����[��l�����&�QC`��+j���.�x�
�+�� ��ߘ�GY�PO+1�~��Xdr��o֦��:&��~!�Mj?k��Ꮰ%8Qڞ8X�B���rd����g|�_F�4M��b;gw;����m8V v�'��u|њut�~ a|����5���0��C�}���?�pe��3����]M��D���-"���R��GnK{��ŬY c=��{�B';c]�����+���[P�lb�A~~�����f$��)�G�9G�����dP��Yr��"sw�b��@�ij�鬾�3��-(�����3ՇSZ�w=S���iჲ���������n/��/�|�
������,�㲋������f5��/∻�`v�N��}�J�Y����������/:�3��� |,�[������l���V�R�e�:$�3"}��>�zp8b�<�B)�DݭoJ�&�US�r{A��xa-�d��cLt�m����,3a~�zi}�].�8M��i���G��s�*��a2cˢ�A�y�Q]e�e��/��D�\s�O�����G�ji��y��Hwpq��w�J��J�l:^4���h�?pKr�ڃ��5�5�|#�H󤆧�w�~�}q���"�V�h��|��Q��}�F�ܶVE�iI �#�T,����Ga�ޑ�{i0lfuRS�.,�iy#�ٷm)��	�=���|0OB��I�E��=�8��C�
=40Q	<�Y������Ս�΀�B5kYN<P5����&��61Y�J))�w�R�e�q��l���p?�+r���]"I�;&��ֹwx&f	�G.Fӻ3�h��m�� k���O'�X�4�jR�ܺ��f\��b�&�#-���̉j[e+�\%���y�ě���0�B���B���K�)MOrbF�x+��(<) �b���d]@�����+�;B���ɸ�X��a�L%���M�|�M�l��c�� *3����|�)4�{�8���!�gZ�H �6Ƕ�\ݳ����p�K��Z<�e��f�tVL+O {�	��{6#�c��Cw��$�=��=�ֈp�
I��uJ��Jf�T:��S�b/��m��-������(��Ě�(x\Rq�0=>PRo�=�MӀ��#;�����*#1Җ^u�Y��5��Z��+��̒`��d���� 5`�+ESa�IJ$ϕ���)��c7Ѳ�Iѳrۧ�x�:�0�8����4t�$�]��'� =麃���D:���ha쭑���&��2'����)�b��k�H.��cl������4{�`*|Ñ�}E-��!�����'Se�Ԏ4,�;����uЍ�gR�O%���犆M�A���@s��P$��%�=�]7����󯄱Ly[�9�U�W�6�-���d�'@�fhA�����|��[	OH�u"�+-ֵ�}v��Y zy:��l�uTT_^$�5/��í/�Y��:��>��,�V�C:`�h�1��#6��H���Q�l�����%�_!�C��bSC&��N "AG���v̿�b]	�A�Z���u͟EU*�ټNJ�9~k'�TNQ
1�NW��ǁ��,��nP:"r�G�Mg��9�~�j��}Z�7Y+���H����Y
�/K�-�rM)�f�Z�&@��)�h�;) �V ���My�]"j�};u��(0̣/JѺ�퐒(>� ����0�b��eۙ�F;��89�ď0!���cP5*Ӌ���r��]
OM����s�]���GV�+F4�D��]i|OA#7UDK��~U�����"��@p�OI��V�M>�H>w���U>ц��s����9��X�- ����V�����K���ϡ�6�N���D����������=r ���Y#=�KD#d1��yN]$偛������fN�=wJG�q[�9<�G�3��֕��27-��R���nAOX����0e����+�Ƥ����9����9y�n9������%yD�SgO�ދ���p)Z*�aq��Xٔ«��&g�{�+���/w*�G־�k� ���`c���*��F�Mr�a���#y��.�W��R��Ul��U�/r*7�����΄�	�!���c��Ȓ��ٞ���y���r���Ug�ǝCN�U�e}�<ͳ`�� G�5�s�kg���酸��~+ӓT4';���'OlE=�9S��F��l�����h�4C?GG=��s>c*���mx�
p���<�IJ�ܧ�#�������ې"�e�X{�K蝟W��_�l\���yN�\�M��~���FWt�2�+�������"\�J�v�]�Κ����+��ҤM!��h���0���E((��k� Y�i,8x���|�P1O/��݁�t�%|���.NB}�N/;�r��~)|�[rl�	�)����N���)�!}�"����|�͘囲y��FʧZT���D���aC�B�I��)�YD���=������[����[9H�*�X����� sM�g��2ؒ��"��-��{�w�)�,_W���{,\��5�;�W���,�* sdi��X�|�}�l�KI.(AE7�s�W0�fu��X�\����ػ3�H�L�7��G�<��G�Ml�R0���0���Й�C�Iΐ����at}>�>R��Ў�F���t�@�T���u�o�G�2����斎܌�~0�N��$t�}��4�R�?�P��<�6#����)2<7�AY�=.����{�RS`*�t?|VF�W���<�ީof�
�q��)��m'ed��1��#��rs;�DO&�\Բ(�x%�7��x�Z��V�3H����v=�->������_s9��s�ǹ������sFLө)�V�8v�C�US ��IR�(������S��!7�p^�d̥��x�y�⻯�J&��N�~��	�����3�_y�e�`G�κ����J���e�9��m����4)�j̃�����#���ׄ"�y�[X�8{���}���sE�L�x"b����	�0�v��v��v��Y����+����%A_�ݥc�ݠ�)�
Ͳ�b�Vj�]Gu�t�~[��
'g�pje����&n�8�{>�Rb��$�8x����(�nX�s,b�k-��K�g,��D!�!,�`�:����J�;���r��&>5D�T'�Y�i�G=Π*4�Lk'�>��ٜ�OµH���Z*`Ç�KT��a��B�ԙ�u��{B
���F��PR�c8�(�C��NB�a6f��E���&�1J�t��)�=�l@�^����fS�)AX�l	87��g�$�6-�7خ�f��`?%�W��c�M���9��q���a������K�=0�r���d���`���P��A}��MV��+�-(�E���7ř����q���x��D�C� �Q:pb�+$�W�t�l�h�� M�n�9����so��2s(��Vژ�&
�;�xX��X�@����	�o�	)M�gјv`�W��VLpk�ۗM��W���Zr��l�(Qf�x~�Ҧ; Ԑ}���������+�Øc��"�*��x�T�чz�xiL`����c�<�@�A��X�`���s��pg�-֍&j���)����9��b�Fe���!`���s�9���*����<�(����-֋7ҕ�̂i�Μ��1��ǚk�S�0	�����j9�l��T<u| ��Zc�Hς�' =G��(�͛���.�i�G��a�]D���A�g�g����"D���_��GWT����\���)7�h����W����\�.+@��d�(�tN���2ܼ��d�bh��»C��̝/�ɲ���C�=�Z���b.��D�-t+b�jx�XUJ�L�g"`N{ܳL���V�յ��+����C�H��c�bBۜ��z�0T����k�e}��V������Ў�DB��}��Se�7f��Җޠm�s,�ܗ�����gv���2�ݨS��;'�ٹ��ix4 x��Ks�y_3���T/�ԥ��E��!=�l;�1<fz��)��c��l�2�eU`��k��)0���ud:�B|����:i����9v���ej)����H����,�ߗ�=y�O�:�b�<٠�o�@]���w�e�,�195!���C��s�㻡R��8�/ҧ�;V�-�Hc�^�"�;y�-)��!.qZؙ��QD�S{�
F����̒��8O��6E�p'�{Bl]N�z?�����t+�y%��\�$c�Al�k �r����6fN)~S���4'�ޏ����rB8����2�K��M�����+f��n�$�T�����`�2M��
~ds��m����)a}4Ŀ�6��C|:뭤�9�G8�@���6qW����xz��)ܣGBM"�D��3Ӯn��t����6�]�.~$���N��;�t$���:� �`a9V��6�j�S��e�i��,nIDZ.�I ��@my��8�����Zs	
a���y����(��X��X�)��_>�1����0�c\g��K���HZm<��/�lEj����������D��(s�;���S���s	>�"�?%lXͼ���HM��Y���jgh1T��]�w(���&���)��%��3��[!��bg����yg�&��n���R-3) 8p0k䭟�O��йB�;goH�J�:�P�kվ�N��ߓ��&B�����%P�Oa��.�.,�A\)#L�?��r���$��9]�Q��ܤ�f�L� �G
�ג8�[�m,cW�G#�$�L��M�~�eלL�
����I��Nt�l��J�["��	|� �H7R�N�zvaxOnxB����-5�R=&.���C(ƕ��їX��}������q�Y��#����������I�����0z�k����z�&�n��.�,��������2*�7�:a���i�6�zha��d�+��wS�o&�,�����t��\2��7ʶ9�]��$�!�)�GAӗJg�]�p\3Z����FR�D�޾+�?�R���ǝu?�C�����T�a7�<byt�@2����߿�D�'��̶j7�Xl��>,��i��0"�|6��Rg��!`I��� ���,�K�H�Ld����@�$����S6�<*������j��3����+w��?��L|�e���jF�E����؁sv\ܧ��O��}\U�`-`�5gK�q炱�lt�w�i�)�ӱ�=�-B��1��ҬÄ7$��e�r��%�{�&�Ex����PP�[i��T�db��|�=lǍ��I����xZ�B�PRW۠S]�w�&]2d���)�8߷�&$(I.��8���h���)bd�$�HM�xV|u5I�@4�LlU���:�ڭ?��u>�H�=.!N�'%RI+�):��qb����C�g��8]��S?��:/�BSM�2��(�����љV����3n��ϋD���Q�U,���M*��/���9EtC���A�C��d���*ȊImb\1���ci1%�O���`ֳxy ^�1B�� Nֳ�9jm� ��sbI�����å�ŋ0P�Z���Q�($ M�_�d���M�����/�"��9�&�j�cQdb%b�?T�tC@F"e��H*[�Z��#t�.`���YN�y{'�Fދi�k��>�l�|oX ��oZ��s{JdQL����;{��\}A��#�`+(�@h�1�<3�S$�b�K2�&C����]�\��C��'s'��#N���4��`�S�Sj1�F�t��{$jH�.�G{YN��ͮ\��A��qO�79�x�Ͽ�	i�}����%�-�j����I
��si�p�a��}�v�J���T�uᮃK�O�mcojP]�b��I�kg��ue˦���r�|�ċ�Y���`\};�w�S�I�b\w����'ad�o�[�(2��˕�t<��\-W����_��[�CI�rvנ������g.�:d*�݅�q]M�bE�����W	1m�yN��tНӽ\92$���[�g��OEG�Cl�М�蚚%x����]3c�d���u�t+& �Q�����zP�G�H�9�����r�)K/^�a��}�?Ţ����s�
յ(������^j��d��"�=���ݶl���6
�{`ֺ�)����c�B�{-h]���؆̹~9����٘,bZ�	�ډ����{�(��EL�Ү냄���eP���=��5q�7L�t7�_��C�˯��T4ϢWR����XK�8-!��/��hJz�\jҤ���9U�9�$��
����=�8۷U�Lx�ۻ�H�
AF����"�b!c"Y���1ؕxT��N���N0�r/,8p���}�U���eW�M��g�&����b�@���bK.��2� ���JM��L0�ڦŪA�\G6�$3Kl��/X5�T/2%��$�>ʂ���[#�&����MZf�/��ezZ����2���$������7݄w]F�-�Hd�0d�s�z�2(�d�2���vPJ(���p�5t�{R�ڐ�j�
�T3�7����D�X��h����G	�����	ӧ�ɒ����p<��B��9Y�����(�k�^�_sF��#ɟ6��[�g�~R��?�d[&5���҈��.>�Iƚ���`�@q4�V�p�5�0PA5�Gꍥ�z�_���|�������5qݪ��V$�op�9����������ld�rS����o5='de����̦n�?Hy>F4W�~��yw��'�UZ��w�;H?-"=�l� ��&7i��Q�M�F�l�)W{@����U|���ŗUJ���Xt�ݲ&M��BP ����NC�Ȋ&3u[����� �q��M;���5`w�ϰ8��y�-,��O�I+��b�%�s��,�)��+K����)]������8,l�/����&\
��]�y����9�t9mA���
��f�S�u�g�l�W0&<�ן�s�F��I���D3����;���Sy�42aUPH� �����Q�2R���%B1fЛ�,v�I-w6�� ���Y��%U���1]0E�?�M_��\��������F����W_�F[���O梞�����hoJX_�\!�V��+����
q�Q���{�d��_8�����04	AT#B��r�k�/��2�~@g!�c-�3XGxP
�c5�9V�l2~�l�+0�!/��9ܭ��۫�֜8����hC��E�^�"L0�σ�b�h�.���S�Mٖ�V`����ݞx�>h��≨���ˊ?���V����u���*R����^4�+���mc/�g]����SHv����O3o�˽��ǽY�����kb����Ř��_J�����{�F�Ls��p�!��s���ћ	�ˠ�,ߠ^����0լ���jmST�vF.�E���&
��е�X���VbJc���y[}�=�b��Ru�
1-1'Pd��+�d����;4:Pu~����z��y,�&H$�ר�1A��݊&��ʦ*�sw�z&���������?J*���j� /3�����%�f
)�p"	��q����~����v���*Q'�6lAaii�ǐ:�J��4?$7�!�ɲ��}�QD�X�Z��|p?)I�S-��G��J�q�w�����0�_���ho�Q-;?�s�9!������M��V�Ӽ5]W�0����{.;��O�7�)����u��!��Ι ���w�ζrN���v$�&��Ț�$E������9�B�)�"<!���Js��<�-���Ɵa�I�&K{�ih���(Pr#�{�%Ȭˤf�"��l��rB��d�H�U��#����U��:�:������Z,��1$��Q�x��@/�"��N=7{�:,�O����*��G�b��=��@�Q�C�e��5�2Jj��!�r&6�/0p��
8h�O`̔�D&6�}���	���mV0n�|۽K��������uWP>���!f!��S�Z�٘�y(4|�	Z�ҸP"��{q��
���^'����>-D��˸�I:��"��`"b@R]"�g'z -	Ew�Oe�b�w�e������=殿~�;͓o��o��Z�UY��Cܕ}���^���d݊3�fH�K!�"-��p��G(sIK9�6p6����YA9k�O��M�T�)m��3O�YX�v��&Yq�Ri�'�Q)ѭ�/|�C���1ME�v�,9L���:À�=eUu�x}O�8�@0Jo����\�F��@���?���#h��=��0�L��'�m7�F�ahw�F���s���b��C�ƶ�p��m�	���0x���$��U��I%�x�v�n^�,���"�>$w����2�D��ḝ�u�]�'���D�4`R%��
O��I��?��B�
P;z���K��qTd!����p�%��0�:.���J���ŝJ��!�DmJE~���7u��P�98�'��%��8�Y�8C2�ټ��=X�ӫEG�|6o�YAXԂl�'���rI2�ɐ+`��NZ�)��w��!�sa>��yʖ�7F5*C%W�ݒ����<ŷ�)�����G�@�5�ޘ4�5c�p��R���Ge�-܄�ެWͅV���+��pf�&H~�庭�s ��6����&V��43Q�7��W��-h_v����o�oSXY�V<�z�NoJ�Ы�U*׏�	!���$���z�����E�	M�<K�xѶ=�Xw�
;g�]�����6#�=n}��O�w�x����G�l?��	%�t��#,��TPQ�����ޑ��U���'��|�Ő��A�KIU��Pk�rS ��[�����e�I�]�����o�M�8����l	+B�AH�<�}M���[,- U:-
�����p���uu��q��v7�t���le�Ǹ�͞Fx��q]rVO�_�T�t��{kJ8��s|5��9˩����o	:~(������g_~A+E�ԐfN!�!~��:�r,ۅz�
� n�d��E���r�j�O"Wz��N�)C�����a&?D�Ð�.\M�,�L�1�ns%�c7OZ�����/۶�奦����6Phk��Y�-�a������^?���ő�5��ȶ§�`�oR��u�֘�61¢,��������nK�s��0������Cg4�����q堈p�b��./f�\`��xa�w��.�Ӑ�~���pf]��Cnq)V��J�Pzc��z�;�������h��97������vpܔ�Hy> N�$�"�W:tva��U��[��G�)�4r��Ó�SD%�0�c�m~��:������c���ak�j yn5��~��N�[D�
��N_ѵ��'.�yz��{@�d�Y^��Q���wY�L*�i�p4�^�^��t�t�8��h�D���������r�n�y��'�,5�km�N���i),�Z�i�5��߷2����ҫ2F~b2�45����w�N���%��ۮ��pF��v�)��j���{NiS��&��� .H@��^p$���g����F��d�+��iz�����;��u��ZZ��7����n�#�=�d�4�� ���2
[�S����������F<H��D)�,@��n��L#:��%��Q�*?.�N�Y맚'\�8@HJ��:�;������~���DtZItW�R�)�Oh�����7�,�sIQ\���D�X�����9f���+�}���nxOu�އ.�e�R]ȋ�r�E��P\? m�'N����hA��;�����á�Å~���"��A������o�J
좙܍�1Ywlk s�q  ����B���X�v�i�~(��ۨ�J ���v@�q^�[��p�IŔ,�(��e��ӗD��%�Y�𤚎�!��T���(�T^���"���>��r!�I�U5�"C���+��e԰b뒆��o��<�+8��e��%9�z�L�O$*�2�H��a�R����|�J�=SQ*�m�eIDV싾��4�cq����p��I1<��Ք��-m2���f.V�k�#E̷2������0�IoN���B��P�f-�l]��@*�,�+��.Ο����p5��p�[f���oƦ`�_��1'q���jB�;7�z�] oCɡæ��x�jYg�0��{R3�s��֒�r���N/f�V���w� ��#��}"/\-����@���B�nȗJ�sa�L����s�0��3�jqC-X�`�&�J��8[�h��A�]�u�$�t�ۙ�>������Ԯ��zg2`P��O�����[b��7�i)Z��&�㱫%y�pam���W��U�F[k񉱠�eH_.�p��J�q�"J��do�γ1x��f]�1�'��Ns�]R�ȋNj[��i{(��z􍋵 %~L)o	���*�G!iC%$�'lT�)��ɷQ��4�����]7������5�B�E=,���r����ϵ�� �oC�_�=�M�A���D$��l�kk��#�C�T�ue�F�"�t��T��gr�C�'��_�}�E5��<�� �S��J"4?�˙�o��7�}Q��n����P���a��3:���͊��mb��C�a��*���b��m�N3QQ6��r|�����m���8<Ψ�j�:T8��_�a�(����v��dh����"��\#J���l�ͦjR�q��ß8����x��o펞��^H9�8���:�3��P��h����:0��hns�d��7j�9o��S�5�JSp����I�-<Č� Kgm+���Dx����\�1B�����n�ӥ�6�Ft���<\y��"����BJ����_��҆����jU�*u�zc�
���:9�:m��"m���oPH�h!��^����sl���@�u|�^)_��_r�~JE��s:<����������a=�>�P���|��om0��\v��
����
j�52ɂ�0�u�Q�j��ҫIT<�>�(��w�>�4�c��P:�O��t��Pn2�h8ֻğڠ~֭'2�sB���љ1��Z��)z^D���E�c�J(S�=���fҽjy��O��nS3<B������Es~
��b���kѥ�y��s�&  9�F�߉��Q�_����/5�ǁ\��4I��tU�n[i~]!� j�q^9�/�"����>/�M�C|� �M�&�� ����f'����O���P�C8.�i��o�_���9b&/�\G���g��{�ێ$4a��.8<ǒg��C����T��0�O����JT� �޵�\nб;���p4([����,��@���(Ց0_�}RM.6���6б&��JIѠ��Ǳt;^ߢ��ըm�����!�ʙd��z��d�����ŀ�G)##F.�i��I���^���g}����ߨ�*!����ڽN�<��ɜ��213e�d�f�ևOCn}>�x��'�,��n���/锻8�Ɉ(���.e��/��M,ֹQ���w���aê���+uٶ���� >�3-H�1�`:8E&�S�y�ˋ�7 OB�L�HTY�?"��[���T��w*��:�C�#��{����¸�;��w����dI�l�<xc{U�=�" �Pe��uf�����hv@��?w7ȕ����	����ev���s"���̇])��Sٮ���`x���.wءجܢ�Xֆ�M�O�"~͗'�I����?����)�������q��I�>ˠ�����rM��G-\������%I��E���`�W�^$!;�Z���/��}>�5Z표��}Q%3��|l��ī���V"=7�-�a\�C�E��I�4A��\�"I,x[����V2�Ɍ�pXk�S>S��SMF���,�dY�u���H��?Q�rD��}�זB��Ѽ�͟�%g�l�KB0Ė�3��-��H6/9$�Oh���w��3Q`���?�i�O�A����5�̼~��ǜ�QaN>�B����+N܀w��waw� l�����G�r������n�
C�1@;O7�=��/�x���F�VauP���,-���F���/8�k�%6\�[-S'����<�B�m!��h����"'p^�0k6(W&<y��b^{�����{�-2�uO�G_�����n`�b߹&bV^��y��ڥ�;ΝSH�:�*��W�Ş�s�������p�{P<�$M8�4"��~H�z���ES'���\�O��wo�.��y�2����4��o;�^���b�Н�7���t`(0������3�'TY��*�s<�q��D�3g'��2�"EǼT6ܨ��,F�hV�dCLʖ�7�d��-�S�mi<��Ҧ�\�b^w���^�H�Q4�Z�u���&~R�OR'�o)�,��aJ�A������(����&�����Y7D8���,ȥ�AA*miz���M�bRAFL���,���!l�Hi�~�w�nٽj�1ߏ���fg�� ;�X~�̳�:��M��t<_,A" R�|U������v/�s�e��^H���[ΦYy��V�)���zZ?P�[��}�an���!���&p%$��Q9#^��囬�F���'Rzۢ�ƈ�$�rI�ۅ�E�x�K�%��V�M|�"n�?����bV��D���#Xu�^�Y��u}|rGX��]AU�-t}�$B���j/�9�d���-���9���H�=u�����`Dr�����,�9z�"�t �=$�{�{R@�x ^� �O:=��uÑX�''�ϒv�Ӊ�[u��~�s��ߘ��Se|T�ZT)T)A�B���hG�����������Wu�4�sX��.�^���EMa=��hč?�|�f�y�Rط _�EV��3����ĭ�N����R]��k������CϔxLr�������Ŧ�������B��l~�����i@���إӘ�]LdIY�����P��5����5^HˍQn���p�,��nO���s�).���tW���T�3�`�=HRw���^bձ5�F�W�<�5^��6�՛p�C~��=��+�CO�PV�����=f�5�l#���A<E	2�Ew�&I��i��g��_?k�0��.�D�"�е�n�ML���%��-s��s7{<�UҦ�SM�V�X��0�n?���� k8����lԂo��#�Zui͝���a~���K"/?��5�F� v$nz�����a�ZS޶ՑiRz)^{��Z�9�<e�r�~I��ێ�I���A�r&eY[7���y��+��t@:C]��V_nJ���땒�Z��r./�~O�3��_�P��Ɗ�b�:_����Hhb����Y�&Ы�F���]��z��9�9�D$�%�|v��(ќ��mq�<KBZ�ZuoH�QI{�6@Z��i�.qOUM�vA�!�f�j��Vu��31���28���\kI�ט�ܳ�x�W�D�,���5��b�[�q�������Xg���~b�b}s
2\T����
��_�4�ݿ4S������<�iU�K�-�MgFY�G$��v� ����3�g#L�z�y��ʿ���Ľ��Xs9ah��!9��y�'���F[!�|���'	_5���+�3�?�Q���8���hMtJ&'��3��ˍϤ���+�*���6���Pӳ�ŜPU@�(9Įp�� Wg�
ޮ+{K�>� t����JG%�ug�o�I��G��:��,d|i�7�4B��QÛ\vC����]�S�w��P�%�^,�\/9�Hl��l�9���>O�Kag�^8V�G)��Y;07�Ҿ��m�-�J1Uzg���
�g�t�\�u�i�"%��8��y	�h�I�w�G�K�_�~f��5%��t��Y���I�L�S�mV��rQ��Ly��о�à��e��S���<0�n����z�;����4,�ܙy��-�!)pp;K�7���2�_���K~�Z,J�k.���t��dU^`;2�=Vب!����6��ز�5!��N0�:��9V���,�o+��B>Zf�6ޗQB�nCێ��yR<d&��A$v�����ߵ����6�3]g�?Z��AsD	?���9�\_��jS�w�0;�(���"�u���}S��O3�+�l ̱BȲ����`[a��:�`�/��$�z�	�C�_WC�`���B��\8i�aV�	i��|�}���TP}�7����q9�P5>މ�@IZ&���KNs�N�@���#�?�����nw^�X�4���߄D�ބ/����K2I��,�Ւu�F4���Æ'8�{-O�A��>t�����N#�m��}ra�jiMN�T<�'dN�L���ɰ�X�N(٧���eߤ 	z��?j���hY�|&�"�0(i,�}�)����jB��\s6f����,�>p�}�񅺥���ج]'g��p�%�f[iF����(���`�g\���Q'���D�����[�wDĺ>#H�����IX`�Q[��&�=�x4���޺�iJm|[��8cG�5�Ug�HL;���&�9D��*b��j������|�T�&?���,�_�)�迒��:ǒX�hb�*�
�7Z�E*K�$���[\ePO�R%B��`�$x=����w*�܀�����1w�$�l�xr��^=q���!�֟�A�S�ђX����u6^�u�A��^�>���<��oz�@랪�����O�D��*ފW�~r�
(� q0�s>{<:f:g���L�Y�;�G({Xi]��^n�OG�\\Eˀ�"���^�0x�EiP��GkOw�fR��hF�c� z#��/X���:f��&	���u��#m�!W��nb4y&�w�������?��#|��H8@�h��i<�vZQ�r��Oad��'6~���q���š�h���-<�π��&�\�u��d;��}�����C�s]�S-!�x��vo0m�ę��[��n�8���>��%�F�$�B�H%j6]��u ,�����lۛ*�ߘ�U��]���`+��I�9�����9A�������G�Z��Z�]u���>վU��O儃3� *5b��eP:)���ˡ������U��2�_�g�շ��o'�6Q�9��ª-'ɯ&o�A�7�=����?���@�S�š��@�ڔx��[�,�0xRm�r���x�W�pK,�3��x���Nd] �+<��7���P~������H�p5�y�ظ\ޘ���r*s�|�sU�m�3��.hfTJ�Bh��
�t`�ܷ����.�gw�C�骿u^��=��_���z���'�� i<�8�l�@����f]��^_8>�ߢQ��
/�[L�=a�y�L)|�w�徂��󑒕?4*	�r�Pʙ�'f}Z� ��
ŏҫ�^�b���ݎC8��	��A���TH��D�+� G^<��B�|ӹT]l�V/w��������� ���A
��~���m`��o�LS`���/�H*��YO?��&`�轒W(���0�����q|����JO�*�1D07��0��[$h�dꓖ:z^��7�����s3�4eļ!�~z�{gH��R�?&��ox`��v����T�,&��zwd���jo��JV�@/;��zF�$�c���[?MVE�����P�n��,.��|'\�6��ދx&G����'Q��,Ǜ�	�����]��l}�zf�}Q �����.B|Fth���Z����-�Xb��s�j`i��$D�����	�=a�D��Ah��턎���������j�8I�V���}coI��^����]'���'W�W=@!��]F�@��4�a%*�v]�(�����v=0���N\G������h�$!�;��h�7^��õ�W��=hW�1���Vm0��f�8t�Uf/��w�M̰5Z�5>�{�\��+�S��L�ZY�3w{�:w��l���E��<���E+dax.�@��#�A�׍��	�Nxb�l]��ܲ<��Vk��5�f���xg��a�V�z����H�^Jm�H޳d���c�RMzZ��"`vL^�d�~�R��6=d��6FZ}�=V����A9N���|�G}@b�SN��ҝ�Q[hd�k�s���.�<�m6�&?\w\�;��*DaC^��%�9^h��a�rI#����Zz��&2�@CWyk��o��z�\���dU�@`��l��Bo���"�:����qׇi�RH&�8c�O�v��.A�(�E&���#Cyc`�R���3���<Н蚾I�s���v��<�^o~��j���)��z�tz��8_߄;ѳkY�!%Vs�m��8���N���:�$*'yL��c����1�9����5�͈^k�c-K;��c�*�1FA��PK�{B�T *����x�$`Bcv�Fpw�L��YʣC~��}�*S�[�o�.�?�(I晽1�����2�G����b���讧ۦ���R������b�1n�Y7��J�S�zS��f�z�qRy�#��IO��޶��U�y5�����\��I
dؼ3X���} �/�qwO�u�(�˙�${��c�෷��G�"D��>k�1�J*�a���,����ݮ����ҜDo��K�ۙ����ynQ�:���ݙ���/�?X"K����Eۗ0�-ǻ�B��o�le���n�̶�M��@Ey��@�:���̤\����'���9���F�Yi�Ȩf;Ƣ���ڐ�����TiS��A�w`inʤU����B�Eu���g6���Q�ʥ�!�)��l�c�+!hB1�f�ȕc��[����	1���]ᬜ�L�Jb��O�l5�o6v��U�~W��q�0���l-%E��o��>���x��W�6��ǅ���O`RϙK��3`ǡ[j���F�%F#�D���t��J��ȓ���@���Q��J�	c�0�,���Ӻ��f25~�6GF-���_��z7b����0�l��'��_�*�2k�྿w]�������>��=�i��rt�7��<��d��]�ƶ���RN�qAJ�[��:�?��),\�;owԴ�Խ���)�*�A��( 8����_~���	 �gS�8(c}"��d�����`��d&Q}?�rs�(���Lc�'�q��>g���	%�6���C*9}{��MϺE���a�՗-����J�{��m�RB����ܬ�SvH�^R�\����z�D�u|#�w,�,�u�G��Jek�w(8�С�A���T��n��YN�g�X/tV=a�/�]�F4E�|�x�O�L'�T�Egg�^�B�T��fm �_M�Ui��?]��=�T�-Gk�!�����x�B�O�`�A���q�؉w������"Tx��ǎ��!�~��3��{�ksR�$�"���uy�UY�]V�w���J�����Q4/���X�uC�n��:��i��Ch�2���J�C<��Bwx�BraC�(v�h1@-�
	��°.�$�|`���u���uE7)�X�l���N��lw�s����e���HS]+����#$�����Y,�!��g{E��-����g��8ze+�b�![@d��1EY�m=�p�ȥ�Vз� ��7Y���1���P$P�M�����֜��!��]_��?���6��R-0�>/���䉯�Y��]ԉ�o$��g�σD��(�Ft�a����k��&CW���<�r����"�~a��R#�L�3��.>��y�����$-s)e�Gr�����֐��!�b��v(M��^F�8�g�y��_�B��x�,?�㖈�[�6=�Ls���+��Fբ��`�����J�j�3��ύ�`�0DԌ#m�C�SR�b��`��ӈɢ1�\Chj3x"���ӑ>�h/�S0��0��Ψn7��#�R�:e���&�􉪗9��ڑ��0}1��y��;k��|���^r�0��h$Ҋ*�9��'`;d�W�����]6�W6|�8�8����1]i�=.,�Wg�����\?�~	Hr�s��T&�ܥ��k��j�bp�V��{�392D.��6Z��ěL�-��,�z��*�������Zd9����)5�t9U/��s���z��3%���T$m���NPb1s�F�u.r!2�Y�F�8�Sk�fv=>ó�>K�}T��K�	+� Q	�;F��!���IK���3^�uo�F`7l��b�h�@mש_G�����q�b�l��v0����D$L�	4W7v�O2��H�;(D\�B!���9PV�&ʐc�ܽӹ��&�i�|�T��Ю3%�ͤ�2���=];e��޽./���d��Җ��-���P���`�L����rhݐ���]��1��C՛?;hd��	7qͥcfNx�ʞ���������-X�v�e��&�[�����!�]�T���p=*�<~�87��q��h� ڢ���-]-Y�Ց<��=�\��>S���S���Lїs"'WQ�K)<=
�8{�,����V�қ��O$L�v����Y������Xf- �ˠ�
Es7�Dª�4zޔ* �TZ���Z����2u�s��h��I)�	X�"F��<�lr�4�\y@�b(��ZD@P`�`��)��p���n!��f�vy<���$ݠ����������_��	:O�cy�3f��&�c\ѧSâ�e����s4��ʳ�?|[���,��
��}�`����i f*����姭t�z�CF��P����n�wo��:-�pZ����j�Ҙ1�C�	��TLǐ/�1]�N�̑�QمX��E�(��fq�;r�z<�<D��������6&�_p.o�=W;�[T��X��g=l����x�DI�7�����e���ni�P1�y��J��w��t�7Eaُ15���(?��16{x�� ��?��֋㘾9u�g�����S�Os���V�z������">���m�'UK��x9���f�0�b͖~��~� �q���ܮNS�4T˺X4�����L��o�.������x��J�46]�Ծ96���T�*#3�,.!eȾ���P%B���7�
���{Q�p���G&*��2����ŉ��܆I[��M����v�{I|Uw^���?իJ���DLZ�	��B�������I�1��c�G����n�k�ݨ��"�VXrw#�����1���	�� �����Y9%`���)��$@���.�VU*�g��=�_���!�&5\��^�T�7�V���
$�\��Y{t>��S�K6Q&��@'���P�c�S��VQS���	���3��AO){M ������b9��x�'��-D+]�P�J����u�;f���i�@,S�F���� p���h;u�ő���!FFۍQ�*jv��'�:���{%��pZCulIi�'Q׻D ɶ4�a�!�����Y�8쪊	+�?g��Zldo�����r9d�Q{��Ap��v/=��l1:��M��7�LakA����ym-��,#-~A�X�zVNjk��N�w.}@<ұ9T��.{�®'om�.W9�E/\��N
��d�mwar��#�DW�4�}�H*��P��5㙃��0xD�q`Cs>j���u=�{��V�����9%�?�1x�0�%N�T�ްAχ��<{y���l�=�/9�\5U�%+��BKolv��\������#rc�+55���
���]�	�#��{:g[�D�ֶz��B-��߇���� �)N�(�[���BU�P����_n7��=��>��]�������X#���a��e5^z|��r���,��/�Nh�=s�g3'�V�RQ0�{���e��Ӧ��v��&E1I��$K\J���~KV׎���S���J0 Bd��F���2��+�#�7�'����4!��D����^W�i�������~y6��J6Sj��I�~06����4&k����M�Lan��1������.L���?�J�1iw�2x�����p�jTU�n>��3����E!���4����n�X�0���~�y��fg*�p>j(;���2)Z<Q]��b�,j�/!��`�OL&5U(sx�M5���ʤo3�},�uHп됨�,)�CM�3*�:@�CB8����hr�Z�V.nYwWWIiK�*I����at TI��;C��K޳��d�(/� ����RH�?������*~w)�T���U�<�sY�2�B��͚zW0�D�hg�3�\��k��Hϻ��GD��E!��`�Bw.{EU�B��a:_�=���"�D`��fA�}�^kU�r^��T�[G��Y�2��i%�VT�A ���Ǚ���E�􄀟,����-���}�+�W]8�!eɲ�r	�:7i-�z(�WvIPH]�^�)�5�X��p�!��R��H> ���ն�����k
���/��5�}�czC�[^��5�"_�����\�i�}|fמ�QLXm]
oEԱ6��	���3=�3��{��)o�@�� B�ų�э��"A�ki�H�zE�OP��x݋j�%d��Ҙ|n31���� �txu>R�{6�g�ʽ+NU���d��:N�(ڟA9���A��nl%ć[��.��d�֬�<��?#5��^'�O���Pox�G��5L�籠,0�<��Z�B�d��X-M5�BE��K��HDy>�ٻ���T�@ft�+&Z��]߂
SG����[P=?F������ޢ�7�һ����E~�㣓X��0GqO��\��	$�po`���t�[�am7�� �t�=��7�S���d�Ӈ4���-�y���>�M���S>�_���M4�%�ZM����W[��^�/�,U�����U�8��:1e~f�Y'���w����^��+��|��K(���ӜDB�X��� pOwߙ�R���nљK�]�ڞ74ױn��+y���ġ���G����g��1�G�yٰ������+7X�9�����Z���!��oiGU���Q%���)O��(����?������r��b2QY^l�ƀ�y�^Bj���zt/fvu�g��{�[����"�xّ��;ɰ�*����FKs�nF1a�T	�/ɜu����k��zxu1�tlm�z<�:�O��U6kodg�h4"�T֖V���x��_M�R��(q��G�g5G���-�D�6�2�/��=�wlVB?ل��V���#ҬK8"'ʴ+S��}	ɷ�ض\o�$X�sO��:/]l�jܰI�o���8B ω��ߣn+�o,���8�,�YK�N�,S�� �x�QUl��n�|`��q�B��Q� �Ӝ�����D�2�	�Q���F�����FBP�_I�vFX��[5Ϋ�ȿd����Y!�bQ5k§{Ֆ �$�Y���`E΂��c��{���Z�ҫS/��m(jL�RN%FH�Gg򑍱-O٢((�2�o�;[�f=��S��f9nY2��1���v>ݫ�d7��u��!KBv>���	�|-��'U@C����_:��3[]n�=8�VI�e�#�-��p�6odc�<�HTdy/�>UN�D�4����輶h��j#U6�dN<�,�1/����f�~�p�2��������R٢ɉ��.�+x՗3�6�h)���ޘ��K+0᭶��ˬ���9����+�9��0ų��s���Vd�A�F``'�xs ���7aD���(e?��alY/Q����x���lA��I��8�,6��S3ؤ�JU��;eI�(C̬NeUQ�h�łh�D�U?�1<�Nd�v��������CdV�&�Bq��`�aۿP����pظd-'�\�*w�1؎���?
ݼde>r��eu�1t�V/�a�5o��:��l��{��》� !�3a�yٓ�5E��(	7|�G O��$���r�p�8	����9�С�o�0�ڛ���0:D&�(�B"�"��le�Q���4�)s�i�̤e��������UtX��T��.�ޅ$A�2��{C�!q~�h�/x%���i�ł�F|�0����`������+<��RjI�33��YЦ�М�3c3Yg���&�g�Φ�a���萠._Ѣ���@�u��a|w�hB�M�x��L9z�37< �ܽ2i`��F
���ų߄�IFr�u�`�j �Q-��q��Ce'�֘�cb�4���-���ya������2
07��@랛�p�e��5�j�.��ܔ^��(H̶��bK��2@����Rqv0��Q��M�����
p��
����xճ�9��7��gp48�F�Ɣ��Aj��U�xN�8;l�x�i����Ekt瀤8��!ך�^1w���D�f��A�2��-�$R-^\�2`pj���jd�,����m�Ov�����`��5k��X�u��B�3�9�Vq�3���I�h���&�7�� �yM��^����Xu)�l<���ȣ'�ܼaR$y�)q�u���rK,�j6d`
(}e�|�P?s̅0psq��b�����\-_w����a;�RCֹ�3�ʴL�n�?`�XYSxDh�dƐtHhü�����3q�T�G�l�h��?�v<<3Ic�]x��ļo��d,�¿�S3�W,7�g�Aa=�T��0 J9�d;f�z����.G��AB=u���!P��:��ed[��'�mM=��&ϐ[Xyw�`�Zt�pu����i��B����J�}�c�ڙ=�b��|�F���U�x]@p+KV6b����*hM|t�����B��ӭc^}�P���ktEd�Tʢ	�T�˅�(|��V9�j���c����~;��_�0a���{|r��YAM��7c�y���u�f�!��y�P�t=a�s��Qe��Bw8�b����"�
A{� ~�=��i7/�c��I��X��X6�Tኊ�Qe�fk��9�6�3��ÿG�k�����T�X܃&��  �C�
�#4��]n��q������j7T<>�X�z�3�iӬ��X�3.���uK�Nw�A��2W��Zf�O�Ȏ�Ll ꭎ5M��sZ����e�����<���z�N �?Yu��6E�b�j�|p��	1)#t�6�~1�8�D�D|�b�( Y�$d��`��T�y����WT��J6^���o��#M2���ڇ���,� ����;�z�c��!Q�Ae���?QK,���a$9#���̓V6��줺6R��&�Z[q��
���V���V\Ӗ��љ%UeR��扷$��KZ�On�/w/:�]�	?������g��*!�0�?Z_����1��4#z!�&Q�ӅZo����e��,�lMý�\o:�V�Sf�/����`$܎s�7G��1�fr��.=K��<R"�;�@�	���ו��G�,�M�O溍c�N�g�y���l�C�|�"<��PM^#�KC��V@h>�M�bZ��ݠ�V.�	Z?�4ֆ��0/8���;Q��1z�67��9�=�3���tN��A�2`�~ħ̢�0�Rv�F��&���A�T��S_�^�^��i� �o��d�Ʋ|��#���
�B�n�g\���)3�DѡX;���T����mz+ H�+�bL	ׅ`��}�����IH$��
{%��� ���Ę�`�6���PFS���	{���u�%w�	F���g5��&�NN���]�8������.��L	�p��z�=\H� �sf%�<6]�y?_O�B C�����]��cg� Xnlq|���$n��}E��/�줬|���{���/i��K��Ēߨ�3���13Ɍ��,��(��,D(���=?5��� �qH��=�,Yj/��%�Z��C�6D�3T�	k�bht��u���1��Dy���\0��irJ{+Ls�)Y,D�g`�>�������6���8a���~��8~�ŭ��z�.)��%��
��^�Vă*d�U��u�j��yT��N�1aF>�A�]P�|@�?"Rw�V��J��#�~�����hQ����?�P�~�;Rȕ4>��א�7���N �\j��]Ӟ�<�y.��g�f�Y8gg�}��
�����N�P����{����]j0޵�]4��ؤ��h��x��Q^BHUN��9�e���X��q�~���jսP��o�
A7��K����L��䒶>�ڙo	8��X�dŖ��q!+���$�֊khH#`���/�|]�a'6G��@q��{�zD���mL�3�����|���F��)�r��ck�a�vk�W���.�1�O�%��?��$�LB"��M�'��2:����$���q���x�u�j*���}�#V�ڍ�K�VY
��tr����V�-`�s�I�I����ŧ�`m���:���i�o9�7��4r����+t7T
Z?���0��-;��iș#&Ha�SX���t��PQC��&�y�ڤ5CR�}{�e"��H����B�e�aƭp^��NO{�s������ӓ]�������X��]>$�g���� ��C������,��;Ř���i_[l;�s��d&��6"�ߒ�&St�)����O�U��T����C�\���?f.{$ɗ�M��y�5��><܈<~m�'�(\�[~K��h��?�m�:���� �qz�E�
*qG���W�K��� 6B��� �����L�b�(��`�)����y��+���f�ml�0(��x�	W��:yY�##�o�1NAk�5MQQ?��h$Ec�Xp��}���p܆�����uq��f��L���y�f�1���Cw�=Y |K��XP�``��E/�L���,��Y�u�U�z����q'�7�-u{�"����]h\r�4$g�+���8�><�5̔���Ronm9[3��[^��j��/F!P�&W��n�[�?<�l���3,,�c�K���^`�7#p���#��M��kP�}���Z$�
�$�L��c#�����t�	�=��Ijq]�ˊx3�Ƴ��=�(dc�������Q�8����P��L l�pKY�k�pN��*̀lb%����>{Ч%�n���L1����}�_Bz
6ǤsR+�u��ײ�F \��Y� ����[5tv�sV��(�,��R����u�%��:qT�i+�U0���|�1�������Q@��𹣢0�AM�sS}�ʨ������ #zk�G�y��DX���8��ڨ��y>QEm�0�E|�&���x�ܼ��cu
}� T�a)�c�Q[��%$����I�Y�>�����}��-��R�huh���cM�I]M`d1����Ou��4���|����Cw~�6���Ա/��:�H�k�A�C�H^���u����b	�T��L�kX�8~X��=$�m���/�V��@+��;�)>	u�ԥ�n>x�ZZ���ZZU�&� �����33ն=��	�gi�B�	U6���?4�ر� �^��?�n�O��|��7�l�0@��2B��/����n+��d'mh�;{2��z -j���� �yj�'�]��^���:��tk��YQ���C�ך�
����=�[b�;x���U��,���D�^]�
��z�.�"o�<D�A�0��Q�L�vx��R(����k�K+PT6\Ds���B��J���~oz3�?�_�_��гST|>I�{ fv�V�IcQ�� l�߶��J��{����M�~�jZD[_�~8���@����R�Q�߶�P���I-��W	����� �q���;�k9�(��\G'��3�W~����>�s���ԺD�GL�YJ�?��0Lͩ8-Jmd=�ܛ���ڲ���[Y���O�o2�c��W�K����k�{�C!=�{B�3d?�0�	��?[aʹ�e;���t�����I����+��a7�Z�Ȧ�YW!�o\_J��i]��H(iڃ�9`ȊQuPቜe�s�E�Íb��XUv��9��萬c�頾��I>{�6���_�����pU��Y�E
U�;�10u��H��8��ÞUj�B������,Y�0=S��SE�'���ƅ�����9#ᗇ�t�x�8&-��1`p�$���"��yE�+�����*jl���LF�O ���]��ϒ.��\��~N���X1��"��GzMm�%�7�#�n����(v�'��<&�i�O��)0�^}_Ȝ���K����\*v��������#���y��]3d�	*�&_/޼�W0)9���lM���V�D�U�h�	���MA�c� 7����RY����K�D$��M\81�tEB���:,� ���3�GA�5�%#�^�-}
���J�%� ���l_z�l'_\��.Z�4y�����\[f?&��N����Q�B��J�b���B�I�����#3ԣ�!x;l�cMws��xz��p����"�.[!��P��!@��I���4�� �e�Q�o��ե��������A�p�Z�w����ǒ�&+ڑ�0��Z|��!�[-�l9����39�e�,.�Y��Hs].e>m�$���@�2<w�pIukd
�h�/3�;GSVH�� ��tS_�ߛ��5����zq��d��R2�R�����[�0�C_�ow�c��R���N����Ρ:5��-�z�Ho��am)-�,ɋå�V��8����d:�����r��S]�:R}(�k��Tm��u)P���h��X�����U�+<��B0ܤ��`����q���D�xC�r���/�A��&��in���&���9rJG�]r�)��rK
�\��9�0Z��������5CK[�0��D:@�l�����Lp ��4	��q��b]���\����H�L�b=�{��{��{��{.D[Z�����̪�7tE����:B��Z5d|��l,%�v�+#-�xT�bǈz�o�x:ۧW��������u❵��+�$4��S�w�X�vN�@��ǉp���`�-`_D� %q!�<)j98-��s��N77=���5����+���_�i�Z<�����?J'�a��$r�T@f���4]�e��H����t�0xp������^������Z����7i�h�{q��z�ŉ\=呟�5H� ��݂ѱ�'���V�+��1��fݵ��9�N��^��Ix��Ş��VZ�2�������7-�%��������(��JA'	�t3;[LAaB,(�lH�c�e��7р:b��qZ˘�G�Mh�s�D\�����cx�����J`�g��g�5�y`�%1��7�Zc�颽1��U�e�#k��a�N\�6�*�`X�G~�� ����N���f|�q6�[��F� �6a`aʝa���/{頕W�"m���b�E!�A�ݢe��(X&g�1V�A�oT����=�Qm�!~�q�|�C�9��	��޿�N������a79xTB4Od�<߬�>��@.�'�Bcv�1(}�#���-x�-�t�Cm(�y�ܴ��#�����L.��
�y6�1��[����34'���M����؝���[�=����kl���#F׆�$+��E�K�F�YcD���Ĵ�{�s��� #�,��d��6�C��6��Q6`}�J��،�+bH%�=�=ˮ��0�  ��u��OJ�����v����m�ࣖ�ZE���o"��G���3�푪|�٨�?_W��]�X
�7�(��1�r��z�yS��p���⽭|8�\,�Ԗˊ��a�����~&�Cq�R��R�;�;鳜���vi�<��
�B�BV���Жk=M���#�ޣ�&��`)KU4#�Õ9��?��o�A.�`\�(�����z�8��� ��\˜9:fϊ��:h���܍2�s���f��O�����%a�AŅ����XQ�{5��YHc �G��~9E���9���-䑡�����Uñ%G��ur�"'��	��6BuyHp��ɠ�qg=O�@���H'�e��K���^` ���P�Ie�#��a�I&ţ�j&L9�@E:�b�E���
�r��p�@��4����GN��j��̋5cK�*��
Ж����VXV,7�N>������;���.F�$��)���Ԯ@.ZՖ���<n0L�8�l��߳��ZD��N���
�K7Jb�f�?u~��UU��vp͝�?�݇!v%P FW���y���IA?�P������D���0����L�*�E������p^*sY�lD>���3I��0��'�-�T�r����g� =��U]*�\��&R�\�|[dnH��Qq�E����t�ס��[�~��W�B��w�*����\�z)�	����"N>b �z��})öK͍,���d�H3�|eJ��6�f�]_s�H�L'B�����"4.��]�ُ7"x�q�lEs��������#���S�b�I��W�7�����b�:E���t�C����1i$��s�~�-��ۯ�%��HJ�u���==�vY�R��`�=���~|\
�����L.�*�7���@<�AX�ˮ�̞7����Y��:a��`�A�kʃyp�����6Լ�������Mo�������-k��w_yk;P��Q���'�k���oS���z߉%9%{. ΋Ó[|�"oҮ��RiE�y�pȅ1�v�]a�g�A��O�Y��Q߰���/��܈��0ǠT.G?�mۉ��>�W�������8���G�JT^���24�"	���}
 Ȇ��<��#^�Vط�~'��11聣�D�n$R�û��M{�H��R�B��	��JZ�����:d��;9���-�*��xwa�|��rԔ~Ѫf�&�^���Y���J���~l�Es�<O�F�ȾTFa���^ZA��au��;��V�H��o�j3C|U's�:3?�>�@ ��˰ít_��%��g^7�i���N��ƬG�G)踘��xM1N4\3jk��m��f��K&�ݼ����B����$����������V7�#D�+2JL�MH��� ��܄����N���D��L<�+��T���m
��p�)uQ��5�Ue��q�ύְ�҉�d�l�9N��-�6�7C&�^\����j�b��V���s�)���)3ڕy�|b�z����z��M%a� ��ʉ8wDY��a����(G!P��&$&O�X��y`��C��ոBOt��F�����~���2q���ϻ���9��Oh|���c[�M�{h�*0INz�Ě5����P�L�q����sB����K�?#�����͢6�f:�o:��W����^(^ܮ�.u��r�kv"?�L[$����EP�W
����Q�.��n�V� $�C��ǹ�ʤ2���O ]��]�rCtW�aB:��E����i@���m(��HL�U4h�
OG^3e4U-I��z���Ñ���VɧAG}d ��B���خ�k.�w&�NQ4�f��O�����d��G�����j=*�"_׍7����hs!�3���0>��=t�����q=��&꒠���ַ������ѵ8R�dݓ�����3hj[�b[h��*����]�9�c�[���5N�j�V�9)��^Er=���͝��%�piq���Px?�m�߼!2m9C��%D��W�������y��T�Ec�Z�眣#�iULR	��aWt������t{O�o�?C�n�"C��ܷ���5�o}q���t��@#]��v�q's2*k�E�t3�����Y�}�b\̹m���~�k�MԴ�5�1W�*{���[���]��c��Ⱥa�M��Z$��}���(�&S���b��'f�� @�y#Ƽ0�� k����V6��E��5�&�I����l����u�xE�"��jt��L9}1�i���u+�.s����G�߶�%;H0F�-�	59s���r0z�>ld�x��p_�msك�.��u���&E  �pn���J-}�^���Ѩ1/;=2�+����í��$��1b��8x��Pd���!��l?�n���;�2b��&�B�ZIL�Z�D雴_�W����w�?�5N����H8x�8M�GS�u�%.�@,���K�.)v�@��Ì�kH� ��T�x2Z�Һ�Ğ�:���H�m׊��>�^:7e��l��u�X����o����ؿ���3�"�b͞���R��"G�����1���$-�;Oֹ㓦���icD
�s�It]r�λ��Oy�˜��@��~�,O>���>�Vf]Ϻ	��{���'�����8��|�{�T��.�����V ����F���l��R]�Ʀ�|��3��@J6i�ͽ6�����s�Z�6Z=7��/�R��x?����^�Y������1Uב4Oԙ�L��R����K��$P���"ij����䏑)��5�4Ч�i���bW�~��#��_+�|����h�}Rc��d���߁�����2�?At.��z�϶<'�`�Z.5�����UF���38*�Z�����e�gE��a�/U�M����PFݕ�D�*�\f��	��H�b7^����-h g�>�7��h��7t���&��=�<��-d\z�I��L�R�� ��ر��?j�;�JG�ccxi+i��<�՞�;Q�Fo�GA3�} +���k��������S7Eg����gI\��pa`�5A:dw�	:��+��pi�%\���]��G|=GU$����a�Y�}��s^I��6�Dw�/>�,�f��Y�
9&�B��۫'�F�&�����^��R)�������L.�	���z���Sn�r���Q��B��u>%=SB����!��#�

^�(���<�X��7�9D�ֹ.�۬�#l���K�0�\>�j��#�$���e�G�{�{�#�I�K&1@�P��epj��E�گ^�g�.l���L��x�w�G.�X)�{\�R��	��&@��5����s�P�/H����_@��zl�Ռ,p�Em`Q�A��x`n�J�R<�6�.-lc�}�E������r���3f[b�k�Wq�K>��9#���{�-�p��dY�}�LĚ�g,}�0�7�D)�:P����iT�.�f"� ����1˱S`!�<����*y1�#_�[el�r#��9�%leP��QjgUX�|>���6 ��2�r񐝻,���q����ABA!�=��T�h .�S����:7C��z{��)�]�����Ł|t�E[�3`2S����_�0�o]��XO��Y���@�l�cC�"�,}��g��3�D�9iJ[Ķ/5�"����|R��f(�n]�\�`i�|1�S27�P����#/�m��8G�t�$5T5X&�M��*��}o��
]���]u�LC��]���W{�q��Ŀ�`�F����@GDl��e�����F'��l��s�����ذmx#*r>S���s�y%�A��=�4���Μ��@�E[Wɭ4\߆��>������&����*|����$���#ʅ�и�W��� �J�;sA\i���ٳEۏ����E�Ѵ�z�ע�?��W84��E��+q������[W:/�SVek>/��g�ɥh%��a� �(0݀�yE�Ce��\'bYD�kįڟ�'�fE4�v|�d���9�橎�z����w�@�ʁ���M��~3Lk�+�u⋵�+�IM�0T�n=��n�c��{/>��E��_0�cXPu�)����=Y�����ڙc:��S�|moX^� *DF&�D��5[�6����)�0��ю���R`Z�yTA� �����J}y��T��:�K��z�z<��9�0E��Q4w��);�s�'�K|\~"��O)�g�1�wI�I{�>%[+㗍8�8e�"�K����p�k�2�)�R�OWp�ٵŠxi��j��`�������{6G�.5�e������3r)T^�9�^�%�⮂&�v��x�<A�9�lQ���DuZ��M0���-=��+֋K����6צ^���DA�D�e:T�_z.�M�S�Ú��� �}࿶P�����6�^%�ms�A$�}y������lZ�Mp�r��ݻ3zu>�S�*���Vlomu�D�V��2j:Ӟ�B{�T)��E|X���v}Uǝ�u�q�Ơ�x'�A���	�j�z`���Gg��;{� Խ<�d�'�{D_F��^3r���� �E�s��(X�$Æ*Sә_O�4D ��P��`�{�p�3\c��P�t���`WGQT=+,4:%��$$��}M��Z5Th_����@��&&��7w��j}��Z/t���$r��$Ql���| ���ɾ��|��do�*�Yt�.΂,�?q[(�ݠU�=ѮG�)I�����۳l��X����w��^e``�����߱X��M�-1P�/�ʣ�4��y��߯>��3n;+#�F*sK�?��׼���9���
���ɧ�D&�b��B�}�;e5�wll���0��#�Q�{(����}�xj�
c��}����j�]#H-Y���*R���H�Li1lT������ե��r��0{�75��_x@�aR�cN_�����	�NG�F/e��gq틴��fI~);J��6�uwꂯ�,6��y
e��9���6f�)��
zM��&l��S)��ѐKW����<�b���3>����T���L�&�ŴG=�Y;^�~d�M�WU�p6iT�2C���9UuͩZ�u��xJ|*v�g����X�N���r�������J4y��h�k��'%�D�1��%ﯲ��ʊ�;�o�tk.=���dw��T��x���I�e;�i�^��<2)qo_����D��W����%�����" ��D�����%a�7��q��)�i�iV��ݔMǆ�b=�_����
�/R#GQy[l�$��A�g�X{Q� ���.ӎ��^Y�/�a�����@����`b���<GR�D-�
�1�+���E�5N� �+����:�g&Y7�/�+Z��t���Zn�7˂�����L���~���L��l!�����tN�+[T�J|��d &᫴6���V���Oh|
<�`�[yag�ԁ��X�"�w�X��9X�\Y������/�*Y�ε뿑��~�9Bm�]�a�b?��S~�@���,��xv ��_���͌��l��5m����Xw0����)�'��':���ݖ�shl���\|��Q�ʹ�z�pË����Ղ�Ctш��L#-���|l�:�ӹ����;%���i~+A�x۷�=��������Џ�)+�,��{
�W hV�I�JiX_�a8�Aޫ�};DZ��YK��T%�Ր�#8�P�n�ݗ[y�^&�Ջ�68��J����@Q	V�Ev��#Y|�%��(��g )|'|����ׄ�[�X��1�"��*�9������c�N�cէ<cMP&�h�$��3/��y��|܍`B����������
� �����,偕��j�
sE���e7�X�w�*��Բ]��4W+���g�NG(��7̥��=��ģ4J�Z�������u�ܣ��-��������t%y;����ez��d��;C� �@�,��w��~%_���R��#({�^W��7R5N�"�@�5�zD�G�uRp����ȕl�R�\ԣ���������-��j����,{N���>����N�b͔4'�N����v���o�����#M��^�-"�!�����e��[gcT^D�
+��Ե�"��+������8#E��3Ĭ�alp��A��(��s'�:�v+wvf�
6W�4�&@�y�N�00�����n �Y֏$�](�o���܎�E�'�+��,2%�D�Y�p�����?`��2���~��r�@Ï�K�����Ġ���z��u�(��,�a�/b��{��+��3ܗ�]�o� �v,8���ZRE�����v�2�����<`S�\g���l[��}"_�ƣ%�Z��� �-�'�DXQ��9�e�X�v�ԒpD��3�j���-4�ׇN^)�A�a_����������B,)��~�e;w�v�6i�pF�qn��C�S��=l��$�(�02%�\Gm�DC������IdA#�l�G����U8�z���$8���x���N���s����Sp�����5{��q;���,��%��l*jmU�`@f�F� �o[���L6�?�2�F�dF����<����l�UW���B��x�Z���qG�vв{t�{t���jo�7����������E�7��Q�m^p-_U��s��pHr��Е�(�!��{�N.�%�h����\��@N��BU�"o�AW�;��\����WhA�*����,��H%��8�� �ZGHi.l-�K�`<����t��$�e�r�t�:M��{��¢��M�r�����ݾ��`�I�鈤�Q�u]\D-���QA;�0L�7K�y%���
�|F��	������,�Ƴ� ��?�BOm�@��fqגsݻLG�@��sW���<YU6�� ϴ�Kt� bƝm��7�"*Z�i�z�4���U�iB��,��R���?��㻔�i@��B�u�&��h����,X��ৠ����#+�c�Y�}��ﮥ��-�30��P�nu�GF���(��FT�Ƃ�O,hsz�&����m(ф��^c�e��9(>h��I���[���E����G��W��;���މX|���U)��i���I��ɒ�T���&���|�H��u�C8�H{�4�M�~Yp�T�m�E�z�@Hu>Y��#���W��s���9��b�	VG��g�L��j=��$��h���'{U�
y�h�1;E��Axt�3��?z8!���Z�(h͟؛��'���'�ɚ��J��ߎ���F��+��"q~�3`�<�Yw��;;��R�P5�D��7�}rt��/�=^D�+Lp
���	��Es�6l���I�ܠXjFF7J�r�"DR�.$J���A"��XM��IF���JY��	-;#16�`�*�:b�<o���'�*Ey��6'���M���p=�[ah,�b>IA�F�U	F��Yy�hh"*CM�]0���M/O��{��������Z�鬀�?L��XJ��4ⱌ�>���?�C䙧~��SYl8=�Q��81)�%m�\������5^A��yJ[� �3� Gg!��&ˈ
>�V'��ya�hׂa:,"Vm�S����@�J�xw��G���S��ف���+��TAM*�~����r�:�W���Fz9���=�lkp�E	]���W/8�[�Qk8�Z� ��{������{s@Y�5XAm��B�F^!�;l��"zYQ(�_rX\�հՖAK$*������[0[��R�[.��Ĩ��()uV���>[:MsP'�I#���xԉ��	
^������g�x�G�+-x��Tu:)wK�tű��X^1�E�&��֭��[8��oͻE6�گ@O���J�&8}��L�XǓ�hW�H��.�F��M�5��ol�\����FA�|�;-���&+Dվ���befw]�9߰���3!Vn,N���J��L�^/�FYs��1�A�)���޵�ۮ��V2f���A'B�C�w�&n�:�V���	u��� ������"N�Y`����
��n�F��ld���Dt(�,�޶��9��ߠC�ڱQת�c�A��]l~���~��}�_��
P3�-&�H�oJa�R *��9m��N��f�Ai�T���� ��%��)`. p�t�j��YA�d��?ԡ��5n��ɂ�w
:�]�"n,
�^'�N��:��M71�K�*��� F��1f4	���xڋ�_S(
5�&���sʇ�`
-�6���w����,�{^ǎ� ߓ��G7�軵��v���z:�ڀ�(z�w۸��#�8�	5���J���Ct��?���>��	��]s֬��{�f�x��ZT}K���Ի���^ޠ��¦����DH[i$qꦯ�,���nh?얀k��W�*��d�D>&���PT_5�D�Zo�)l.�g=��W��04Հd��q7%���(��������o��9\/*=��� d�Q7��Z.5à�*����#�K�n@|�z(|vgd����Tz�r��I���C��FP b�5!����(ҧű�H#��7Q�9��p�b��R�  �~A�6�d��Ʉ`L+�-����R�K�y���L:(s$��ɛbzGp�[bh*i���I�2S�IE��Y?l:nU��;�[��+�卬<�a[	��-��1��9U�p<�'��<���b{��ω���6"i��u���u�W� g���b=\��&�A&0x:�_��å�Z�c�8����c��=eE�__@�,E���9��;-�٢�׊wg��� �LugT�eD��d���͢��2a�D`��|jc+��3��R�� BF t�Ӱ9{�+���~*�޷�B�x��Y���I�X�ry����
���(z��Yȫ{ö�ݞ�U�y��\�b���d7D@�$� ��ߢ����>+���B��,��2K������t�u�"a�����h�v�m;_,�qi��߼�~Y�L�	������p�/yܒ_�k3�d�&>u>J�dyF-JN!����M�d�[& .��W?%���=�"���#9p5�G�SƟ�����u��3� )#��ݽʃ[A�^�g�ڒ(Y�T���������D��tȅ鈛iӏ�s�4���M[r�ƀ�z�ؿs	-��ކglx�G�X�m��˜8a)�O�o�[���SO�';��M=�͙w-h�	pF�����'��Z���V�-�B�$����>ڎ���^�E�8�G�����/��Sb�2��ٮ��,sׅ�����:*�Li��9)��a����_��b��S5�������Fo<b�^��h4B%�	[��]���5��F�Y�=���XQ����TA��<�nצ}����e饒�<��?�śM?з ��DٿYO���2$��&�^�^�i�a�VML.���)�ǮR�e�ǔ�����`����m��I��dW���U5�U\� q��	/��j�v�>�Yd�t�\z�슯a��:jm�mG���eKdɦ���|��x�j�mW���v��s���@S��Hr}�F{���(Smy뻺�H�����BwC��9�������ܬ��/i��ëY�H�{24qw� ?Q�Bu�z��ܽ'5s�6�\�x�s�mg�s�k�}_d���mr���ema�f]`*��.*��t;�iw�"-Y}$R��O0�@�j�9BS~.*�u�b�Bo/]՚�ƺl�-8Rn
5�l���%Z���֨H!�4i��o�� �t�YA�1@g��`�n��#Ycl��~M��Ie��.(�����ӐE��yJz����1��h�I���۲ҟ$<��<��%xM�_˛~��O�~witn�uE5M����W�0 ���Dt����$�%�[�+q��H��2��tB�a�8m2#��P����Zs��M���J��-9���^cx2��Z�lb|�i%f5�F^���E��%*'ٜ��;6~�h�|���(�#6�8],sR�{c�����ժ���b�k�#�]eN�}���d���l��u��G0ik<�u<}R��7G���o�ī����(2!�ʈo~�@&�	0�xC��V�[�l�zV�� Ƀ٨9�w7�> i�I��*�a�Z�ī�o ����(�˘���`��"���`Ec��
���m.�F��NL� ��w�|�o�/��E5a�>P��X>9��̎��h���XM�j҂ #~�$�/��Iu}:�%��k��zm ����*A�E�Mq�+��y��JMN����oq5 ]�\V�j*��0#��u˝�z��*�Z�9��[�[�����w�ϵ�6����J�1�.(;m�o�[�m��^�^(�Ȱ�C'�����s�z��g8+:�"���(Bmy������E /E��)ŭKy�3�R�^M^���MB �� �e������=$r�l��d*T����P�G�˯���ع���yh�tf����8*l;�Lwހ���	W �T3�`|��n�m���{C�Ù�Y��8]���ڌ�����/u�����b�q��;�f��؅�7���۪��W5*��	�#�9�=���E�
k�?8���^�f��f��w�Ihd"T�\��L��4
[��#"צ	�5��44�)q��|�	���n핥A�w�t�����>'�]zx?>MX���F��83���nx�G�?�Y�S�Ab���N�h���Dݧ�N#%�	��Q����~�dn����0Ao~|]JO/Hl�~�\E��*��ǷM}8ƐiǱ4��%QϜ%˖V��ӗo��o6��ZXJ9<|nu���
Jc�4�z�^�9�:��(�[T���i* bL�+�#ݬ�p]���\x���<�Ham���w#��?��A�����BC|��r=Z��[lª�Ɉ��2|���#�9�d�'=[[e���^k.�D(�xH�[[�6�xH�<���W!(���&Ax\
+�<d�bO����������c���d�Q\���ɛ�L)�h �KQ�V�%�9C�ėF�������d��E���ob#���vuV88���
��m�U�Lq���[I�����ǹ�0��E4���U�U�3YS�V?f�����]��Z����.I�7E�fS��kAǟ<�7�'10�MԚV��E��/�dW��vx�u��_M�ܱ� 0x�iq�x���p{52N¡5Pm\��H{��A�:�u\����������
���b��8���YxM���q��]E�<|f�e�BP����O�F��b��lJ���� ��ХQ�yX;Ѧ�l+��":��c!# ���IZxM���-��w׊��M�[����2b��|2׶� d�;}!S��	���ށ0�NT�L[��@. ��+ᅇ����� �	갯�|�bm����<���b���.2ӄ�*���S�:MJep�Ʒ�zF�PwchK�8�Xl}J��?��Nʗ�gWV�m��2�8�|\����b]k���,9�T�%�j��j���2���uL������N��~�m����d)�1��%4$�x≳�R-5hw�a�ql wc��4fKi3��@�����CE��5��;��b�,~;T��!��L������"����h�aE���T�	S�"_c��D+t����\5  ���R5U@|��T6a�b�6�|B /V�0�����8����꩹Sr�2lwZ�ekh3�|9�����
�x:
�.��g��t���A�B��V���F��l��Z�d�+>�lv<�CC�1�]��̲�^��Q��Q�� -C�*��	�F�m�u:���l@�j���q��5�z��L�O��+�T��'�`���˟�S���\���NB-ǼTJ�u�¾�l�X�4�Y!��ӻ뚒�=}����y}~[��A6��߸s�+��-��*��gU{��U�9�ʻ��آx�������t�z��	FvKNQ��^�����í|H��W�O�A���IrL=���Ԕܣ�޾�H��K Ḙ̇���PI�">\�V�����E�{�<��H^����Ľ�\�?1١��Ќ�j�mDXW=��CUԆ�ۂB�=ǃ�ֹ��%vf�Ģ݇��wx�� ;x�3���X@+�>�R����W��p�w��f�(7@�j������[�FT�/6a-�S'��m����!{�ʢ�ǿ�-,r�����ө�dn�u��tW�W/��ԟ�Bj��/�4�)�jAu��w�^fϳ�Y^A*�K����Wy�oslгW�S!��U=�ԉ����i��.̧l���v�d���+~:6bd;��[ڕ��i}������ts7Q;�g괁 �U��8=(U�v{�}��|[�u���>�M��t4��Sg:�¡L��Ҽߙ�oi7d�����F^A��ci2Q0e���v����,pja�zXh�Yev��YJu�11a��C=]ʰ*��h �ѻ��L5ȩ�F6�Ӛ��n�Ӄ){Z1��s����Y��\x-�'��!�y+O�y�������$:$Fm���o�3B�9���0�'E|�m�zH�����f:��G^�N��i���Qg]�3����h���C� *�nBG��K'n�F%����b�9��s�6|u7����>�#^sDI�Z��Y���t@�\�@�n���	XjK�ұ0�d��6z���ך�����ƚ_Y�t�-B����i�$ ~��{Έ���ݞΎ�# �I0�������[f�c>!:$�����Q	xJf���֝?������NT�H�i��TE�N,/LO�А��QRv�^�׏��!��*�T*#h�~�C��dVE���htk���/m�a*380� r����#���_��GS��ZKLj^�|A��7ߪ
�1����8�Ї7�RR1�ŃŐ�H����ؙ���Ir0c+8�F/`0Sӷ�J�Y=N��SV���C{����}#Z�������ș]w��v)jq:=�>�[@q��N�ݎFϚg�O�z�A��� �E�mGR��̳�����'�\��?����������y�\CD~_h��pI�QB��)���q#�ÅB��&�]���cz֨3,�Ӑ.^�KUP�d��P���.���!��;T�\��,5�;e��2#x���M��$k8�0�ޥaՓQ��\�5EJ�1��g3q,���w{�x�3b%���D�9h�9ԟ���x7y摸F��Ȋ��޶%;��/������cU��1n5�cs��!�V$r���8��	���u�u�F����,j\o��s� ��Kv{�,5�,��s�H�z��ٿ�&���e�kI�[/��Ke��HO�i�7��C���G�.6��\�jј���Lv.���q����M_�,���4����O7�U(!���J�z�|s֔᥵HHph�bת�{����U'��d�٤Ti��w Cw�����Z��,�uKb/�J��K�΢'�SĝD��"����c�� t4^�QI;b�j3�B餻4̱L������zC�Y�r�*2�<�Q5Ź C�?J��n��$���c溤T�N>jw���@Y��QC�����M�U�8�r" ��J��<�e��Nq�@d*v������!� ��j+�Ƣ�#VA9�� �~R��v��ǀ;R�4�%H�p?��o2��e� �y���F��7\~��䆏���3��Q��=��Ο!�d����S����\�`�ՇRa����a�!��-�ҧhKCF���CD����=�������ў3dֿx?�cz欒G	����n�7�UO�V@�;�S\1:�P��O��-;d���lW�1 c���̦ޘ1!E�4eY?w���R���!�8|�DO��,�W޿i{^���M��g�!����r�D06r���>�:�b�t,�*�s~tg���
F63�*�0��2s��2��g�Q0ѭ��w,�Sh���d!�s_��?��'�2�g˸�g_
v\�v��V�����~�
ז,_�FcD�,���R9};h����BA�H��L�{+�=�ki3����t���+�[���fC~�����ݳ������Q;\���JO���C|x�=�����%�e����~τ��A�	��gVc�����h�:*��L�Ϲ�띌�0�W)��:��N���wb�.It37	&����/�ۏ�P���6)D7a��m�f-E1�./�I}��W�h����EO�����N�k%9Z�J�\$��t�F7��E'܋3���&y��%�@1~��� q�ߖ���d�Ԡ(hV� �!Kt�`1��ĵ�w7�g�a!�Ԣ�,ci$P@����wpB3�d���%�,9��yK�7!��8Aȉ���<v��n[�*��,�lnz|O�.���䚹�o ?�zs����:��q�D)Rp����c&�<�<��!s�/H�Ϻ�2�(��҄�h�Y�}'��`g6{Џ�`��@\�6�ď��i.�X�皬s��t�>^H�[
Ч��x���F�|L�����K���]�q�L�ܬ�Y8�E����j��P������P�v�)E\��RB�W�أ���t��w�����/���U�Hdx�Ӛ�?<�G6{�=d�Z��c���u��H�*�?w�N�t�c���r��E���3��H��W�Md�
�
�[R�U�Z_�`��W�#�N�ш����"�Ú�;�p6�V�\u��H��EΤZ%��'����(���vw�ƿ���p����᪓�5�h֔Oۈ9/va"=P�diVJ�����<nE,�#��:lqê܄�0�$��llq1Ǿxu�7�cQ�^���n�`�����unC���oFnC;,�7F��۳��ePB
FQ�*l����v夊x�|/Ǘ�Х:��*�,Jt�zD��ژ?�R$؉�Fe�A@��li�bOf&�=��>]�zy`i5�~�B���BΕ1L}1;�ܚe�
N��fw��p�u��?��ܡ����^;Eo /��K�Lt0�}=Q����Y9V	�@�����O9/�T��9�����؇eY }��R���	�x���bʇɨ���|[゗��iA=�"�%��������x]eG!�E�Ӹ`<�|���[���<��E�U=�!��(���U_a8HrA�c�y{W�X=F;��� lhd�Gj�wyZ�	��3~��׽4�\r�>�HI5�?,2d�窬-�N �c$:h=��gVt�}="9P��V��ҫ�>�Vq	�HCC9Hs`��8 ����z�2�`��]��{t9YC���ZS�W�j:�F�~��!��R=1���Xb@a�+�2��H���߆����'7H�C��{�ap丩S�����2g~�v!U�sE�N�_Q[�fk�<�hyOV<�sp��Ϫl~:�tW����19����.	��9��^�)��I��9@�ψ2��e�g�������ʥe�;!O���xiHH=G�C�g���1����n��s�yٟ�\���fR.d�FL]��{ӕX�v#-8�RX<�ԅh�N��2��ϐ*e�Ĩ2�Z��!��F\_��bMD��=A��d���'��oY�0�N��Z�^T��.}���R6-:��q��E-3�s�T���ȱ��r�J��neU���c�����E��.��=������ܫ1k7z�Hg:���J�#�Q<�����i���"�&2�`E�^a��2�r@�!�E�&�����Z�f��@����*V�	��s��8S8�C]a�����?ܳԀqU���إ������R�h[��nvN��'���Ʒ���v5�قMf��NJ)��5Q]�_w_l�Ҧ���?y!� YQ�<����*h��eX��ꏷi���);�d��s�J�G2�\��:�k������5+{��+��Sp4ӪZB�Ap�/���p�4���(�5L
D�ER��ܗ������'��]Y��2>�/��s�j����Γ>;�3��q�b���o�{J��h��C�w
͹���h'���]�##;�a���ޖM�e�H`~~i���VFڏ{��k���I���{�v�'�VZmd-C���y7�5;�M���E�]�:�����۲tr��ȂQ Da�Tn	�Ҿ���  �w)���7�X�h��*�xrl�L�ܟi�M��ՙ��ky����\U�y^����"�ӪЍ��c�J+�3������e���)��[G2SǠywí�;��:KwcE�e@�7�5XȂ�0���%��eN�<��t;?->�+�r�_;���F�U4s�f���QCmÈyf��12�W�&?�Z����ƐҽC�y�B��:���/��m�T�G#U���NƼ9�(��f�����)�>������&Q�X��v\Z��T1����{*��Nݤ�'�b����CL#���zIx��%��xsP%��Ҍ����$���h����Ϟss�v��5L`�yzk�W�uw%�G�����3�f���A��8�ؔH��(]�5a5�7̵]�똧U���
?�2������%����;�NS���r�1�ࢩB�b�PQ���~d ���0T\&���#�����u�w6�lˬ�X�8��]�%��#Š<*�#D�)��L�x*2�Et~���TF�Y���)��Cl�Ⱦ�ˇԏ�鲭�;<}� �J�P����~"�(�&�8tx.��ٲn�w���'Աr ��\���j����>�(1��7���2D���n*
���H=�z�\��D�#�������s6^���Wʫa�ӓi�A��Gd�sZk�)����L��fO��͢*1r!�_�0�N�TF��0�y7�Q�ck%�k���Z��GzB��C�w����6�"\�ݫ}e;���)x�I��nE�ADx#T�ods���@3T̿p�K���!KȠ`:������*�uv-`K*+�܈��SN~h���@�AF2��V��� U��"�?=�&W�9>wŸΣ0/�o7s��w�+rg�7;���O�����3zMмye�4�q �'�zbLm,s2
����0� rD[1��
�뛕���. ;�2����I��)C�1�u���(s����C�(%X��$�|O���]BBE��* @������`:9cB"�`B��� ��v�1���೜��yˑ]���t�%�Z�1or��j�N�<T��.mi2,���+�l�vV��,����}^@��鏉l�^���P�9"�,E�0���:�ldR����n��f�'g -�T��)P��8�opY�Vh���4o3�C�c�8���Jf�~�� �<=����"l-�EM���͔�/��7ȞtjgG��O�Z)?DD���ߊ�	������>��`{A�s �Uw(��k���L��$r��t&f��="y�X�k��R��N�D��k��ͪpZ�,�;��"&��E�T���>�L���l����f�Z�i����w��a^d�S���/qj�Զ#�Q�0���W>$��x���4�dbn�F �;�7���������Z%m�J�or�ဪef��Jc�������nrEa�$&k���k˴/��g/8@jR$���C'�S��"xJ�yS�Q=GUE�|�ۜf�0w�" ��k�x�Mc��ܚUb�u�V>�R��d�d;?[
6>~�ܧ�'w�
r@�
�"|�դ�5�a�;+!z�֝f�2�9�����0�{oo��g����l�u����!N�J��[����<(�LR�'��r���-t"�AJ�c%�[��X[r6�D��,p��)�o�����N@\��Aܺ6;V��sA[>�:� �[�F�j\;�d4+���i�N�m��A"]j�I�<1 ������#nNw�'��]�u>D�ۛ�i���_1�#7�]�k�q��O�I�"S�6�PA����h����4�w�Z6c4JL̍Z�zO�FP�m1�6�T6���o9]<@���Nj�,�&+��s�6��f�Є0I���6l�:P����/���m�����c�}zc�T#���-h/�_iz���WJ(ؘ�D2l��Boz����կa-��«���WLʚ�����U̜��\(F��y�h�08=Nb��H�>1�z����P�'1�i��"�TU�:g�k����Q���a�eu�<%���ht�����#SX �x7ˮ��)���"O�(�<cV��
��������``���Cph�.Ƀ��K��ھ	�Xw����U�`wT=w�д���~�¶OPr��B1�'�k��������/ȖK�)�����:4�9�t�����~!��-��}����]�Q'^�-�ay�|\O��Z�S�܂.w
�[Dʀ忴�KwC���Td��(��V��ަ��A@��݀�1Ke�@��f��D��4����һt���a���k�c	�v�*��av:���+��0�+Yi�Re�*�P�LKJ�+��߿�.��S@��'g��IFUZ���-��o��*Q.V8��YR�r��D�1���x.���7���ƧpĞ|����q�?��u��O�
�i.`��{T��h�ؐ�~���M�O̧��`f��h�~�I��^Ve�<�в�P�1i�v�m�!��?~V��f�W�"����
V9�y�p畫���}Em1���pWn��8��߉����)8ٽ��qQ��i2.�5�p��L��S���٧7�(��8��Mԛ�Y��>����9](oŜ�u5{`��K�HG�Ѿ���׉����qڤ+�E~/�"A6��*K������c��z��O|�7�:(X�H�O����f���>Gg),��v�k!:��a�+UJ�t��J���L�͟u�=p{�yw���;Q} �{U�������is�ܟ������)�Ա�t��2��6GHd�,��:��,�����w��De39�/80�����AB��O�QOP���di�EoU������oq��Iu�d�U;��	�t�½��8e�Կ���$8%����ۯ1B�[fS���̕��'<�[����F?7�2�v��R>V?�l�;:-�@$���iߐ�� �������B�����G�BƲ��J�S�z�?�igN c+E$��:�����vh�x�;�Ri7�k���Sx�z��Tv rEW�A�{U�^�ބ�p�h�}��N��m�I��HQ땹��?�%ĝ�˒�s�&o5���r��qD�����^m�c�݀0+�xB�U�ԤD�5��n�5��Ɉ�~j�~��> dD�����/R�h��+n6��_O<�?��7D72�[�-B3����{��,`=#�-���;-�7��̔��XI	:�J�`��_�wr�7��ymJK�%�e�$U3���I��59��A���7���ݣqe�t�G�Ҩ�Tk���s֜�M�1��F/���Q�79n,�-Nq���:r�AO�$4����R�V�Iy���ּh�$�)�P ����1B�]����Ë=�� ?;��g�����.3��!�PY���5����G��s�o�:iE�~�
W�F�ս�h���n����^��f�С�܆��x��ƺրܑt�tP	�l���r��?��m�0�� #�Ϯu�u�Y\���0������J���XJk��i�z��GP���1o�-����K��K:M��I^v��N��,�*T��}=~���<�l� �Kt��)���˖�p�����y4��:��Jsvu��K��-�-��o�f.�	N�l�!�OBQ���6�b�3\>�ObщK�R�4���0������TΝpv�,�d�{b$�h��m�8��-A���5f�{�Hq��=�Q�(֙A���H�@�����QO����#���,X���z�nA����Տm�M6f&d��(����\��z��.������W�;D�=��{��y�<8��\q#{�m:���~�k�$�P��0Q�����uaሉ��+�G=�&ƒ< 1<'� QE WK�A$ѯ���Qő��9o�Ǔ8y��ۅoē�/��\���x^l����o�#_%b�Ć3��Vy�4	[}X3�c���3t���C0g�\<���ߩ9	&������!��g����h>��uvs���-��PZ�����N��S���`�!ޱFV�o4A���I�>�W>�[*<�^Qg�6�����d_�r�$�Ռ��`�f�lƋ���2(Ӈ�������z07�/�1�-��gD���[H�������������J{�Pj#:���94��2�'NPTb@ʜX����M�(����q8�����So����^�ᨽ������v��y�~����};��"����l�xs#��l8uX>����o{��'�ηq]�̺L��oћH3JQ�u�Ś�tA�>!JGO�h%�#�Q���M/���4ܷ�=�P��vEn����"mԁu�״sɬ�j lڣ��]N��M�}'2�c��S�>��X�F���-��L���ܓ��xoC�Hre�D�F�� Y�N~cZ���'P�0��7{����jf�3�&��mIC�Ҭ�g��Y�!@O��*��"?$p�bߖ��gd� F��_��b:����j(����v2�>�aT-�@~6�<~�Lt�)q�-o�m��:�=*NȻ��=3,�HW'~[�!�v6D
�h`�g����-��Q��kDu*�O�Zr���:C,+���I�'�x�ʦ۷�*6���h  S�PtcN�$��6%�Vg����Ӈ]-�+�/���f{_8(�WV?�� �\kGAoR��NkQ�)�y��h�h
_W���X��2C��Igo��X�j4�4�?\�l|U\�|��J��Վzj�FѯL�c�y�����X��9��{��L�p��z��}K��-ֱ$������#Q�E5mj 5����xp�FO���ӆ�i�Cfz�3%0�������,��P�k,LU77��R��{�2��c�g5�y�w���TV��m��.�"���>Ft����_y���(��[~0��HAƵ>?��&��da��-Άi���F�CL�f:��`��l_�8�8���z�������;�_(���"i���\����֓�e(4LA���cX�r) 3�dɽ	�s
��" �COĭ�]b>��}�Sb�u��-n�y.
��?-��t�Dy�w�����e}��cނ�/�I� h+y�����7E/��@kW%�7[������s
� �R��@���͚N��$6C�������`�m���v�p����-��X����:��{W(S�c?h��ҝxsܟ"2�(:�R5�����<���dc����z�}I��H"�PS���lF�֕9��X#J�`��j2v�Gz���&�xS�.A�r�V|�M%Vc�:�7�Х��e�l�[�;O�l��Ӣ��hL@�ՋU�R"��8�FR��J��A��U�fmY��M�r�����.e���|X�fW)�6��_�O'ϔ%�Z��7��[�/7���q�*�0��N�:V�jY����ϗ��`0¨�1�@wҸ�� �QB翴�_��\��g�{�yPOVP��$/O|�o��eY�H���ѳ��h'���!b����$pΩ{�$f@���B d7|gu��U��w��b�AY����w ������y���� �4�Bi�[�B�f�k��F
C�0r����7�NqC2(�������6h[���j��ŝ�+��Mp�M��Qȥ��j3o�	s�
l���R�༬rG�Q~�7غ��^<�����|�A����0�5}-@�}�_������������$�"�-�YW*�1�����	����s
f��A��7	��Ϡv���C�Vb�3�����{!Nӗ���2��]��~|��5�ȋfk��A�bw�$�q�0b
`'�ŷ��b�ܚ�x�#m5�qb������Ecv��c����߭�>G/�ɚ���T��oe�_�˱�Wjrm��ԫ&�P<��&\i�]���	�(fyെ�&)�0�N�T��Jzs�5+M�*-��o7�a�DkN�`d���M������E��#��^؄��!+h�y���ݍ	:l#�浌&rӴF��F��7Ȏ;o��4�����J��"K�`I��t�y�q����o�����i;�4�-� �c�#�>�*=&I�F+g������N��+L_�\S����;�W�|ž7�h���E��;N��+��G�-�(���>,n�~^�	b������bR���Ğ4���GT ��rKȱ���oi�EU��
$��(W�q��w�P�|��-7ͪնS,����BX1�VK�d()�q��ڎ��A�{�#�Ѣ��S�E9@L8uz�_Cl�&�E�QjdD�Q��ɮ��x^�8�i�j`���6jī �*�����i�p�,d=�Q	z�/�:ږy?N卯MOY���^ZҬu^B��j����vE/*F� �C;Q�:ak��?u?��r��$!��bXGʻeԶ�~�� +�?r@���	��[v��t�z�՘|�j�����ԹN� A��<�k�;��5
���(��Lt�i��f�)-�I����a�H����=i��"xO1��5t(��\�[�E���b��2�������7�d�������E1{§�M�� w��I�Yt���Y���Yg��G^�%oG}ߤ͕��)fo
j��_ε��$\Q�_�ǂ\�����+�&")�)�̯>o��x��[�Pހჼޡ��{k��k�s+%#�B����2�z��DLz�)�[fk<|$���M�؏�>1����t����G��s}�s�K�]-�li�r������8�?�;���S��o#g���i�y� Od�B kAKBGL67r�Yl�Y/�t�U%1�u�!�� �&3������{�hwk֧�n4Y���y$��,��𷠓����c�'a�����g����cmt�Ht+li���R���{�=���2ـv>}X���A���[�O��i�Yl��mv6�\@f ='��� =���7D[7��\'K�Y2�ċ���f[<釪�� �t�8�$FRs�`^�К���u����X�-�ek1�o�nÎ�����%`�;��j�5}��+��	ȟ�)8^G�qB)M�5�c�\�i4-l���٩ftaO���l�jf<W!n�+�#!v)LJ��J�,�D�f��בֿB�� �_��Iu� �&�Zd@���~�a��(x�h!�(Sx��Mu�����.��g���Υ���Г��,K��57J�ɳ�جv�O�� ��G�
J�`GNҎ�חt��,nI�V���X���Z��w��o�׉�l�GKJ�K�!�����i��_�W-D�"� �M �;��WX"�2"�fY�=��j�K��J�˙=�þ֔6�%��@�%賣�am�b�w� r��Z?�G+��0�i�E��%8F�����<��S��m��I3B3�z�ۢ����5Hn�S Rq��W���Yt&;{Ŵ�=�Fߤ��9��M-���h����X�ɀSc5f�I��P*��O�d��rPh�݃�B�$E��>X��Ύ	M��n�{p	�!|�.�!$�"6k��VW��M2y=C����v�Y�w,�� ?}�s8��y������ګ��G�������o��`2R�@� 铟���%01 �a@���M2ɯ��[p## �:�}'�#	�D$��W$��%M+����k��|��?׷��Nx:���h4/J֔I'(��A��=�Xw0�'��P��&E���smN�Y���i2�Yh�d^���K���_!��4�#�p�܏:2�霋�����rRQ%0�kG��\�\>�v�mQ�v㿑�����N��gߺ���Yn�Y��x�ʮ��.N�� �C5��{e�	N�-���,.u�z�7���֤�=� ��H��ؑ��7�	�P�ZO��t%���Ea*�-h0򅑟�\��6j����[6�4��\M�Y���>5�{������2��Y���zլe�e���/.�<p��:�(��]ɉ:���<M|�qh9L%�9��ȵrDh�keT��_T8�a�A�������I2%1��T�h���/e�6���E�0��^Wd�fv>ͥ�.������{cDa�C[ŀɢt��a��A�P�H-.fi\����n�T���Dc( #6G(U3(�R+�M�tGi���KCe�����x�	u*'�N���j���_�~R�сTU�2L��o�ژ���eLƾx?��)�r[3�RL�z��V��Y w� s�IM�%3����'�fx:�w�~tF�ӫI���(�`o��U������ nmA������l�m�c���a��~��d@�\��q�6����B<� S��7qAN����P��Da�x+|���/��ip�E*OS�OPs�x��?��*�}�����f�U��iX�чRi���_6NӨ�ZZj��jS�h��/��gb1��J�j��o_��u`��72�>�'������ 7�m�<3%i���׬����Z��k0/5�^��A'"u\+ggo5��"FS�cdFpnڔ�=حp���W<i"h�->�@%����`�L�2(� u+�RĤZ��@��b�BM�,FZ��}�t��1&{=w�R�ϱ�KI)�A��� �:#���6J��OR�t n9��e�b1w��A5���O�a6Z���h���!%�D��$i-&��|{�>Zd�P_�+���=5ZQ\����O�2���d�$)¡R1�h�^"��4�_溚#g�f�R��D� ������:����1�`�	�~��Yx}�#�x2�.�s�����$�L�#|�Ă�ޜ����XMĳ?���AI�O�� ���_���@Jn��RyM���%{�^�q���aEG7oN�;_�!�RP��c��-�I��Q �!��ˏ��Ӂ�Vh�w��@z���I����l*붴`nhk� �6���O��*)�nԇ׷c�ӆ�6'�DH�g��O_��fh��W0|J��^�t��G����w�N���NI��Rٗ����<��e�@� ��D�R����[_���DW�Ĩ�K_�<O�ܵ_6F�p��b�S���I ~Z��N������-���,�J1������Z�r���cSOc�R�׎,z�-eX��D�46�j_� E(0#f�=s��,��d��D"a]�a���KkN�9��p9��j���
&�Es���M�G�InSM^�q0~�+U�$���6�j!��l*ң�U�[>��a��{<�z\�Q� �/�a�h�{��=2?�Fp���ĄVV�Nd�L
h)�yo����A}�,�F^��u9	�6�B5�4,_�B�6��;x$���
V3s�Ck��&)�u�$P������Z?��!G�[��O�li�p�\�<J^�#�<�x%N>	�." �7I#��sCK���^�9����2�6�t�0
�k8���i���~l�￾G���./�� ��.��xѲ �� 7���s�S��Y �*3a��Y����M}�=��f����N�w�n��a������D�ϯp����Y����u/(hK�Fs�M�1Qhg������P��\�yd��?���T�=�_������LI�c��"�W�|�WrnϢ�+�ﾮ� q�;G���_��(�Z�Zu�M�J�ۀ=�J�/"jmI�I
���,�Aը���/Nw�u�/*�^2�ʋ���@t���S�㡆�ԥvx}��O�)���e;1��?؟��h��퀫nFxU���Jy�G@�)*��\1s�E.�ڛ�/��<&X�L�h��I|�jP�fz��i�u����=̏2A%�f�1�O���O#���{U� �����ق����)��,�
aI$����b�`���$q��������Y�`w4T�t��V�Aq� ���Xo;*�`�
ua�	�
8K�W��\��C��$9 `�V'8����K��|���ҍHo{V�mi=��H�
����J"Ϥ0v9]��ߊB	�}Y�w�õw�W��ј[IBS���G��B����yH#�p�6VuZ��LU�C���}/�J����
J ��lݐ�s��M�AB���f�RQ��}ϫ�Ϋ��!������ő~c��۽� �ul��v�	$������͟�(;����C���Tz�'_����o��!?��	A�w9��X�'�KIȃ�[!z ������[(-��b���#P��E3e'=A��j���Ҕ�0T����& �3H R���|����5}D.\M|�x���<x$��538��3�/������1�zO��/�\("�7h�x�x����cP8��8{4xd�?� �ЀYS�2��qɽo �������N�bϴ2�v+�zf��߽�-�?�CO��2/4��&c���YK�o���
8�����Or��G3I�A�oD�D��zV�Tłb��b\{P����sN���yhd4_A�l��e��}R_�	�P��H�"���le�%&�=QG;�H5y�/j�NJ�{��D肘������(bA�@ ����$��\��'W�ST�����EG)��UB���y�^){T�O+�b�E,=��=s)[SX]K��Kl�{ ��g4C���$u�s�������`������p�$#n���x7R��d��?Gg�²�Vx�%��E��}O.pT�����L��.N�4l8����YTK�����#�蟲<�H�L�,'�PW\^����*w0cb֟�����]� �@�T tx�Դ�Z�I��|�E���g�!���U e%�<���"E�����[/�)�����צÄ�f���m?o�c�ٕ8E�(�V���R��ir���E5D'�	줋Aщ�ɲّ���'��Fvb�Z�a�r���4DżFI�7x-�"����b�9�"��	�l����&���9
�w���f,�V!�=�0HKV�6yy���=��]}�фa���v��m�o���۹�
�Y@��Ԇ��@LW�J�?lE6)��%1��V��;�P
����z�V$:��<����#�﯈<2<����6z�a�@�L񕼉gl�2Y_�: ��ܺF	c�P����f��+BU�Mj�T@����ݘ�/m�O5S$��n!��~7�Z��д$u����
�i�i�L����/��
�pgχ��圈`{):n�ɔ�hӎ��l����PUk,,'�}��NG�v
q���k�zgO���[�C���%�;���͖j���\UX����0�E����[*�p�'3;�Q�=X�����0���H0�E�bb���4��u�jWx���°!|[��`�%�43��Y����/��iN�����(�1�](b�K�,�s�8�	��n��q��E�;f55]���|h��-�:���.X��J�0yuf���w�Y0��ߠ��~0����l:��2a�|�<����T �5���X���;�"@˳)�ݵ���#a�&R^\�j���;��:L�T�Q�,ʱ��
;�pɸ{�j5bZ{r�M2�h8S���d��R�9<CV+��X���=���V+9��u&�t[����1��h_�1�b��ǰf�v���.�j��w2��уT���O�d�Є�GV=l��+���˓��*�ӈ�jbB�T���SW��I�&�&�K��a�kAlѪfr.���'��f�ܠ�r(��<��GP.�B��ֲ��I�ޫ�:�:6��S���B��X�g��li6������v�j-SS�JK�"�,�?�1��7�ȷӬڷ�rF1gI	���C�),i��*rT&ޘ�9�۠`�#}��-"��҂��Ԙ�^=��Ծ�ܞ����_|��JZ։ς�'���]T�����3�@�"Au�>��w^����N����F��l���c�1�b�\��m�c��q��˧#�P	�"��`���i�����6g��g԰^�������̦Uo�J��sRq:Aeٰ'�k�7�W��J�O�W�B&~�ё��/W�dO`�ұ{���R[���{Z��q���!R��"$)}Y2�-��z� ��h�!�f	���
=�+	�b�Α�ǸL�e EP�tm���U$~����|Wx�(����G,N����W�Œ:F���05�)֌��>�( �t��N�ʅU~R��Ml��25*ͥ�cMH:L׊�c�E��f��Ug����=L$A�����L������nձ�`�2���;wÅcN��-���X��"�ga�z)������<�[�;Xh��fP7r��!
�����9�Z|��/`�5x��?ڲ��$���#����Ѷŉ�;�O��h�9០���:�1��ॳ�[H	7�V0rc~��T&�x�J�����*���r�����-����d�� n��J�|g���q�%�=�p9��l���a#vV\ �[C���1�օ~q�4��u�{\���NR>jй�"�W2e�Z�$/�:���DA�/ylR��,��/��-�yv_!]�y�}������9E�6��k���R�:�����qaJ�斶��D0ֆ/e���I�2Npi0 GJ�7�����ɥ�r���X7�c��0��k�
}k�C���R�:9AC��dbzTfZ�S����y����0���U~;ï�a����h�ᦍ?�d�,�7�.�ۥ_��E�K�9iɝ�)�:�(�*���@��}���ɤ�V��R�1��R� :_���`8�:6*AX4���y�U��,ޔR�)�	��]`ẇdħ��	���tP���STǇ���!��'u�&Bw��83fenN�[�mM���D�ӟ�HN����&��M�b�&ݗ-��|o,�fH&����������k:�p��T�mmiُ=��	�~)z�xqWI���D���b���Tl*E�{�F�K�>��ȁ�kc�HY��#���`��7�hR�Ѯ"�������N�N�u�ӯPl�7Zn�8o|�6�H�R"|�HC��l�!�׷XmL[�a�b�����>�_?V`,�~po
�O�t%��#I�T,A�[0��q��u�,0n4 n	C�^<�2W��@飴F�k�(
��v�V��K�H8�� k
�T�*5��5 h�'_�sڪ���^TB��MH�bo���o8Nrh��73�|Xs檯�X����8?���N M	��2ۭ�����y�c�J���-~�T�h�F�yG�h%�zl�o��GI���^�6�^p_���(�;R�t���������4RF�����y-m���r��J��f��:�����D-[4o_�zL��!}�N�n�T�R'�\J�(�`�Մ@�&o�9�G�0zTŒ�-dK�X��{��P_#E-�gV��Ґ��.�u�"������j����b֪e@x� ���������U6�G���P��Y�軱x6�a(�^|�9I�(�ؓM�M+��
%��ZY�]jD��u^&1�<�/�����s@f�&�USWvS�S��G�[٤�'���1� _,|�8���ذ]�H��R�-��2Z��J��M��r-[d����7qC�^�l�5��͎m{Լ��W�7�V�Yǻ�j��O^U���w�i���2%yƸzP�E6x#��Ҥ����l]�
�>���ޛ����v��g�^��h���}p��%�r.��4Āt�n���*E��6w�+�:��Nu@�	?%	��N�՗�^LNU~�2P�$z�o� Vc�6�Nr�B-�_�ehN}�=�6f`TX����j��ާ�ߛ�f��`wU9���� �����7�9-�詬!p�P�&��÷�9Nk����ɷu�AQ�O�^qMM�f��\�y ��P��K�4�S:�X��k�e�x{.-�5~�7�{9Q��y+LO�-l6S���K�h�iV�v���S�$�s|�������Q�կZ����jf��~�廂6gD��G_
[��i���PNA�oa�AXjB��� 
U�6��Z��6��v�wm�ƾ1,�]~	�<���*�f���T��,}�T������ ���i�␹���ƾ�Z0*"����qd<���$����w����*b:Q���]��:�q���6.�;iIH�X�pw$fF����lZ8�eOE\���/ge��
��W������T�����%�0i�M�Y�����m���Q���?�W����*d�h�7�eIN�&))�Q��~���W'5A�7�y}��Z����t�a0�X{kg#c�7��A��n�i2�~�E�g�W<��P�[�Ől��� ����x�/����jYH�����U$����Dj�^Ѩ����Iz������9� F��^�b#)4��a�� �+����ٽ�7����W]Ě��2��}͌<�>��w�ͯ��yHE�e\ �Uh�? H�P�jş��NRO�ӟw�v�\��~�6ơ��*	��S����;@,Ŝ��,N�r+�\��H��Z�6Df1�3��L����
�|�c2�m�������X|m�(2��2���k�({�l��ֺo�U=G�}Ø)6�oܭ�w���H�8�5�>x/O�������zj�f�� �'����ߘ�ATx�Ykl���d�W`�H-Q�ND���uG��{��%��E���5�K��]s�0����GW�?Uцr鼾V��ZBM���5@y�yIe�x�B���$�`�$�԰4�}�Dc�� �}D�P]/G^8��M�F.X��Թ���g~�!V�s}��}�mm���7�+
;/�E;!y/��L<�i���B$Y�kT���)�c��`�^$���t�/=��fx-�2��W���BE �Z�G�}^ԡ��Ni|
�l��S"c����.?�(J�s�8�Nz�(xk �r��w�K�
"�,��(׌�O�"��. �C��C$##�_N`��0&"���3C����#�r�e�jbg�[C�$C�:�b�C~˹d�FAmkmc;Y��H{���oQ��J��#RZ�G�p���w��O2N��ZZ7�b@�a��mw	+�䍖͌t5��`�+��7���ԏ��0�w�=5}����:0���lR�i�Y���NnY[[��]�vwh�=�s`h �n`����'!y4&��P�M��1�WX�۲��wr�{�t�br׎cq��+컴�N���j@܈�����O�a��&�GJ�����3�IK7vr� �&&�-�*���<{��z���o��3��M=g�Gv�zm_�W.���[�wߛ���Mw����1[��L�fx�}ta\��E��t�� .�۹�/�M� Q#�9�s���c���F�%"i�K��Y���R&������&��ʊ���#nA�A0�*�Z����ӟ^J����̰ClX�l3�4�ڦ�����	��Y�C����sm����Cyɜ���`:�T4�9��avR*����!���j�Ƕ%��Z��=S�Jd/�����Z�cCɡ�����h�XE�y�J��e=]�r�`P�R+�o�gt�hKwp%&�3�͔i���� ��({=aliX	���e�OR�s0"z�Qz� �dE�����7n=������d8��/)g���NJ ��We�߻v�(U���L?���z�]��J_C(�q��\��B`����Fa���{+�����;�P�l��#K�F�noϯ�!�veYz�@5���ߥH�}�ɝ�X��D)����:��S�G��K��_�aֺ��?�k���UˢAAb� 2��%�8�	$"�k���1�sqƑ@d=���䰳�ģ���_�C��JN12��~��y�~]&&��)���AM�9���h)�E�-��󽁻�r�ӷ�,RO�cP��D�[�Ѥ�F�58��$����JRzt��d�ՉY����ׇ�ȉ�/A��kh�p�l�(��J��-�3����DϾ�r�D&�BaP��μ����i�E1�@�}p���8_p;�`��]�g�`�i�<����a�9�ںh�b��u�kӁ��:�2mh�:�J.=Jt:��}c�{�yw��*lO��!�].� 3I��!�u��G*%�h��l�R�@�J������O@5�hUh=E2tA0A�s��W�aS�ܛ1,�J��\����J�(�E=��h�V!s�Ҳk-l6��^X�F�d'�ٔ>�@���(�J��,_� Ւ���^�Ե	a��k�(�^'��Z%�z��/�r���x~�����֮;�ۤ��;�s����R���99K�K}�����ɍ��d*��c,���Y���PH�����,�^�إk$)jy?Fo;Y�u���A��xEh�]�D02U ��]U�BL��[��\�B�]$?޳�r)bi+�7�NÜ�������w�"�b���
�pc�nW�����7�.�5���c)�L)|�G`������n�L0��(�
ד���s"�U$Yi��srn�9DqM��o7��e��5b���wW�Fr0G `��ۇ>I�y��[���3N��w��W*i���@��?�Z��I��>�}�)K_k�9��c�"��G�ҹ3[i y��\)5�m��#<l��H�������so)8>�Lʈ��՞�h�*��Ԃ�)����
N�b>��� �d����Uk��i�S���F��	������q�$XĂ��(���{#�����3!d/�ITs��q�t����a*�K}�;��Ƌq�!�#>nCݬ��+w|7�}�0.��%�6��I)ݬW�Z��+k��$�}Op�-��e�3�p��bΛ!�G����m���06�op��)%�������Vi���8�yMh�IGO�S*���"r��{f���_"�{۲��SZ�4a���L��f���	������12T ؎P�:G�G��q�"�sQ^�D(�0jdК2�*��>Hh�Ll��CC'2�Q����h)g3Im�2��j/Jpb� �ܩ�6�/ޫ<]�%�jo3��{��O��s�c��^�>�cJ/9%з��+�I���x���g����ɝ�����^�2қt6�f5"�qiTKh��������)ҫ�el����Sw��ȸ�Ν�0�4ǃr���B�S��x���E˽�߭�����>;�ZX��������~�N��TێQ.2b�R���Wª�"5���S����.�0B��\�EZi~0:��s���Y�˲�(l4����+h0�CM�K��E��Vƙ�E�-n���J��݆	��٬ԯ�5�`����\	H�\��5<�V�p��w3��I;9���޸ Em>�~�?/c�ppmq�;Х���h�H����'@=�8�S����N�	9].�5��` �۴R3�z�Ϳ`��P�8g]��j��"u��E��h=�6���� O/�*zƂ*���,��Š��(Y��`eM6en3>I2z��W\����Z���+��e�g��+@W��EZ�����S������_-U��N�f��JJN�2��Rm���wT�����le-r��e��Fa�煪�:���ewj�r۔�>ʲZ���Կ$Ȓ�P���W�}���
�ؗJ���e-�R`^qʵ~`��[�b$,���=�G���+Ne�5�t�7`aiW�[�.^3�+������s���<��e�a��L�a��v6��{���G;��.倵��kr��Y0sGy��"��9D
��]��!�U�4�@p88�r*���:�h��ė���?S�ƕ�$�'�-M���������i���l0�t�"y2aE����N���Pپ����_L� s���t��E���l��],�������D��vzK�=-��������c�s~�� �,D���v����.�X��J�C:�w`���ⱐ��;Yꃗ�xQ}l�h ����mY���ٗ�c��=g����C��A��z�A��S���2΁��C0qB�UrmI�'ѭ՘6�s���v>��ȇ8a�Y��)���Eڼ_b���a�;���&r����D�_+������1Aۄg.�f4��nBsyM :�1�%v\'bx��>�_,�W���>Vf�Eӿ�P�E���yX5\���x#14�>O�l����Ęa�r%3n�<�+2��.*��f ս���%!�k�T{[,�ʂ�$�Gj#��K�.p8��G{�3�ǯ�7��/n�ӕ-��g	�!<$���IU;����/�ߝ�{�К�,�J�'z�(i$A:p��U�-7��h�t>޸<�1�AwG���rU�16��s"�cha�rܪ�@d����i�D��}�JTP4�?eu�RI��X�R�y[��ޮ=V �XG���I��=vK-�U��$l�NI��"��٪����a����T��ʁ7��3z{�O��x*�����e���hȾ".��T0Ċ�U_v�h��9&�c�ό��|�#%�;�j�osz:��9J	fo>�T���;H�8�:�T	�S�m�r��M����Q�S*�Fߔ�  qŹ�%��F����aKL�nټj���[' ��6���^$��uk��[�[��r��3R�d�����d�xF~K�76V�l�����6��������g�fD�,���ޟA��q���<�PCr����Jg�?g5{ރ%�v�LP������
�ˌ��#�#��qD�3B�L�����f�4�+�F��[��� )�h�GP`�6��z�7'>M	ۙ���W-�%4�/��%F�t�J�.ԾUc2��6�8���Z���q�Y���]��">E 4�X�hL�\Q(я8>.<=j�"���k��Mt��ܽ�A��K�9i�Y�U{%�ə��ǆ���ת2?�&�:(���H�;��4�2]y��&b �Ɓ�� .� |���\0�m-L�G~�_����\qT��/�"r	��l"c����ivy(�s�DV��x�P�i3���۰w�.�
g�+�bl�}�G�N�y@ʛWV�hN�0�u�F)��n�}�\��xlg,r;��LHw�lG���A!��0���.Գ�)�xmO��E�4��H^�/GtA�7�rxF$�0Sޙ]`���-��_� p"^�����2�^
��'��͠XmE���v�UK�u�����A��F#�ҩ�:vw��p�*JB�{�����]�oG �!c�ԁ��ڰ���G2K��v+R�g�^)�L�RU�mO��	�}� |d�QՌn������߁s��y� ����M�s��8��s�Q����R��porЈ���J �ܿ��w�{r~X؞�z�Ĥt��i���Z��j�T��I���զ�*�6&��NHMM��s%��Z��{ 0�Ų����E�Q>�&��&'\��7��YSB�X1yS)�� �2�6@x�'�{c�f�$�$D
e"i��e���OcU.co�"�Ire]�Nh�S1���!�L�ז=��2�=�;]�sV�U�X�&A��uK��}�}��	��6\�n9����\��=��{����Ҝ�?ҹ��"_.���B�����wȴ���g&��\���/p<_�� ,6�<8|���V(��:;�#r��|B���0��]8-��|�T��y�;�v�����&Mb��ӡh6Hܗߢ	Bs��%|J��ƹ3�����C�e�����T�IQ�9r�v�B9�+�.e+��U	�hn[63A�Q����Gp��R����;���i}ǹ�X��By��������n�k�͸Z���ܿ��C��w}n���Mc���Ͱe�|$T	�]|m
�k;������W�]Fd�8��B�]o�Jv��V���q������נ�{�T�rc���(�ܝ3Bq��m2�ߊ1�?3��#LvX����'�Y�~N�[�hi����$	?��(���$�L���^y5��A�$��+���s��lQ]�_���.jE(z�c�ب�CV��Kw��! �����4G�����u�4]�P8" ��\��0i���x����<��;\�J���	6'����N��+)n�6FO��׉�@V�q֘��PXo>�p��Q�����:�=rޓ��Z1V�cŒ0�򜽢h�</���d�Q�)�J�S\H#�g�\\�����J��$��p�|��?�}m�789��5�@��`���j��J|6���ެ�@ta�?�m&-��|��7Vr�������%��8�7o%C:�����0�Uw4�lQi�K��O�P��z��P˘�xg�p��!{���Ύ�c�s����b���{ bPkS?��	jn[c-˄�Ȭ�6����>��ci
�,!-賐���-�,�{�/(�� .+B�� �\u7�o4C`�"P���yPm�y4���{�X1���N���/��l�d�,&�ıH�|��~ʗ�6��|�n�T����e:`Q�mp�֑c%�#�-G��}�Ś��Q� *�fہa%��`Qŗq� GW��{l����Pۺ�t�� ��jM�%�4{Y:�p���r�9��]v���i���*�|U���h;�����m�����F���d���`n0�#�#]%NYj��F��0���:��ޚ;+w�9~�.�i|��C5�=���r&z��,mv�cu@���
ϼ�6�b��9��\	w>Pnx�W�r8!-H�98ZD��2���aUE�FOb^#@�tpN����vOF���@I��ã�S����|l��#���@4���9q){����nFT�4D�%�����������MF�#c�eF���Pm�$K�P�*~���dM�k8&:�
�D��.���u��M'!Ќ�&=��֊ca0�|Q)�6��?�إZ���_!u����]���il�	���88:�r��x�����z�	gr��q�Mzvu;n9*�כx(R��C����G�nJ�L�)����'<}y�If>���_�����>U2^Dud#�k�Yl�:��������B���7[@t��W�3y��%l��S4Vm/l�9��Тb�S��Wm܃;M���;�*3 ����s����m5�50 B��ÊJ��H'?��Sq�Utjn�nۥ�18���=���Ӧ���م0�;�̵�^�r�X#�C��)i\j�ֵR:���7��pFu�I��pY%�2ib�Xה&C�
<�vQ�I�d����.sz�Z�J�t-悈M�1!���°�i�=i<+�i�yl#�U��w3Սk5s1���U�(Dk6�޳�r���?��������a�H3M�d7'���w�����Պ�-x��qɇ]��j包)�h�p�}T��E,�3\��q�d���:���}�r�BJ�)T�=�k����> �uD }��q;�:�u���]@&�8�w���"d�4�/�����j1�p�T�:����2S�qo�����������}�����~Cs^�X�5�x܀1�+�X���@Pa���
�OT�!�{�^ӿea����^�����4�+o�~3V�����NC� �=�Լ��t{��X���(��7��Y��wf��m:km���i�m�&-������D�J�?��'��D$+[�*�����&��I?��o�">pI�.�=���1�]���~���K/�e��{��j�!"����f71��:i|u�.��&z�M<�����#��{̠�y,T�E��\8^K�.��a}��1��aH���I�Z�E�T���'[}�(@��GXm!���[@�Ô�=����IWG|��Թtn.au���J���&�"~&�py��B:�[���ʌ��$���+�
:}2�_��4��G�H����x|V�8����IB(z!B|�FAv!�THE��r{��|�rJ������qtE�$��*r	�M��vBfԂ�a߬�4^��t�y;{�P$ƃ��>���
�T�{��gh�x�;&vb�B����듵W�K��|
��%hS�!���fllM�p���m�\�(;L��so��g#�i�r�H���}���5�z'�}9=q.�`��P�M��Zᇧ�Hh�`��Y��@�T2��pP���s̢5%=�ب���4:��&�����Hn�w�&��^��&�o@p�=���Y��b��OjP���k������dY���U��6C�pk��{}����_��Pӂ��MpUw}Sz��R���ZO�l�?�X�⍪:�Y)X��YL`�z!=ߘ0� �n��"9�n�we5Ίz��m�r��Bԩ��7g��-��a�[������7��`�;}�_4���-�8�RN��gg��k$ �u.�j�4x�W���qٔB��{ 'Al���[��94Df.ֲ=C�NӜŪ��gp�;���	�A9�b���`��Gܷ�g��O�a�P�1�M�{�;jm�����T�����H/�bE�/,;(����õ}e�w�kQ9TQ7�2���r�i�va��.�+��/��eb�$Ys��$2F�����$�W'�'��L�� �|�H06Ѹ���1Ԭ/�B�nA���+�O`�,迕	�	T~/�lO�.�-(�}�ly�۸G=�8z�4ϊX�9�n��}��HA��u�O9�r�K���E�/H��t�`��,�7�$��۰��h��G��D��<�A�C���������l�(nV�#�Y�0�%;<�=���w��Na�'9?�*�
�՞�H��.�����3��	ї7u���� C����A:��F�n�<��N�������4��C�+$����?���j�<�q�PL�[ĂUM�)�jĄh��2	��&7�����:xX]nx��J�M�s���(�AH ������+�Q�gi��f��ET8�L�2�9�o+8���j��W�&ˎHlն��7Si�G�׋3�h�:�o^�.�� x�����S�mP��
��d?8�V$0�A#�n���)�Գwv��а!���E��^W�\�Z�Jvɧ�7������0��u�6_ڶE����5Q��a53�$�J���2D#|nFuC�0L&�Ղ��M5��^�m�s��y�Iޕ����ˀ�e$�IZ�?�n�j�f=�V��n�aĭ���Q�"�v� 1in�6^�GhPJ���[����~U�w�j��ȃ���5�GZ'	�2�a��9�ޒ�Ϯ��/�d�7�#�^ǻ7�ޟJ΋i��$|�Q��
v��x��-o�ot=��6X FX斟ؗArH�l8`)j��k`6����`Ra�\gƏ�t�$��e�d��l�P�do(��A$�'0���80�|������Dh0��#'q�:�7��"�������S�h�>*��=�.�y�`�"P���-�����ݛG��*z���}�\E��wp���D���DLE�5�����V {p�����r�/���<HG�a��~�(�<8�c�'��|,я=�n��!�=�{�$MU%G�8r�����OtI�Ķ��הM_�z���qn"��2�I���a�	�"��� 8�	|���˼P��w[����f�.+��	�?��1��������%���}�H�L_酓D_��r�r��ф,�5oi�+�R�8�+&���abAA����h�<z3MJ��o8��W�%o[n�R�brbŽ\q��ѵ�g�YT�^؝��hū��¢��D�&�R:mM�z�_'Q�~�r�g��듘��qF+��}��x%�z�͵�mƳ�-Y���w�y/��L�݄0�%/�H�to|���m	P�ͮ\9���\�j�������du��8�>@��H�!�
}YM�
����z���z��3`�'�K��hKܹ���+e,�}��
��@�i}�'��C��TЂ����9���ꍥ��l�9����e�su��z�s�"����s�;gm�N7c8f�M�bp={a<�[�!1C8�gg�-m>`�_;CK�`dqر.z?�88�*��[T�g6��t<�bb!���чF��M�ʅ�4aA�E��� �K��V��n��4��I�<]٘�O�'I^3�g�W"��|w߰PD<R�eI�L�Ο�h�.�f,*F��WڝSs7;ygt��q�f���q�"qUP�i�P��^\���֢Py�7vt�r���I�W��]�Mf$B�ڢ�2:%|��5E1j$-�CV4F�y �b���g�6po,;F)i�%��ڳj�l��"�{��
$~`(Rdn�C�������˯wa�ӏwZ��_�+\
�V9�SU�j���Tk
��A��F
mr|�Uo�P��:�Y9q��eW�뉝��_���|�|����c�jK'z����Oа���IA�(�{�c�(W/�c�%�&�E��B4Z�]��Lnv�>Kï�����U�S�$���%�Ԓ0����S`�$�w�d���-��󠄨�����4�n��;��g�9{N��Gd'�poF_XＧ�ɥM� �MIꞙ�,B�9�A|��`���{O���S������KZ��h��v{c?�/k�	��X��_6�so'���H�*"��U#�v��d}Ҳw� _�ngu��wz,��8k$rUv�Z�F��)e+W�i*	u�ؼ��<��$����2]R��g
�H��F�V|f�u؋.(Y��v���������m���G�i�j}��p��G�:Q��޳O3��R��'���,��5�N4��o�3tw�瀄�və6�I>�����._x���=��+����!��ܮTOj��/
(U�մ����s圛��ۙ���*�+��%\�	�i�V�֯T�����-��e���.�x�b�嗁�>�I��f���e*�@�����\�wڂ�.�K�Q��<�D�h�J�s�/Ȃ�18�
@%�C�X��(��.�@wr���+iT6��)"^�x�.8�	��>vc�z������.��-OݧHaO���|��
���eX��#8�j��JΫ�Ӎ�z�E�u.l�+��D��u;H�KJ�8pc$T $�FΒ��Nu�Wh��o��^P����Lޫ�eL��9���u�'����IJ���K�q|K�YB���h"��r8���(�E��~Y^����9< �Ӑ0I��)��+�0C�\�a� E�%/�I�O�9Gc�1���7�:�3��=�$_Պ�Q�L~�����Q[O][��3��&g�ߤA؝Yf��U�_���>k-�����|�N�6%��7_@�t���h|.�x���[��s�H��F��依����=o�h�C%õ�yE�$��W�i�z�'�SS����"��Bt�&k����G��#���GO �*�X�&���r��޵q��-6�o};�M��o�;n[Ճ㽦�k�T�ze���Cf熼�ڎ�
��L�'	�j�맬���˥}���)��4�r*l���uz~��}�6pw\Mxω+N������J>�fo�U�qA��L���j��+�c*b���M��"�W���+��;�8�s&��_�f5�=�,מ ����Fh�S?�5FAK����hřQ��67�+�?d��e��z�]�^�0E|]8� ;6���K/�^�b�0+��9�rH�m"o�Ŧ�!ņ������{��yp�&.���>,����yH s�"T�����̔9�^xЭZt�K�jH���g�Ӭ�2�Jk�A�:�W��CWB�[�`���W��ￂl���-�rFY��L�b<��.2��𡺴0	�i���O�s=9^�$=k�ķ�2������������#W�̕ �L�����}0�e��ؙ��V0-4���KN���Ÿ���)�#R�M?�Hh�z��� +��j�-�$���1�W��qʞ���1槤Χ\>��Lh�kh��
���~�*�1�8=��HwI�:�t��<��Zr<B�h�z��������y��y�Bꖇh�(Y4���5��?\2���ʱR��W,����G>\hp������ЁY�T���׭���$迮_g�uq��}�쒀�
����v��?�>ŉ=f�}��o��u�� O�M�Ab��L���3CBb�;� ������u�y�uy~'K]��lj2�&\B��ip|�U�o�R�Cph�;o�"E��S	C,뉗����!LM�v`�00 :?ֿ| >?��p蓍xE�-��K�y�@��#�Ǜ�N ���m�|<�/*V���*�ʋ��~����P��r���@�E�#d'�?Yڼ�}������,�2{��ny�&��MFbm����&��I�BjM����Ev���HH�i�j��7&���*d��~����XV?d�N����Z����z�L',����e��ۘ�ܫ��q���ή�ICh�J�F�@��/��>�O��&�2�X;]�����0�3Q�"�������`ǬIϕ���I;v"�G�����7`|R�����1�|/�*i4�qq�@��{��y��U������B�W�?ѿI�^�	�xwu�X�y�ja�) �~��̆ ��:9��3�{2^u�@u���i�o�}�N�FST:V?�\�J�i�o%0��yW�a?���!]�ᖼ��~9�����)�3\sH�nB������2��搎�u�*���l4W��<�+oq\GL�M��[����!�(��P<�v����
�y,��.�>��x7����P��K���S�mf@��zH���=�-/sL��|�� x=��exR@�^���8Юǩ8 �9��*�Ŝ<�tU1��lt���T�F*۞�ܕ�\�O�q�2�c��ڡG/1����jB}����d/>:�\b�ƈ}�ɹd�9��6��9"�oT"i��X�F)J�J�*˦�^3�z�?IN�3ښȸ��
��jLrF7�mB$�z�ev?0%q����-��1F�`ʩ9��ؿ��A�DjމЭgaKk�{�/+�h��k7k�ǵ�]f|�6�����	9��7�٘׵�V�?'��z��;��S`V��,�����y���j9��!'��F�|���Qy��B�d��Myew�JC���p�MZ������� O�1��T���:P'�)��&�����3�;��k���<�XR�� �(����o��h7l�;��xm�~��2;'c�Q�T!kf�vT�9%j�9	��D=�b1ǌ���%|�#;���Q�O�P{��t��FYU~�2	]��B�;<���e�����z'W~�'ƧT���^S|3�2����}i�H&�0<�.�:�yd>Y� x��7n7���u�!"�Tu�,�!9-$������2��B��@:ʳQ�/�lB��e{1�z��$�]�܍�įY�Q���8�=^:����^�aN���35��1u�v9�w2��1ن�7�[���iq�Ke��ǡ�w�/W���3ў�ؒ������=��1�����_W�rgҦ�>uG��G���a�ȶ['��X"fPe߉ȡ�1*��t���jx�h���qz���o��ٶ���D
���������ة\�'=�.���-���
��T%�&��~���s�K�U�u��O��^�(x�� znȚ"	blR`�T��2~p{����H���p!��!�8/!�t��up�*Z5��dSc�:���+�pN:D����ȶ����$C�̠|�2F|/EKϴ�	.Mt�����^ZuZ�3�����ĈcҥD���������YBR@>:��@fr��bޟpt��'�ec�@=�Х�vҧ���w4�AG��Y�X=B����@��eV�:|9����bga�G�vU��� b	�Ϥ�态�m�;B��gE�i�e�s2�F�d��o^4�sVQ�q}�i������	��*C6�uɫ���M��-�|/�v�<$�����5���A��)�C\mU��PW�L�|��|Mօ�Q��&ڕ��F���*�?"�a���}$eG~_\�^���ǡ���L�A��J��k�$Z�L]�G���[����fKJ����;�N�À�����%��S�.������9�6�u�l��C\�:��:%(jS�"�^�ׂ�j;�8�狳3f�&m7�l�ևV"j}m�{q�"/7 1{���Q�еp�����%��Tb7�ch��
uL`���iH�
'��@qPљOQg�G����RT�2](�����a�h!�ەԼt���Oʞ[;�O@�&��d���~J%_������2�QI�n
�E$�j��� �`]���|U��j��o��2~��L�
X�7ش�M�M �WvV���2���8Q8U'�&�z�z:xV�����?��qO�<|$��8/��Ƿ��VP8�j����x�z�{y��Yl�^an����������t��1C���4�����^F�N�TV4��i0-�V�����ﲀ�#�����R�iFd���T⩚U�r6z��P�g�f¶O�rȧX��3�����P��ϖ�B�>��q��"Y�Nr�M���4\�{V��P�R�����j�;���5���?'�6��M��I�H�
Ep�nC<r�y�[�y�VP�:1uݼ����=0=WZ@!ml�o
�J ��:����±t�c���\s6Ϟ����870� �F[Ga�:g�T�n7�R_��Qj�����kB^�͐�}�Q"���_JɘŻ�������Xy��3!���3�c�	�Qم7�@�9b�O�*���{q`%?� �j���$ϥ<\����s�*�5��g�\�ꛘ���|��E}.k"d�(�cG?����j�_��?�k�RU�����]�jb��Ђ�DòG�ӖؔieB�/�OU�ȯ�"�*y��q<C��Mh�M=�����*�"��p��r,*e��91��V\Nչ�~f��$:��	RT3
���+h!2�8lR��0�A�C���\e��yZ�%�?-�c� u�gI#�ƃ��}�N��gР	�C��:*� ���-��f�jT��Y��q5�d�G]On$�<B����2�h��2Hg�������r��&�Կ�|�؂w8-��A�0�FMg��M�������}��.�U-Y�}#����َ�s/jx�4����H�VM����ŵ؃���<ʓz§$+B%�wh��W���?ˎq�88�i �+U��|�!�z�u��}��v�``��R�v&@9	��ey�6��}z��1�?eJX�қndzc�j�P�7�u��W3Y�����0"o3uu�
����3
ҬԵ�O�
���fZ�y��%S��K�ȶ�xA�ͣ�����!?ڋ������X��'
N�s6�ȥ�7�L7�FP!��s�Q��wi�$풥��NY���7��g
%Sx @jk�NL��%��ݠO���.�EŤLEu:�|��]y����^�Ȏ��V��%��Re0� Z��+��j�o�}�����9k�s3n~h���%�adO;΁��;������p�Rܳ���ڜ����}����=+r�ǎ3��=Z�e�,d��A�3-�<�����>�VHxt���6��U�ݩH��ld���d4� �����-W-�8Gi
`S�:z�k�b�1㵒f�O�9��q�C��.��J�d�Z&Yh���즗|/����}-��2�q�}l���hh��Q����,�yU]Ǝ��Hjg��2���H�gǼ�(^�m�N���cC%���/5�~�6)��m_��L���8�n��"Un����-�t7�߀V>v?a�^k�N����{n��֔v-;��q����rn���g̙۩��]���i��~�_ȑJ{�.EO[|V�%���.�`�\�M>D��\�]�d�#G�-Wp�Y�{���\"�i��L�P�Z~x��h/�9�ɶ~�'�o[]��$�
�?�?N�>�����	sE��!��v�/������h�	�=�M�V��y�D�a�ϯ
0��t$}堿 j��$�r�ag�P-<�-�}��ުr��|S��d��cu[u!�1dtӬ��R��5s'�&��V䓝]���v蝌y�kưx"Je9�I ѯ q���9�ڌՀ�
�{t��]޿��%�����'�����}i|�!Jg�1ѫnm�;c���9�KJVq��fA^��C١5ڢ����E�'��"��e�{l�;���z�+��fg�9=�u�V��s�)'`(�o��Q��!�0˲[d꩚8<�U��Oс�d4W��p� Sun��J�*�l��Ei ��˙@Q?��:y_柃q��p���m��j����9/�N.�
O���Bi��MRY��B�cD.�q�)6���1�{�I��K���APl#�=�e���d!�Co)���V ���[�뙱��dS�4Ji��������\,���eX9vs/��i��؂�y4���ՙx����E�XaC��?�5����@a��i�L8�M$ߕ�F($��Կ=� y��HkLԋ�I�h�n���,�e\�.F�/HdȠo�v�Ey)�И��v47 ��Nٸ�`������M���iДj���^a2{[�S�#���Y:����?����G�T�:��X�����Vׇk�y�;�7PU2�AzӠ;�����61��ɒ�_�ohA�e���P�T�X�z��f+ZA�p�֤U �
���V�R�+�$+�:��Ly>�z�mSUd���ݨ�r��o� M7\J�͢'��៏ֽG�F@4��j�֥�B-�L8��<J>�N1Y���:r!�xu`q'�~p�b`{/��Ɉd��%��~0�V�h�['��2yЀ��6���H�7��7 �'�c%)�Q j-�g���5�D 9J��E�KAMDb�ZJ�S��	�A*$�I���p&y�A�K�HbH��C�6 b�p�Jt�>FUٯBc(v���n�N�-Wpg��p�G2f-��g����D�S��"�YT~F����K/��8��
PQD��M�ac�� b��Y���&z��p�K����>b�o9��(����+�P$ȣ�gL��E�lzg=icd�(A�o��D��������2�����AX��acp�='lOS����*N�+%X�0����Ab�i}�ʄ�%:e_�]P_l:�XsKS}5��_`�.����N []�#��A�;�Aw����,����#���̲�C�BG��%y;	��Q����v�a�������5 ����G�&��h��GZ��R���v�� ��҈9a3��%x��3<[��!TIK���N��k��-����^��D?��`ҽ$�;���𻙥S��x��5�nQsD"SV}aCb9w���k�5��P_$1���gG�B n����g�p��38�����as�e�VW��rQ�\����G�i�+]~��n`|� _B3ﰹ��Vp5XL�TPG_v#�"�F�y.��7݊ԃ���2?�;������u�$���!���jf����k&h;`ٓ"<ʃ��mD������ ��&p��W�MA�/u��hq�l�qK����� f�@|k~5��'�L�4d�� �t��<�t?����)�(���:!eO����;:L
���M�����D�!Ӑ�b�Il����x��y�m|��ɭ��):����̞C*] �ٍjZ_��"��I�}��q0�3e�w?xYn�l��a��'ڛ����-+r����Y(a]y(�y�����ѧ�(�w�i������X>Aj�����9[3?w���f��H���|�}�S�āF�H��>�sf��Z���J_]�_����j��X���'�8��^.����!�>8W5D�A�Zܶ܃��<�"�W�+b6*P�S���˕\�l@�����
y�닕���?��Y�!�y���'��$�X0qB�\�,Q��߉�(�,1v48��v��9�f
ݼ?@�mn���䠄��wl����X���b��_�D�)L���婚�<J����-�Vq�9��)�g6�W������{�cw����iXθ/⺳��[�MAXy8�0wP��Y���鯟A���l��z��b3�Z����R/G��QC�$`�v�\��F_ۺ��@_�XT�`��.(\)/|&^"U�P�3Ʒdy����Θ�Tn�Su�4����/�@��C�/����\��8�8>��p0��O����a�=�NC�]��y�#�Z0��2��@�mI��*���JZ���5�ʪ;��{�f��E`��uؾRrC���יo_�|��f���="��&�?4�lb��8X���&2PcG��~P��<�+��a��گ�5�NV�R�D vVM_�chi� ��}��T��(�Lc	�S,v��(����`p��jN�=��TU�qK>i����!���\�3c����C;46�D��$F+����O!~tY6���!�g�9B4�/6���:���u+r�W yrր�2��j�qA�j�ݽ2���������g�={Ԗ�AU1����-�$$�~�S��iJ��b���V�Y�;�]�tDG�QO�V������׆ul�D�X6iK��H�7\
q@���Q�~�h���	�2I�;��$&u~Q,��~!��Yo|�� ��0u�ί]k,�:�9s����@$�[ϴZ��$���ߟ��?���8e=�ŝ��O�'nn���N�Z�`��.��Pe�+�E��{�t�ݻ� 9���, i�&�8i��sǢ�8p�"���M?�fIR�w�0/ c�8���%�F���'��Q%��82<T�hy�)몯�ZJ�չ�mI|6�qm�'s�W.�u�=(ѵ����xD��m/��k7�?w�
��ٚ�mk�-	!�E��:���
>hR"�L�~�儲�S�r[���Ĭ�b�9���C�����H(g��{f6��,�j�c���Ȑe�%�� Ngp�"uDV�б�:LP�2�4*�<�_U�m��o}�!�3(4��{�K�Y,V�ۂ�kG����C��2��h�n�qm���Hb�M��=�V�e~轳'z+d|Ҝc��Es�ǆ'�wL�ݴ����/�6���t�*���v�����9D���p��(�t�f;~8��7� 1��c�R�O*4]ww���I��WB��� �*]T:�`pi��?惲�����R
���r#�kWM�6%���
|ep�L�3�Mq�\���G�
X���r�H�Z3� ���qPHV�dO���}�'$X�ٻ�DxH�s�A{��!���K��o�9f�
�v��NV�>��4�
{)Qɧ���V�3���׊6o!�\aS1*���}�_�C?��P�U
��]�	���;�'��M�^H�g6Que�u��B��`~��)I��F�6a����!�T�NB�I|4`D���GM�[��݈�9&�����_W�E@f^��E���ztJ��ߧ��+��po������+b�g3�jW���,7*�e��f�< b����#�
'��2�W�`�D����f��k2�9�j�
پJ���gG�Pm
��Xs��QXf~�=t/�9�ɻ1��?����"�%�o#��pJ7�0�(���RP2X�1�HC$Y�f�Gi�敯M���o*�,Zے�A��T�l�����S����񞠄�b��P#�Y��N:ہW�H���쯺�K�'�5\𭻴m��>��q� 3t�6�z�K��j���~����V|�NXܭ���$Ѧg��y�1� jeҸ��nW��!W,$�����l��4�g^��Ө���tB��(jz����D�lw�^7H� �tr�^\3?�c��e`�ĳ�=Z�)%��}� �[O��5cN_��T��)*%����y]G.��`>r&P�c�6*)
z�[��eԻv�9�7*�1��+���*�۸���@ՊbE���B=��܄bc�2|�!�����F{�>+ǇQ�0�W���Y�)��A*�̪�>���oJ`��W
2�P��P��W�d�<�wCv�_8"�.�h��LHI����2SĪ9�w ���C1���?yׇ��Oר�̹��`��ΐ�������S�vQ��v�.@���e� ����ImE��H�%O��N�l/{��$�>d*�a��x����ռ�w��痓���D����4fp���Ty����'�r �v���F��au�)o<�BJ�^����餒N���G�u��Z}��ľ��Ub�[��U���?.^>���'��4��6〈pW�t��Q�����OW� ��5�JEpPy����аt�L�QC;_w�����ʊ���p�/�7s��e��G�8j:����}������o�c���|	�m�C9���})�"&Jj��刣��e;���fIn��?��f;) S��q��*e|[�	��EC�*$�s|pf͚k3����ʬL�;M� 1{9<0�d������BV�O[�>u���E,V��:�i��G��w#`���*�bv��\F�N�Z�B��O25���3�&�f�Ҝ�i<��yBk�՞�u�!=��`�{yz�x��dI,�8~�q*&���#`o���]{Aڽ�	S�������UL�$���oRe��E�cș,J�+<�o3�o��l
�n���<�4K���#%-yU?��b�갰B�Q�<G����-P���v���o�@2 �+@W�9���<-�k^�n�����ݟ�lBhg�.�G;#~4�m�i|�����Ў�����s�}	��� �Dx����$���ty�m�Ȕ����;|G�/#i����k��Q
JAx��)+��E�;���&���|����n���t 9��p2�y����f��N�FnWI�n�w����;1D���:d�=��:O���<�Te�tbv�}����I�\QD�u��*��.�,��UJFȴM����w��0���<F,Z5��N�N��J*yV��sH��ʈ�rژ������Q�G� �B����
��(
����%}OH�k�&�0�'ͥi��e����/,H�����%A9��v�O)0r�yN�}���{1	�Nk�H^�$	'����6 �4g�_�Ͻ�^vɭF8RO�`���{������<�Я�p<O�S��)Np�ej'>*zy.t�W���l�WA�ک����R���Ζ{�\�6�{N[?=���)b���b4���Y7N��w�!a�@����.YNIg���{Ʊ��Ll��b�A1M��E�G������d�f��\c��ldKAf>v�4�[���>\z����_�*����GU�͜`d�����N�W�K�9[�I���sX��B���ؾ�8� ^�4.qZ��_�%,���dܱ�7ճ��W�a�<�	�u�2���y�B�������v�h,��mi =����S��0��6�<Tc�e���1&+#4%��&,6�Y��{��T��tA�W��"Vג���|w��?9�1��[v����WQ�n(��&r�3]|�a罿f��y��[�u3�� �՘*,�*�.�|Hs�����d�Պ�G�nM��.t�yˇ	�.؏��ʈ�#��g��T��kb�����1�C!I5s�N����M����_ڴ�s�nsfΫ� ����U s�ć�J��ytI��gr'Sm�u�JQA�V�������Z��wu�)���Z0�A.����/I���L�KSz���)�k�Y�8��b��~����R�)�]p�F)�'�Z������B��$����9�Q�*@dOX�ٺ1b[GI3�i,�=D�� S�����>�0*���\���#��� 6 ����ϩp��q	eiK5��Yg���Ka�+'.<��o�A.���Y���I�ٜ�\v��77*�wA�0�6̕�#����ѥ��1��٭i4� sT��qG\��#�s�'}���S\��R�fEI:kB���k��q�*���2 ��Q*��[*05� �N�'�l�f 	1���8���ZW�orlw�S��~��ߕ�xx���/Q��6'�/�T�ѕȝ�b�H"�0u�P���j�Y�D��	�џ�2dw�c:޸��_��Gu�dIz��m��0��~�/���)�=�P�Z��$�ю�Ba���6qLР�
	B��U+	��]����vr�����p�<���,�b���E�	ˇ���� {�+��}�T&D��GN�J��4��f��B"^��iED���$l�<I|O@�]a6�g��׵#�iݐ�v�QkX�-<��j �x{�%����S��~�Wi��A�ƪy���hw�(j�bir�6��,ӏr�oy��A3E)n%v��'��*���>�޺ �����&.rgߠ�Z�����\���:���/Ua�7syAUDt��''z�XFGq�M%��Ga�C�GA3�_�Cvݽs��J�^Q"x5/��j�F��;�-�2��i�Z��.��h�A���+<3"���2	���{v\����+�E�T��1���j�B>��K;6|.����6t�H���q�`�YTR9�)�n�X뉭��=�y�_X�8���뙰�m���l�Q���Jl���A
�%Qw;�kI�1tK�*�y 'c�&��_F?��iώɪ�)C??n�ٴ��5־�"?OY�`���O�7��1�-�3W@�X���{!H��ۻT�t4���Ԃ���#1��������5:��p��4!G�m�:�E���b�{z��<8Qaf�P��s���Ol�&�ħ�'4[o�Gf�����>2�������KU7����Q%��r�&�a���gT�R1���0�M6]n_+��#A���j�-�j]�2� ��'{�Cu���@lz��o��"�|I��P�}t�Bix��e˳PrM�)а��N�.���j���]���
F�w�&qau�h�_� �6����\���J�B����N�N�Ld�3B���qN-��2U�%%�!��V0$�?�[�fM�ߘ��yp9m\�/zyy�ZTˆ�'F�c�w�'d��.���x"'�o1~Ơt"����N)�6!��N�!!:������GJ�o%x�ЗU}#�6ʰ�S#d�����wו����ҵ��V��2��>+D�s�^g�-� 8�az]Pnl�O@Y����p!Z8,�^0c�I{���N�sO�a�S�\�����n�Vr�C,w����%�N�B�0��ތKH���l<�ٍ�'C��fH{T��a=+GK�5�OB���A�_�Q
� c4�%f�@�	����G�7�F���Z�����Eՙ�R��b�iM�Dm����5���'Suºt٣Q�"�,�:11���ǍXl�[~Д�Y,�!ʸ��FoR��FI��t�r1�K����&U�[H��~7amω?�r�'(�$�����,2 �-A�s3X�@1��F4C�����T��XD5�+�I�Z��Ifq�"�
`'��u�+cd�	��<��զ�J�����@�>U,�0�᤻��@�vO�{g\����9
HǍ�YC��1�-�yzSw`�^kE>�8	�9jח&���c��V���^����9�~���i����{���<���(����^��w���	t���@���S,�PfU&�jp8]T�Aۇ�o�f!�w�r�ϳ��}x�L�?�4�@�NxP&-k�;]^�,�V�r�4���N�}!��;n�p�!~�<��C�+Q��)�TX� ��1j'�%vM4�ѥ�	L�"��$/h-��zO�	w��6��|�8"���4v�sw+�ރd�N�D������uӨn�!Xn(��#վ��0v��"��iN3Ь��Ѝ�[Y�@MP8 �F�N��m��@w~3� �����P!:���&�xH�ye��������Կd t��/4�Sz	4k������K���9�eN���;m���!�kH1;L�T6�j�P�s��B��"�ДkD�Y�ގ�î�akD#>��x���O����S5]~Ny�L�0��j�������+���|,� ӶbڝˈQ7���Yn��kH�ƍ�yd%�0����o�멥7��;<v�W��Tu}�����4\�N1�<0�X��J
��"Wmc�\U��ݕe{�ثE;�e�1�ߠt���*ĵܼۇ��57)Yg�s!��	�g���T
�������i����)��ۓ{GbY�j0ͺ��wuf�wm�u<m�{Ĩ[z"*l�� B��?��	 Ȯ�(�ȩ�`�Q#��/�j�_
Nō��&7�L����,=#-�`�I��[Ls������q�V%�c�EҍK���`ާ�]��%��f$��<�҂DR˷B�
u���z��'��a��lzb��OGsY��Z=/>`V����"!�x����7��+:��U��|�a�cL�ݏ�A�
TE%�'�6��}��/7�9��G~��Mh�|V�xP;��h6�1_.��3��1���i�k<�B��c�
)��%�)��&�:�A���ԇ� j(�昹_M쵓�����>�@�_C�{
ld�,	3d�6���ib��ȫ�H.��n�7=sIk�r����[ޏ���|����a��Adx �\eW8��lD��UO�N�l�$��Dl�'d0��������dÕ��w� �f>E?�k?�|��c���}���6�j�<�<�]�;~��-�˲���\SD`��!u\��!`���z��0�f�D����=�TJ^��R��%������ý��y�*L��1I�Œ��P�$�����E�ZM��teA�\�X;����y�!����?����aoj�i�er�.��%TCe�ؓ�56�K�`;�W���/7L�,m;]��FJn=ǒnT|S���i�2��ьg�q�+����Ξ�Vm�ty��ξ�$���=b~霚�����r�~ÈW+J��S�(<�#�[#������oI�k��P�Nʋ��.�s^č��Ia�}b���hd�����"�׽
0�t��>Yk��P�Q�-���Lg%������'��!�a�&�I�՜8���P�dú�C�{t׏h��A�\�<^L��W���������ca�]�u���A�/�����*E�m:����et�-шLO�����)N���S�j[��*}���L:��/(,��r����ۑ (�|����\&��jܔ����vb%��?r���eNt�ga}�6�����H<�x1���|="��MOeM�8"B����E��ē#(�W������p�#��/�6a����i_�	�e�*ҼԢ�ܠ�N'm+$�Dq��"�43�e��Q@:��َma�Y�8���d��I��;Fi��9R��Zt5��Y� �R�6/�y�|��Ω�#`���;��	�D� l�!H�[|z�7y�:�8�1��l�<2����R�V������ڊ����k�����alR�Y&i��z��9��1���~n�t��8_�Ll���)j�\�\�,\����濈#>�a���>�dzW�b�� �m��4�x�����V}�M�uq��
⇣�㝫9s�Q@��l��AO�J�7�!�nR�|��03��J���)K+�a���!��v�A��{�Z�鄅:Nr��:[���y�����B�c`�o�)P`���]����9�H��t��\AU~'�W�ܳ�;��:ZhAٗK@8�ϖ;�ŁG��љ��(5��\�f6�}�fJ�w��+�%��5����3�����=��{T"f�ގ&h&l�\�0vw�o-e7�?�*�a�QuZ��DڎLcM�&$�.���v�|˔zqE��|6H��zÆK��L���Q�֛�ں��Fs�Eb��!L7F�Y���1.1aW������`�����d�P���(���-<l'�����킋�Q@kRe��X#K��N e�����!�#^������u���{q@?�<���rJ�
",�=������:��~WΤ���>�A��K���}�|�"��T�U��r�v���8`Z���MYՏe���Bz��|��a�9+dIv=�˲�#���N:��*�������!��L$TݹEa�a��e�i�J.&�1~`u#�����vu��,�EVՊZ�>rb3��=�!Z�ق{�9�כ��>�k�$;�K�RW����?�-������+�A�!�3L:��l������;er��g"�j�!5>!����A���l��6yV�!��$��a��Iɫ�j�(�k��}�d��8��d(���=ټ��u�'\T1-NZ����0k��~Rca�[��c��b��;�L=1t��0���wV�h<F�[C��u�X�|��>��F`�xi��y �k*��bqx��I�zr.��Zh��&�`)���N�r���Tmi�����NM��_��.��`�j���B}қ|�|�B4ؠy�S��� ��!��J��o�S-Z���Y������~X�O��	����,���ׁ�FE�=�D����C���Q�uD�A�\��o`~�媮��fq�����&87`(o/��P�@~plC8S�B;�4�p����a;m��*�ݦ�:��x!�!@	O�M{���E!��#0�Q�����:���Ƅ���9yH���MH�� /.��nQ�f��_�^ (V˲��Oy��АfBb��Ы�|Bk�2�QvXL�\���8�g7F HX���)Q����7E^�^��x6�%M�_��x�:�
yg�m�%0����J_��f��^�C�en��O,k<������ԝ�ys{Ij����W�
9�/Q�.Ź�̝Ġ,*��T �ZF�
k�:� �δ��ʃN�cE��w����mF��f��!a���&M��ȩ��zm^Z���B��1����lW;l�٦\�"i�<_>0tf�X.y�a�G<�36'_]$w��\|���B�p�I���e�=0a=,F=e��M�jKƫ�F�J����P�ST����K,�6��N��b�l�>��Wq�GG�;�8'���D�v���wu��i2�K�%�sb9��W^�S��gM���\���T�f��T8bv�[/�U	�����}7Un��Շ<O�K�(q�����;�� �2jѬ������\KyW�����3�!�T	���ٯ�|nf�N��*�s�PwA[���;�C�����}Z����;#/��A���!)�ӛ��!�"En��3eΑ�Ǌ� 1s�YP޺9�Rʣ|{�����_�ɰԱw����/˙�q8'�w�{�r�Êf��©�:x��CAF��,P�Ď�;��7�|�f�~�/`
/d�
'�I�z����p@�ء���P�z0�]�;n�L�Ϸ�!1�&����r͛��+i��64�=��.��t@Ȼ��d�@)���M-�JX �N�2�,s�pJ�9X&o�U�w�-�mz�΀3E�4�J��$@�0i)�� �7������d��YD�_��.�ۀ��,�D4�dvň��򸏄��9����O���Nɛ���2���hv�i�\�AD?gF�&t��;R�f�5���>���H���b��R����>�.u�;��G�ѡF�,|���c��D$��
�n1�ʐ�-dC:zT���y�Wl����	4e��\�0������B��ao.��z;z�D�c'�3��r>ƃa����xY���x�`Qt�e��X�L��ԇZ���/0P�)&������!!j"M�=��6X4������k!�T:4�Vgd�-Rԣg��NBJ����Ó���A�����0��w9�����Sp�����4�cwÿ�׺S�v��=;I{�F6�է�o�|;.翹�f����9����FHK��'���En��Q���p�ê��A�K�gU����{8�o�GZ.��trj�ߠ��.�w���=��A�s��ڇ��@i������ⶮ ��D��_U��"0p�����|cB��w��Z�]p�Nm\��hN�������q��3�C*kC�U�)t4�m�ҕ6V�����r�v�/�
P����#Х�mC� bq�j��f����y�p���ڠ�{�Q�@�q98��G-��X�,����-�q���*۸/�P�Sڨ�����P�vǫ7�i��t�����2	�l��B��k\����Ha��Ǒ��ޔ$<��Z�Bw���&�r�`"z��Gok�?�m�d��"��,�����nG6�,� g;CG��<�Qg�{Zs��k;���=����Q'�5PB[;Of�M�a��nʱ1Q��w�p�W9]�Lߓ7�����|�᫩�y.;�[��o����v�Y�.}"�A.���RRy�n]l0���H.l�$#U}CQL��w���P#2;e����n��z�CU>F0b��A)Լs� e��  :L���]��a1f62#R��:z��s��z��S]{���n+�� �d��=���3L��YJЩE�g���L���8� �[�Y�
m,ğ;.w"�5���N?�heY_�{ƿs�7��n�6����s�6���8v��R�t��L��*4��6�,}wr�+IB���!E8�`-��Oo,�V�<��~��/\O���9㑤2`~6��DH�֡��V���&�/�_������/�)A���|Q)���
��#BL�����;��#��@�e�W�v�$_�Y�(;�G3�ec��ܸ1��T�/?��Õ��o�(��S���Ə@�Ev�E8ԘE3ڔ���{���L�gy��png*pW$c�-�W�G���p|���Z8y������ <!ߴ��~t�����%+>F����'�>�:��1g����|�Xo��n	u�]2*�qn�˱�D�Y~n� x��������{|/Jj罦
��J��!�/��!��%�!�=ӊ����@�sG�S��Ƿ�a̲� ���S �l�
,��!e���kO��y��Mlߪ�K��=px��L��w�<�9U*�Q��r����#V��ǳ/д��$L�IF��F�_������ʤ���ܷ���E�m��.������t3�6��;.U��4,��h恠��ګ;GW'����~(���?��䊺`z��ꂡy:&F`{Q2�}!�g���k�I3�3�&����h�l���I4S n�e9�iZ��X=0f�J�$^ܵ��髐��|r�h)e����
;(�������K���j9r����.�.&=�S����3ۿ'�	���lG��`{j1�I��$�2d
�cA����{[�;�i����s�ӫ4�e�F`��Y��{Et�	�y	۷�������9h4!�A]�~��-�!��z�s�C���*�ϗ��kE�Gs��T `�����]� 0��FGVu8���?����D	���}�r�?q�u,�"��-�>Ơo��LI��Y={.I!F~�K�R�↖�d�ע��K�6��	��φ�6K�W��]g�]?��Я)`rx�R��F"���%��m�T^���!�k�����`�l�Ӎ�X5�(o*�읢�l��6-`�{
�G�^�k`�=�50��;�V�4�5p��'�l韙-;�S&�0Q���E�ܟʐyF��},}�bH�'��t� ��>;]^f�)���DFKd֧i���)��%k��4�W���Av$HUIC3���(j�ރ�hs	_w��)��h�1H���YA륱�|���'�u~�Ux�5�s�f�!)����N�ܟ-�o�NxX���W���#�D��LD�4�QQQ���y@��� �֐�z���)��A�r�}�[�����*{q���e�*�w��n2��N��5\���!�(R�x�I%=�Y'���.�5Ί����9����>/H�d�0��5��+������Lu�3����?^��8T!�%�Ҷ�T�$v��a" ����m�2e��Ո9ʐ.|��OX��e�^�3,�1_��P�NLI�[�T@[���s�<%v[5<q�x"s�#<d+jj��{���r��ŏ$m�J	�}iD�uϞ�:�Tx�j�H^P��V���/��;Η6���8sM�T7�h�V2N�p���[ɧ#JEtQ�sP��3;�O/w�E3�/s�G/������[m�P�4�$�z�?U�awa.*i�{�H�H~�9{�M�u����_Ξ*���ra-΃(A�p�����N���ۓݟ.ͤe�)��_��x�b�
����my����'(0/�<���^��er�k>�'���3�/��T�����,�� #��!pb	K�X��S��x��)Y�H�L�V����3��1/Ju�l\�R0��gh�o,�3H���ܤ�������P��^�G��t!�'�5�U��l�5�s�a��� ܒ������)��O��̍Cs�b�u*w�dY�#9c��Kx�q���I6Y2���Y�:�U���P@0���B��^)R�Q�*�^��+��$��g4�c�|ׇ��X��^2>�m�ļ
F����?�jC�hn۬Dx�xo�T(�}���8��	d㰀 �<�F���5^9�h���e�z�ńy�)Ic�`��u{}���F*�=I��f�_���:�g�*,:� ��&c�$@�-�5Kc�.z�H	yAYM۞&�ё]G^P�6�IN�S�+W�ԇ���j��#S@�����̃�:�7غ�F%�l9\�w�:y�������S���X���=L �r��@-ώ�o s�\L'd"��Q���EL��.Pm�, ���Q��'D��BE�X5�La!�u	H�J�EO-xy [�5��d��d����xEi,Q�x"��Ԍ���|൯�
$��fBD[ն$�ja���oV6/�9_Џn���@l��9s9��?���j�?�)iZ�l�5mt�Ra�������|��%�����썁^Ļ#����ˈO��y��힅8v���U8�р�DV��"�J�zՇpZ?�e_�����OK�����L��O%�%hyzB�.c6��q0L��p%�����a/[G��G\84�#jc��olg�6c��)\��.%��n\܃s���Ql���D�
8x��Tg�[�R@���vO[�X�� �s#�i�N�������.��-a�Z��`Y�	;q�m#���!-�~��®�#qB`����Gj�qe�B[W�/$����[|��r�Sո�}܊� ��Ntj�B�X�����p'$	�9����<�kYR��8�b2$V���Q��̎�.�T�o�����H��Q3��}��ɿ�o9�.g�<�\��KX���C:\M,�.z��)/�M�m��'eb�?��/Z��3�7
o��=��	-�>�H{�N�t'Ņ-P���_��$X;n�e�����}��l�����*�z�����"��Z��+�mꈔ���8��GF����z�4�}�L�Q�<T�/t�y������hJvp;D�#|��/�#E�D��*�Y1��AND4�d�qGG�7E��>�ڻV�s����tϓ��S�V�▨'?C5ќ[�B�4��f%DD��/.����,Ů7r1C7�$���bGL��/A��Li������H�|��H?F%]�i�R�2h)���{})~�e0ʁo�Wgr2ף��n�.7�["��H��֘�V=H2����Tߖ>ر�k����3��7����*����̏�~U����)��٧�L
&iU�6ܡʓ�/�0�n����
5y�&6 >#Q�\��Y��ϒ�����.�n[t�d��dEp�5ꨋA8�8}RB�g��!��[� �&� m��M������K���}�f�Ⱦ!��(dh$l0�B�,P8D��bfȎ:�������� N�=H���R��3Fpô"��G*� ENhy�/C�%q�Js��e����W�3̇G�����<		4�e��%�H�Lr��Y��_�SB��Q8�d�S��H�!+B#��u�t�K��D�N�Y�P\��.�;	ǋD�JژN�2�A�M8��Dm�@~#��A�.A��<�GHfVW9V=���oQ�X}鹇h9���p
�D^l|91f��E:V_ޜz��g�����/q�C�)k�o}��/�6g�=�� x[xBgʹ\+�Dz�c��!�b◱�>4;ZH���i�g�^4(�k��S6��`��7B��ɝ���U�;���)�O�`n5I�BR�ᮿ�T֋LF�Cb�[��p�����	|�ϭ�ba��
�-+���oEki|RwC<�ٟ#�U���͛d�_����H��#Д�nb���Ds��#%���_�XL��r\A�����8g y��|� ⳴� ��-� ��!v��ͅ���/��u�u�ͳ�HhTL&�h6�i��Ud<�n\Rm���B�k��
�=?���j}d��C;�����3�"5�LA=v�`�x���a�X<|��P@�\Q����4��?#/E�� 7w��)��ן��h�;Rn��7B�G�_)�S��������: ������_c���:�%S�M,��#���w-F��|���]t��&���Ȃ�ml#]0v��_mz�
�A_��&�L
Ѷ��'�C`��KQԴ��?<�Ni7�g�g��NZ%#%���VwoD�K�[���]w����D�y� �����'��t̞�,��B�j�Y�;��ĥ��*�li4(}OFsUC�cํGڒ2PJ�œ�W<9��ĕ���Ir	ѷ���^���̎>`�Ti���[*.۲ow��W�A�Xe�ԟ"���$�`�h*%&;Y�`�/!���h3Ź�wv4E?jRr��l\DΖcaH2m��)�y$�}瞘< ���Q0m"V�Z$���#����#*���L>b,xG톋�K�̶�����۴�"���ڛ�$$0�^��q����&b]�F��4�0����?2��A�Wc�1/>8�mQ^���I^��p?HQm���5��.�S����2��,�&t2�=GR@������p~v��Rj0�wx��rEMAB�PUS�'Y>_���`�,���GIQ0x*:����!?�q��ΐY���h�Fm2]ʝR�`�BPy��}ٕ�O
`����%ӎF�ƨ��$
�A7��8�7ܜ{��$4��I�g�!�H�u���27(��sy�&jx�Ϋ�_oj�V#�#Y�#�I���$�G��4]T+��l�D"Șu�r��6�}nE3bV�L�3�E���茖��>�xFeG��Ws'���q��9�bk+�:��9��id,/3;÷�\+�B'�$��o�Pb�w��-:���4:"�e�����/7(t��ա|+�Q�|�9�.I:Q<Z�<�r�g�HG�FVL@`���.br�4i���%�I�26�
K4-���X��6��FC�=���ڔIsg�z�rV9'���(9�25�疈J�=���Ȩ��럾�����}�*)�6e�]^y�LY�H<��[��Z��ɴ��Ǉ��"t�v��Dh��+��/ˊ���F;j�HT�K���a��p{$�U+K�����@�۽����;��3[�W�r��nK'^����8w���6cR9	��ػ��C�g����+���wq�����nG�un%�@վd%Y�6�0�����ƽd���q�b���*ʧ��W͟��Ε���+;ӏ
�s�M���)L�3����"��ø8�@��V?\���U:a]`+��R�n�b�f��)���Bbt�j0����~K���Rp����:�	�\j��Yg�=�	�g��f�E�Rw6���k
b�Ç���Έ��GlN0��&a)���"}ưZ��9)�y�ʕK��_����Pa�� �DN� o%���?�={�����9i��r��I�Ӊ!��ƍکnGZI��~y��xl| �M&��7a�ؔ�C�, ��u�y�j�N�|���g�}6(r2-5s�]��=i�v<�!�@]��yd��Z��[�ӛ����
����3��#�I������O�@��Q�)��t-�zW�c��:X��z����ˁ�pj�ܣ����y�.]r#fw��uXR��z�S2T��˰J�Ӹ۬�]���>dp�V�����c[;w"W�)���R��sq�z�z|eW��Fx����Ԙ��6�ʏ�s:�ɸk����~�H2���d `p�Y��.�뤦��DIBj����-ո�$>߲^J������Ċ��i����tʖ����U7k��f�
gnF*�F0W�fE� �Fw�����(�6=&E�<�zm�:��`p׺�r�8z�@���2|M+}���J��t����CV{���OP�MX�|xv�Q���䐹�^���ӻMQ�$W�e�A<�,���pj/|���焞Y���̍u�-�¿
k-9"��Ӄ|�����u�uGpP��� ����B=�s�;#���<�ac�Oce�����]Q��N=���
(t��/��o��Ű?G+ ����N^n��3�p��i��C�9'�j��i]�!̍����K(��-��X�.�ؖ}���O&�+xM n�I���0}�{���n�zG�A��)h,H����n3�f<�Ⱥt�V��?ˊ�&i�-�N�����@�Y���Yj�_N×�r��f�1�m[L燇�ɷ�5����\�E��j\��X�d&�J)��Ü~�x�����c���B�	OD��&����O%�{UH�W�uM@���<a���  �*�|N���~��"��r����w���fG"E#�q�3g��A�|�ո�A���G��\\����BB��"�ʒm`��c[�"�|,㕪�gMo�8ٮ�J�F��\%�	�!��.;���Ϸ���߉�� ��8�jq�І������o����r��Y��2u��eHS�+q�xW%�~P�ɣ�Ww)�S�n���ݒP�N�����^�5D�q:2tuC	Wȃ����G�o�
�_;HX�ǦS��� Qg���&k���V�%]틭{�|g K u�J��J�@���C�s����E$�$��r�-�R�v�+=�+{-a,�c�&�����,�'DF$�9N�DS�]�o��K��JH�Yݾ��FH��'��WK)Bt骪�u�z̟����^�3�$�v�F�QA������[N��h0���$p�@;�!�"�<��r�t�Q�q^�1BB�L}�ʂ�>�m�t0�DO7X���tg&�Mo7̽yx@<[�Ƭ2�]Eڍ�
h.Qw��`S�t�9F�����ۖ!������&��`��3�&���ܝ;��	�g�t�
����t�?����A����r}����*"O	����$���DA�_�aj�tW��3{��4�����"O¥���T�Y�$��G�dj��U� �wx'��r_�uaժ
���_�O�;�ZA�r��ũ1�DI�՞���'tύ="ӷ��$����Z�K�*��:)�|+�E��/�uI��rs����cL-���!���Dݬ����WX�`��ې06O�ǔ��� ["��&���v�c�!9���;>�@Vz�)	��i�w��}��}/P �&�oϾ�-YǛ�Ԛ*�/�>���h��=S/�g�Z�!I��l�#42qXTO>dχ�k����B�&Anf��^���z�i�4�r �X��6�o#9��G��h��|y�Q$����up��LBܤ�ۤ���ruc�
�Qч��8��ᢰ&㫊���h�%�!Dk?f��D��Ӷ�+`��c��*�'c���7Q��Ҭ��^�k5��𖴬��U svg8U&�n��R23F���5�����V��[@2V���,f4M��7B�H5݇��'7R��>�W���� *'�Vf�M`�>����q %���}5`��7C�@��vR�h���s��,������:��H���� Q�E﹋��;��7�*"��-\���N��d����s�P������)�v>6+�ǆ b���ieȶ	��د�0�e�jǫ�C��ۑ[�K��`�c����l��镒�w��������~4od"�,�]j�l�����~��uXaG\�U!�������d�`�(r�K�m����Q��=s<&��_Y�l86gRx�P�|���1��o�޲��>8PC�`���TA0���o,��4*`����W��#���H'F��WZ�L�E����}q�.�Hc&;*��Py��V0ZN�[})����kC��c�G����%ƍ���;m�D4���0��X�m�q��EU:�.���Y��U������G��9s[/0���ji ��߿��M��MwP�$	z�X(���N��_�%L�����°S������'a�k�h�j���+z��OG��d�5+ -nZ���L�K�dJ�+����L�!b�����UO��� ����9}�M�M��N����ׯ�d"�ے�ͤ�`x,֓h��^3$�B�Z[�FJ� :D����w\��5����C�U�i?#<��Q�i�[o(r�|r�p:�?��7d�v ? beɽ��"���VS��5]#��P�#�P���s뙻.����
T�I���+��3 �Z�9'QP[Z�3{�,��v- <X/q�^$�ٌ���A \l+��h�т �E Hr⌛�qaC j����n�0DkuD���)�E��'��b��-1;���D߻=��d��s��X4�6��f�����i}i+�]��u�c���!���Acps�P���|�	��m �?O��7�a.M��S�
6ܴ�V�o��d����E�3q��3+6t`P����K|F���M�w0������ܼ
}��~���YI��l��|=�O���cA��5ճ�<�-2�i��p՚�c�:��D�ta�@�y.��5��=�%a�J%��ۈ/�Ur2������m���l����d}���9�U��Oj�>|����ݹ��ܾ���0:�����eF�>��>I�xx��Ɋ!�k�1��^�{)Q�J5�%Y%���})�a�}-]�=q�s���	��e��uܷ�f]JiL�MB<VG�D�@���<�B���a��Gfn0A�w0�P��"2CwlVh$u�E�8�@Ǔڴ��%�j/�trT�F͜��7�����7����c���B),C�^����B��4�W�"�X�������X+#U�����R'H��|zp+WRRO�^PX�X}]��|�C5k��.�
+�O�����$�a��%=i5�t'��r�#��@ƒh��l���N����ΐ���Hj�D��Q��I�c�@D�!7rB�W� u�	r�����8�-�V�Ȍc��Y��jb]����(m���{��qF�ԏZe#PB�e#�gk�Yj�d�̴�����Nz��k��,c�;�I�� 5�d�y9t6�?dØRb�uT����ȯT:��_�fЃ�)#ͥ�D��<
3���{����Q� �PP�Zg�S^��X'&�p��H�:_����B�\I�ݮ`�9���	��F�s����OR�U�EY�)�zPt|�!d�_Sں��y��u����M`��~�?��_MF�C<~h.#u>�w�j�xrj��~��{��Y���J�C�<�X�C��G zH��p�p�1�݉�*�z؉���|��B	�"%;M��F�������Dn�������+��=�^��{�g�� M����TÍ��u��N�!l��"O,I{�F
!{���^��ʘk�UO<��N�Ȧ��M+��yK��q���06�(Ш��ױ����2�S s�bY0�Z�W���f�No$%� �����bQ(6t,��}�ʹy�tl�-���yߪ�q5�D-�R��v�@�2��ޙ�N>t����y��)0�	���9�f>�j��Z�G۷#����/Lf�I�n@i L�/ߧ�� �72f0#�y���30��B�k�f�J���Պ�Ws���H�]{)uU��C5�����'̈��1&U��{Ė,%��~��y���wH1%y�r�	?䪐I��#	?5T�������C�I�m�v��2
Vԣj��'j�V,�&�JW�߻�q}�)ɺ�ݖ���Ӽl��\���ӀX��5�x/���L=2�+�	�U�1u{�H�V�B�G	Vί�V�;�� �@Qz��
��jjMkL(���	��q�n��C4��
�f������@��Q�5?-����_��������
��mu0L{�_�rp�8or�*�<�x�
E�k>YkNq��J�0'�,J����z��R����&i���b�������Kc��!�}�����@&���~�O���jz��y�m���<j�J�ܺw��
��k�vH!]U��oՁ�_���ω�qZ<���>۽~���j���y��0��@l�z�%���a�f��gԨ�L��wத�Qu��'|;��25W�i�cK�gx�iņ7�V句�)>d<l�0�Q����U;`���6��� -�����L����K?���=����)��.��s6e��ѹ1B���q� Vb��L�u�y߭��I*��֫�l���D�<#Up����afT�E��� ��Z�;�3Cz�tlky�҅l5���&�;������nϽ2���o��5��ы~#�Hn�+6���f��8�*죖��9�6��fɮ1����ө�?38,ٽh�7ay'��WtCʆ�MaQ���U�9(o6���~�kuu��*#��������ٸƬJl���9�� v1��1>eF�BY�M�2��� �ns��Tsqw�_˪�zKGpdo�	]Dc�e��t`z����9�S�)PE��*��I���]��@���z(Nû�W��D����ʊ3���˕k|S��'�ek�9ZH�Y�稭�<}��F��K(������������W'��b�g���*�w��e`�9�\�D(��P�0�R��p�H���ܖAe��}�\����4}6m���n��b��Ȱ=��}_��BM_�o�n����n���%.��CΒ�K�!�jHF�|XߕT*.�w��,�?i�9���Ґ�z*,�����c���|%����H7vJ�<�N"�8��Q�ʾ�k>4:CY�c�x*ֿ0�a�"�%ڽ!yJT��S�f�M�b��M��)����()}}�f忙�����h�n��B
���	6}�����	���孽�����r�`���	����������F��6<ꭡ�$|K)-�eBO$�!3@�x�o��~F��_g����h�ǝ�*���-��L)��TI�Ȯ��E���������;C�(��E�
��B��S;'�]��*��S
�7��?=o�"����% .F�m������d�sCB�8�=bƗ�EC� �8��^������ۘ׿~ݛգf� ���>�ea��F7{���F��Z&8ޯ�w܌ck�_��MOW��m�;)�����O���E�)�Q���m�q<���5��-��2�AT�B(�Z�:TT}�h_�R�!u~ٻ�Q��{�HX嬆l
RO���ʖ����lh/5a#y�d��X�A=B�I����}�N��a���#"��'>���(��0�a��)j�'O�ʮ�z�	��h�5�V��\�^>T����J�Q�:�y�~�+�A���-��� O��o�9A��E�?�y�i^�E~S����.��������׌ή0.̔��R��
�B7�H��[+�7��oN�5�q�D4��M)-$���H�x#b�Q�־�`f�E�V���n�e�"ہ�J���u��0ڡp&�Y��R]	[A|:E�|c�%�&�t'�!V]a5�?�m��G�*�g)��!�s
u��	O���=?���w��%%�M��p�!=p��*�YI8�F�QT���spI�Y[��H��pV^��f��M�I�+(u|�G�r䮢]��mDg��������Q���H���b'K�uL\
)Z�j�l+��!�Xk.93���?�L��xQ?}V"�E�������z����H�~|���sIӼ4R_:��C���������'P.p�����F-U���ﶹ�֣�c��
=?7O^hQ���!�����лt�d`v�񰐆MM8i������MB��{��*ه�_
h��p�H�2�eY�)��Yf��ݭDG�%��E6T(�F�)���o�!:��mA��̾O��_W���[����x�2����zT�UmՎ�^n}|�*D�qmS�$%�~��F0���ɑ��Sv܃f�B}���n
6t�3�<B�}<�m�F�l��qU��b{�*�wd�\�E0�Mv��>^|t���Ҽ(�����3�3��U�H��N,�K:U~z�(��?���C��,��lʰQ$�v��}JT~i��}�x#K�!��{)��E&x��.�F�Dk�bް'��)�? 	�������Q��"� ����D1�^���(n��!�}����$��o�ah`�'t�:?Ao�}�qѺ���@
�t�D��D,�c���}�76FA<tئ�;"�I�pY��X\���N�h���jx{��ݯVg�z$���pB(6�>����d��ָ0[����z\*Ct۾@�n>���~xI	�Z�Ʊf�ot8�%�pN��<���[9������IT�GgW:�T�	t	'��#��na���y�K�4c��J�gӸ sj�Q�.@���$�&��k��'������I.D����+э���t�8F%p?�bIa=^���w~]���v��oi�7��fZ���u.h�6n#�|e���9&� W�&^��g�v<��9Q�[>G{�R�T0�R!�E���-�P����4ђ�Ln ��-�
��
����AQ����}����5�(�F°�����@��M��|*PP�1�S��`�s����p��< ����$���X�&+�uؾ�>Ʈr��cw*�̀��F�me���~������ �nG!W�&�,8�?� ��4���*�ܐ��3��=�`�4CN�o\V!���������$D���=��}t���Ւ|^Ti,�g�5�Fsx)ؾ��)�߰�!��7޷�����jg�����6Dԛ�>�^����𩞃�������l.h�����I�U�n��}3g��-�^�,ք��u<X�$-s1\t��eZ��8����$�o~�:�Фa����t���[�M��_9C�J���χ:��%�A{�����z����L,�E/������kd���Zm!1?��.Q���dqA�2�G��vX�9:9b���]�W���$*́	I���Ju~���h�@��;�/�����)���T����Z��di��C��S��J�a�3���C�0�/� o�h��>s�ɹE�C�-*N���"�G3Ap�&�-hb���?,��-��EHI
����(k/�dSK>�փf�Vt�Ut@S��h\�D�
|@�h�]�+��C��|��	��v�s��Ɓ2���Y.`˜:��!}<BlZ�������9��#^�^;#'�;J�~�	^C�Df��6XQ7�j��m�;1����B�[R����{�Ĺ !X��ƌ���n�Z��	48���^rF��/`��T�E��ކ��ңH��Ik�|�x$�Ly�2���=���:u����H�JW�a��u�<���b�b���\�wn岧�!uͭ1-`�0 �2��L�	��k5��*%1��/��_��]o0z�t'��@T�ˢq�t��j��<�6��qz{�H�k����0�4�m��T�B�����i�띧��2R�C��`�o�#5ӗ���ـ���v�&R��F2����1���?��N�������* ��EQ�eJ>"�`_�^j�ޮN�9���9(�?H�)ި35�`�4�#kK^p�� L��94�ZD����z"�h�-��߀�*ﴄ�+�����J�w���@�Y��c��})i�x�H�nH���>���m�z�
���j͹�}t�������ʯ4���@���L����|���S��JXV"
1�U��+���N��Ɓ�����oyȠ�NT 9�Ln<\ҐO"TpI}����m��lr����u��(����o;�9�tW�_OQ�{�0�N֖r�V��;��o�&@�ME����ʤ���L���5�F�Eq�뭫��Q��c����5�/-���@˝R?5O�.R��N� )��U��>���+�����?�B�->�G�{�N C�TѷE��{���3}^k�����>4��JH&���|>ф&Ag��y���o����?g��	�Jz��[6�Wn�tX��5Nh���/͕���9F���o��`_
�����\rz�ά�*Hs��0�S�h�H�P�	:L��!��f�W��zCFF3;�ܢ�I�`��>�hz�2(K@�;m��
.K�Bm��^
�kģ*�vb���R��o�9WG5?�/r���=�²#�3{���O��+ 	� ���2[1�v�8�un&͐�
a�󘤃$6�/�_L3�,ĖU��S�^+�d�^�2�)%x�l�� �`z
�C�vy��Ҹ��zìi��e�U�<�^�k������l�]�o�*V�2�&�t ��P܁n.��VLp��ơ@(Ǎ�R�A�û�EꎣϢլG�&i%J �@b�U�_)��l�d�̡���L�,���P��U��qz�Ð���S�L�g)�K��{r�m���\���,�1�zʛ�h�@� ���!;�������{~Q�O��!ߩ�%C��i�^����<��b�h�(C�$de�N��B�Y��S_�pR�5w{�G�֝9��u�TX��9������Q�=3v;FhW�Z��9��,�5��Q��(w��f�D��4W�2�1;��! ��:�fO���Qʦ�� ��_�@�ŨU�w�Y��zk����֪���������'�a*��M�N�� �NZY�pu�B���~�4�m>[��!����f���iN���?�a��/�B��`��W2��QXo����,}d�K.è�U( �/�9�<����\e<,n��o껯��� ).RIPn�i���Y7=��e�wU�G�W���
5GıaA���T���8�U�=v��O��[��?��cG�-]�+!ₗ+%`*�.B��)�6��u|%]Q�*�<UF�F��u��IV�&:�^fb���;�]iK_��E�C~���g;e�o%բ�%�+���_�	 �&8U��~��_�x����;8�N0G	PX�L͆�VQ޳X��ό�e󶈔.b[8u��a�A�Ķ����c}T^0	�$�q �d���y�ӫή� ��g��'^��#�S�Z��{��� ,ex�f�E�*��-�B�N�_%灲����"��^�b�d��������"�I��+��2�*�Y#+�vz?鞣8Ǟ��GwQ[D�t1��PW�P�b��X�K�=�������伷�3��vܒh�W����}�?}8z���}�r��/��\�M��S�Fv�tD|�қ:Z8$8����\�����o��������&���L\	�|P�;����<b�`4u�2�Cd�"��h �'�[��m��]<'������$�)�^�ʴ�c�kf~�W���̲�M�iCP$�����w�0�6�8D#;� f���z��o���Uյz�6[l�Aw�~�6�W�|*��4��s���	�U�,nu��m�J`��v��o3�@{����TV�l*�P��8�Kԗ��`L$�y�8m��F[ְ��y%�2���^����������3p4��%��)UPy�������eb�8��z1.�Y�����!�l����Ȉ"7��������:[���If�h��L�Fk��S3<�0�As��W1��Gûʣk�\jar�S{1�E͓ ��ı���D[���7x������7k.H� ���b1��v&L�g/
iW�n��XL�]�����>	�>��:n N`��b`p����룠*)l�0�+B�K.��A��d^E����C�:�|�N4	 ��39;&?)'
�����u<��'t�F=�jI������^�ۢ�!.���=l�2�ϧ$d(�jp��Ɩ�c�I��4��"g��q�
���2�Ш�o��ӛl��|Gt����'B�8��b}>���̂��$��%�*�e�k��$��_^�C���=��2�]�� ��-S�2����8��v'�+�2����T�X�=�W\X{ �C�˴1�hD��@��i����t�eqJ���H"�br��F,��m��6o������T��I�x��\��m�і��@&����ѲU�~�pk�;���z���;s���A�a��F�Zgv���t�8@�}Y9*�vrN�7��������Q2;I�gbI���)Qj�iv^N�������Oo��|]�X��;2��ؾ��lN	K`��|M��:
���0��Q�k��0�2��ݡMM��F���.6]�*�kZ�^o������F��S�`"�#Q�O����{��u+�fo�s�!���:���L|K����# {�k�C��j�WQ��y�}��rr.q���� {��-V��#����3 ~4�j�{��깽��)�^�l�c�(��P����z]��M�s�.�����BwyHec�Ō4�����Qf W����tt5y~W�O)uzq���x@�[���5辧y��θ��d{j����i&��ɟɶ�Y���o)s�YhK���+�ڍ���K�_��.K��t0 ����1�q��&�8�JS5��%B��NP���ʋ[���QO�S=�����?� �.�8%b��1i�Ĵ �����T�*��+�:�^_�EɊ��Y�ӜPc�(1�[B�j���{�7�SZB�A!;1#5���N�X�0� �S��� �z�
�Oݛ�1��b']@P%���(�����CN�&m�u\��"�6�LL�;K��*�����������d���)$�3H������gn�t�*��ȀԦ!������B�$k�N`/�v�S	�z�&KI3�Е"[��P|>��.�5Q^$j��tcLOI�?{�M K���$��z����q/C���>c*>
����b�FIe)1���J>}����4D��F�i�y����p)QV��5�9�)�0 ��G[i�g�����i݊�t:zS��}��N�����W*D�y&i5�z�E�W�\�}��]�+F�6��@�����'��_�y�����L�q+��wV���Q�V�S����IMN���{�<��cM��sp�)�"Zt���;ۡ5d��V�dￏ�^N����\�N
�H��N]Y�г9�W�q
8����2wMi�H�\ED�����&?�F�[*��o�_~�l귄���͸��N^{Ac����a}]_�J�P��4����I�3�{�vI7�!�z-G!���.��n��lX]c�24g�8���,<w�C�M�w��k W��f�F�XA�O����Vw��Y8���NK9k
Z<X�Gc�Ч1A~)��3Y1me\%y�vt�4P���6���
��0-{�_��և0h|*�Ƅ���E�w��HÇW:���&�)&�7Q6�R������t�8�3y+��~��	��Lvf@��x�1��T;��"�0�	a��Ī3mB�O�cz�{b��+��D?��
����L��c���B�	���ʵ�� eTm�|����3_^�ش/�]�Tיִ�����e�ȩ?�]b��y��� Щ!+D��|>�����wϮ��yu��q��X��$�ᡬ��ȭ�F�`�O��~]w�x��Z���1�3N�V��/�oX)ؒ�4����#�XC��18�'�,���G�벤'{�q =�o�u"�.�M�2�ľ�D�5���E-��Ux�]i�2K��}���$,�愤Qq���]�J���2����1��W�A|�Z��F��H*L�<rD'錇�_Yp޶%��	�5�;� �rwc@�(���@HX��%s�d
�g�Z;ﻙ�x$+;&՟�h��P��y�)SiV��
C�w4�:�5&��pC�t��.���?$�T+S�$����+���w��NNA6f�ƙ��/�sN�:��1h��h�����>!葧O����c�z"����"�ҥy�J�H����� �{S*<P	�w�7Pq��Y�}�=c����&eȯ ���\�r+Fs��+d����jW1H���k7�5�R��Χk�q~����F�������ҍ)���>n�0<Y�4�&ծnZY	R���%u�)e�1i�b*���hҦi�Jj�p�&`Ȥو�1�_��K2J�Oݹ�O�n�A���#ŵ1M%�$�E���ޮg��*Y� ��"�.�>a�@��D���?�b�*��G� D�X�\���7���wy4i''�l���/�5u3��=�Q\���	&��H;��.��Ǐ�?�*��D�R�|�ql���r�Iu2"���l�C�Z�<��Gf=S�)�Qn=lGǌ��+�jQ�2ǦCD<U�ڞ=�F)kl��}�~��8���덼������ᯠy��9f���� �����a�r`���̇-U�>Rs;#�{kR4��A$��x%\J�iI�6�Z,7Q,&<��"�P��B�ӫ���/�;�`�10�=۰�?�9U��O+ H[���? ��pc�2X�Nf7�m�;m��}BL
N��^XҢ�c�> �MD���XP8�,�|�|�hBE��q%�d� �B|)��@����4G�x���V�0���X	gDI��_�9���.��3ё(WJ_��z��$z��0�IҢ�.��sMS�#0N�� �z�b�QlO[F��!Nu��
�I��E��-��is�s�;d�$Cl��2���hLB�R�2$D�Fk����S5!��*O��C����-.��$�Jd�?���4 ܟ�k5ƞ�!}�>&i;������i	|��p�~?�_\����[�P���j��_;}?�D��*NAB�6K�z&�/WߧF"u��~b]8aZ4�ה���6#���ˤJ\�eYd69��ҍ���T�&�w�g^��'�{������W�1���P�pܝ��`�)�d���OD�}CDf�Wmf��L���á�?���
/�{�Z>hZ�^�SQ@� q��7����FI�?��&�FR����6wm�e�@�zLB"=X:�!2�ڥ]�o�D��S�y�veH�,���	}Lz�/���
��j,��fN�����9X�����3f<� ��ӫihQH��~��y���6̥G�y��>�+�R�Jw��V�hv�fѧ���:����y-R��nB�]���`R�(����$��~�η�o�����B+���^���߫��"�������;7'	H���X�n���T�5^��^�A�l,�|s�	|��Y�����)�' 4Y�b֛��,��E��YBF�)�
����&�+��v,�΁D+a���8�������8�����Yt�m�W���s+cw��Q�rN�(����bl���6��̑�5��]4���-�9�~�=I�A�?z���I��g�\$RC��o<�k�tP��u��Q������ף��c���^V��&��w�P@=5Ǉ��ɴ�l���R���!�Ҝ�89U��!�P��ς�3Q5s!5[ b��	�oi��#�� ��"�q�әz?�A	{��qYMWU��ʘ-��=���w���3�Q�~�*��+)A�:ڠ㰀�8�؛��Z�>C������&/*����A�` �R����1��!M�ZFc$��LP����<��RB��1q8\Yܩe��N9�e$�f()���B3�
�ҁ�PK�-�~-g�RY0J#:�I��p��?F??�A~����
w��S$(XJ�M�8��ɱw%>��K8�:�E�BjTZ��9P=��&��Փ��S�m�eT���&Y��-2�:�
vHff���%��|l���y������1�I��i��g30TH9�&(����:[������F�!l�Mj�b��p�	<�
�]��*���}��8ѹ�ǞL\e���1�ؑ�ep�Q�S|����.<h�"��~\�PKUVb���EA�����(��?,>ϗE�;���=<��5���	|'P��_/�'���BC�F"��fH���Ԫ��My��ʚ# �YZ�w�j5��|I��I�	�2�O�ut��^����$��C�������B/h��r�����|!\}�9[���wzBF���W���}쯓���k�i�7l��� J�	��y�%~�B����a}�Q>�4Ӛ����Y5��xmS���`s�O[H��^�����k0�����N�'�M�8R�dO�"&9�w1��C5��gf���(�{��Y��	v\Cѵ�0�����}���(�CF
�?�x����#	*wL��2���R�ZS��s*}J�a��L����z��Q�&�l���=�Kd���9:��k��U����|�(XR���f��t��J)&�_*k���os}Gp�.1�v����ؔL���{���>�X���;�^6~r�Jck�79p����־��d�w�vZ����m�2������Es, {g�H�!� �NIד�o5��y�Җ.���H�=�W�iY�d�	鮁6��2���oOOa�P����Z����y�4]9b(z3���\NW䕔��Yh��{��Z�孛�� ��͛C �ڪ��M��n�tU&l����R�e�c���-�Sܦ�r��7��;��/�w7�v,ƹ	j�i�r�t�K�+ﲿ<7փ(�H_v?�:�A:��V�+:��!p=R�_?����)�2�����	�c��'6_�1f���x�]]>�L{I1:XM�Ϝ��
�Qɼ�-Q>u��O�q���iL��d�(a�`�[T��¾��ݩT��Ѻw��~ݟ��A[}f��� ��-ӌ��" a��S ��c�9L�=F]X�|���Q���\Ŷ�]g��luĹ��[� aA:�2�o�2O����k�*6X׻�Ni�,ш�4&X��gؤ�O�8��"-}��b�B癡��U��r�H�~�̵���(���GS
��z	�g�yϻ�>̓s1�nX�����bؓ��N'�s�A�L+�שּs{vq��YF��v�q�b_���hަ�R�Ƹ��B�x#�F�>ˀd)�{6F.	����P5&ܼ{pNv��4�ܶ"�Z�'��7{*���LW��r:Vg��ߦ:��۩�����WOcB��0+ǧ�$5�J�y&Ua�T�Z ���K&%��sl���:'�#����D��E��P�س��
�*洟����S]@t��^�B��6�&��Ԥ��<�i��>҆��+h�?�����%�^�%�)�����r{{o�9 �l[��&�IYo�ᤗS:�C�n�7����N���!�R���t�
A �Ͷ������"?�B�~?��<���7c�#t<��)����Mx�^�%~��,�8�j�]�=��\:}���@��� 9��'�e� H�d�p���Ue�q�5���t���87$}i�s.�ԑ���-E"jKx�QZ��)F�����P�X�����"{�^�:�Icr�&3Σ����3�Ċ��o�3��������r�5� ?��H�>��q�^7�"E�gOh�` Z�r� ��冕�R��T�J�eG6j�Lꚥ>n/�~��2��+e����lNZ9�)��=�$%����S�Ex{J���74����꿠nO�I�&�;R
v_队�����.���$�-��E��I��4�uU?4�Yyb�Ѐ�"�z��y��arˎ��\}��uN��Ȑ7c@�6�P���)��5����rI\��L��l[�[8�}��Q�s%_�jO:`���l}��e��AΠX��o�_=7m|Ł��(WTZ�ҢrB�h����n�o���s��4�o�S�� P���x߭N��_/�BE�9SK+_>�ǀ@�Y[��Ν�A���1g��VR>�b=�4���x���FY\�)aـ�ן��!%���	e���'x��@M����F7��H����ÇD^tj{�����~)yDە�K�k��R�8� T/�Q,��*��� RB��_�i�_eVa�ڡ���&�e�k9�T�b�C�~�k�%���'|}yԑQ`E��1:��05������a�4��Z.ǲQ�Ti2���u�����w�Q(����fhK�в������;! ��"{��Ŕ�`[Ĩ�f������wؿA2�h�c�q��P�l�R���NM���.�K��m;r�	�~�+�O��%s��,A���h�q����qr�|ɺ{g�@��.�hp?g�nY�xZ8r֎]?WA�n�lR�o�lR, �uF��ڝU���΄�'XA���k ;k�`lX��z}\�9�v�9p����L�7p���TKFyw)�b2���	o^߯z_�-t��5��\���4W�{JT��%h�.PT��������9fhߞ���s�[q݉���}I��gF��*v�-������Y��iz�1�_kw���n����	�V���(�b"��8 ̭�N�'v	VC|Ѯ]�/[F� $�>�I�;S��)[ѩ��eF]}UÜ��G]%O��q���O]^�S>m�Z�:��$�I��V���u�}�[���|�������}�)Pev{�;H�.�����UF[�݌�#���(<)X�A�b����^�$M]¿	��n��$Җ1�a�ʐH�x�Cɀ4��ԧ��cP&��@T��)=�21+|�P&��|B����߉�̲�P/��sd��2�y�'�li<�q�:v98���	�s�S�_O��8��h{F�.H ��of��`6|F�u�B�1���1/����s��h&�\V�)��$�����wh�D�NW�F�r������ٺ�)k�ċ�u �ExZ"��"�7E��Fd_���٪�ʘ� �&�e��5���Y�+�[���F:�	���k>t܌X���� E�=�@���3��7���\���!��\oy ��M��<c�b�_Yl��u����n��&�C��'�㠝��d9�@�zG��2��¾���8�`B�6��P�7!��C�����Q�q�L\�T�|yE�x��P�����X�ͬ�~A�Ms���rLY�8�T�}��
b�^y�)���}W���6"'����?n�֝�?����.�0�	�A�,�������<������dm�*EB�u^\9��.���(�9|][o��lxO͇^�$�ӷzxT��K��IT�{�ò���S��gVOp���0�:i�ﾤ�X�(`Dƛ�����㽦�@�
���	Fr��*k�(=� 3��:^\؈�L�c����$Z�sg���{Y�?��z��P��y�V�`����[
l�Ѓ�M#��T1��(n����)gw.Z1�X,��3�+É%#�1�tOA4d �+��P�1m��g�`h��6�L��1��5O����m�zf�x&��9ۑ���*�/�&B|���JW��[G��G���AV����o�z�w�C3�,�����$�y�����Z@�fX�_���ܮ�U��F[We���������$�����i���LK����@y�2��;qԍ�eɘ�a=�u�GI`�=$���qe�S�� ��$>��l�刨�T|#�)��~���r�C���2&2O�/mG�̍_���?����FC,��zzw:3�95eZ:�.5VP����L9�x��)?6aƤ�J���o�9נP^�M]-PPB�#X^�Z�zb���g�+%�0?���K���J�;�������Q�O����5��V�f4D�_��F"z1#9���:�2�ln,�0�1Ij��@}d�;b��Мx����O+�4����C��ߋ�UT��IF<N�`�y��'��N�{o�Hޭ�s"�B�A��d�P<���{ǒc���ncq~zG��!N�g	�25�ٯ�|�u�R���\��e����,/���f��'���F�ҋ ��dP�~t���ĽQ��#���w�SA�Q͈8�A��P7�2f@����c*$	D�T���t��i��5�ކ#�c{*j���~�ýl �a�i�X�W����c�9]�3�?�.�l�w�V�K��M���f	'*D`P�Y�!!�V�pk"���C��� ��C���"���V�%��#^a~�Jh�?�i�}�~!<��j���؁�iC
�eB��P:��W4�c3ȁ�F�v4r����Ź�D8���aX����,��Ǟ��s|��]�H+���A�b"ʱK�V ��
���3E����y�~':��7��	s���sG��D\ɮv��5�c��U�F�5��(2T�<���+��%��Ǥz~$_R�길��PlA��%�C�� q�,����9�:�����U@~K�gL�w�<�%IƹR�XR�93��L�E����Kdk���!� �J�(�v_��N�/��m����p����~�f@ۀ����R���� �����©gr�ԛ�!-b���q�/.� Y��̈p���"���z�l��*:%m�A���O���QW�'�QT�r�=ǘ����}��l��٬%���_|����i��n&$�s�$�C/ԝ3��ԋ���iWYK+ϵ+p��*-CB�N֧�l�q�.��P�����������n��Dy��T��E?-u�jg����G	�|e����Vߏ�Od����B��s���܉�3��#�1��<3��(
@��I��9#W�5�[m�˃���O i�$Ly�� +~�ͦ�D��) oo�`ΏFd��ɸ� ��F�Ɵt�1V�3Ѯ�9���>��U�&|5xk�B�uʲ�+��vB�G� �'D863?�V�s�_��-��r�\�D �$�e_��E�Z�wd	#9/��ɯsᏗ� pԅ�G����
�;����'��c~h�[
e\��ʸ���64b����
P�i�%;yI�v����#�a%bh�!�j�8y4����3��Û���%������f�ٍ�ӏ`w'��=IY�:��76\s�.4�<-.C�!�j�I�G���P�R-t1>\�G8�h�j�ᣰ~Y�L�	��`��y�1j���E�?�֞t7�a�c���G��W%��-��YW�M&����3p��j	���G+�'JxZg��K����Xϖ���(�ANEZ����iwyEA6w��֯���jCS>s��cUQ�0���l���޲�*���������*BӠ�D���-u���B�N�Q�g�=m]����I-Q�|ۗV��-����=Q���꜐9�����|�*��Y]��܆1*��2�9�Uw�rN\��DM�[5��c�T��RQ�?�f��mBY����GZ�ۮ#�����פ"�/M�f�J�~��]��>0wD
]Y����M�O ��7���
}��L��U/��}��@>9LY�ZZq� �?���8!k�� ����^ᶶ_��*8 D�"b`��������~��c���4]���F\-Ѣ9
Z�񻻙o�c�>�ƈ�,$��]���%2n��Jț�I��hfc�p���i�!@�-�*�IF�нF�?Vk ��[���R.��B� �`)�@�����]�l���u�QW�&�|��G�U��TI����,���0C�K*4|v	wCx�Hݼ��!R�3'#w^�Bh)A7�	���9���Lb�M�:3e ��0$���p��_M��o~UR���� Nm���>M&�ۤr��괙K����v$�
��H�6hP_�z[G��0���%�FSa�
L�Tf�F-h�UrEJ3�)����j��X�-~��?����6aE�)ە-\��,���*/��ֳ�տp�
�D��<W��Au��f�Vt�_+�
��2n�����V����R��i��6\��H���,s����D#�e�d
~gxګ�Z�(�:��QG����(N�K1!���P��R���Ɓ�R8�6�	咩z�ϒD�������T�ˇ21it+N.�uW�+ޤR�o�V>O����L*�r5�p,�s�%H��	!�ۖ$�?Q�0y��O��PTTN`X�#��8�,��)&��9�`���W�FG�]�1��?xhL�(A���,p��������bK2��q�������d��T;��6"�#�A9��o���)�\��_�z�x#�;��Ѩ퐝rD�缗da�^�
G+&(M&ا����<�7$Fo���_��Z˜� ���>�:A�t#��Jd߅�e5,�b+��� ?/F!uw!�˙ӄV�Lz���9g%R7KJ��1w1`�ǲ-I���j�F�E۶-��-��F}���2'��\nC�\��t�Zm%�Y��n�u:��moc���(��'�q�M����5�%�#ǲe+[?TW]v�u�Bw^[�޳^��AB��\#?�Mm��^�zÕ��w�0/�-�P�A�k�UA .���+�=��=~���A�qW��r m�+L���7�=1*��)1W�y�Ùe�e��C*�-&�飿�R�vYρ���8�FO����:�txh���g۫F�����PI}1*�C~�1^����"���LyYp��Wo�Qs����
�_{|ɰ�|�T[+�&z_�6����c��X���{4���{�97�ee�{�*�N�l`���/d�f��yU��jj�&qc�}\�>�*��#]�z$$�o����� ��Qo�O���~�4�2gWV^�y
"m�~R��`�R� �y����uP�ܦ�3Bł�����u��/�n�u?^��6c�aM�l�R��;���5��nKb����p)lV��v,��\��'͏�R�{��D{���Z(��2|M��@P$���A-�kYN}��;�{�Ù����Z�l(��st ��%���3V�>l��H�ɒ�z�O���K&��x�t<�a`(|G���/��'��5y���5I�t�ܢ��8�m�b���_|Vi��r�Vk���k_��xp�X��0���%6��:l5i�YXM���U��~�SP�E9��QH`F2�s������.X�Q��ov-�.��1XEiL'1 �9)�!*����L��!�0O9�;��QЩ��b�g|�Ȕ�#
J;��uֻ���@'�\Ll���
�ȼ�5�惏�Y6��Oإo%s)԰ݟ-���Gyd,+o��'#�?H�r)����ĸ}���]�4,7U5��^E��8)u�˯�I@c������Z��ZX"���{�H���/u��G��ͦȘA��&U��� u͛�C�|�P�\*E���}�5uJ˸�Khۊ���n�n
�Zʠ�c�ئh��f�˯b��{�b�
��g�4:���m�S��^��DC����O_�8)I�є<��]^�{(9R�P$Kw��A&s	'�������}�8���Es���OD7?�cA�b<"n��R'8W ��T�ҵE����92&���"��莗:��?)Ue���U�'
��rTA����a�8q��K��T����K��}�$S����,z--c�Yc�P�������*���0���a���Z6��Z�A�@i�F\uZ�sR�XPmЩ�V]H����ٷ+u,߂#遽�����;`�K?x���V]�:~E���,�K�i?���<Uk!1�!��d���)�9&��J3;���ů���聑zˍaUl��I��	���ƺ��]U�c���5&��/`�Y�CZ<uH�eq@g�>���][�b�&�m�h;��b��\����/�%�r�=5d��7�h4�z�Uې�Va�Zd�AORw7��ǿ��$i�rZ��Vl @W����QZ�;y���g���̳]|P�mW:���-h
2pfx�	~{])!�Z���MSt2P�%�DA�hJ�Θ��Z'ۨu�����@~@�CxN�/����v�4�������@e��PޫM@�����#���d�����U��f�P̬��Co�	�7��Ӷ��;�9`����1���l*z����ŵ(���e�*U�W��^Ԇ'o��tV���a��C���+���jx���m4v��\@��?�����Fv���R�X�k� s���P��9*B��Ax���n)��W]D%�cT�/{�_
����L���8����#�рh�f�C;�V��ᒥP-v�~Ֆ�T�e����?/@��i̵����Bo����u��<��#N3�r���S��#��i�r.�����/���r��]n0g���XȪ�"���>���\�?���",��~����Ke{��_Vx�A�D1��($�Z�L�aQ7�Y��*�x{���*�ax!�b!Z�� �9G�dbl�c ���3D��#��SO���ݗ���,�(���7�|zE���.S<ˑ����~���V�|��c
.��*��_���!�ݞ�S��գ��2eë�'�K2�耷��[��ntE��=8�⮪�hO��a��g����+�2o=�G���/���X��'Q`�C<H!'�֒�S g�J�Q4Y�PΓ��K�IZbM����	#��X�e��|M�E=���Y�uJ�R��C{�/2�ph���`1�Ν�mzU���B����(��F���e!���i�5�~.5Tq�~��`�.��ȖzѤ��J9~���������BKШ?�i3~q��OU���d�)��,尌Cz���hOu���[G�&�-.)
�1� ~��C�p,ڏ�9����'	&�sh3�B�#(��+tTO~�d!���<��x��C6�I�'�Mńx�����;�|KtSf4s�#��H>K�{� ���w�扩�{����s�������n&�T��bF{=�n-�	m~(<	 V�����a�6��)���Sn�G����R=gĮS5����^'�0H)U����BB�,�o����7=S�\�}X�Vr���U
ډN)S������������pyD�l��փ��ɜ27�A�:���?:�LX��$ߌDw����5wd�f��p����$��}�U�Q��X2c$Z�����6��[���6����,�8��K ���K)D�º$�l�[F��soa[�w�`@_�Aަ����?U�A4��;�`����(��5wX���=TVx�#�B�2"�J{�zϜ?[�i�=�I`��l�*Q��8� ��������Qq��j����'Y@;jR���tv42�y،K�W^����j,p_�T��a�Cs��X�x��|�֩�6�O�!%�Ց�o�N܄�u'�`�1H������vS�֩bl��x�#ă�(A�U��*f�}y|&zՉj�@�fҠ�VW��PK�U{Mi�}}g��+0��R%I��$�L�6&@���B��+�RA-���]��.ηV$n4�Ux+#�G���4��		��s�~�T�Š�5s,��F6oP��aZ�����	����q��:{�\k��I��/ង�@3�����Z��B��㒜z5�� VR�)S�E��o*g�Ag��	~��~Ѽ��K�fG3U��,a4�*����s�6���p��EǸ��X�+�.l���_��ʁW��ie'��Іt2��ڕ���Mʏ>�%X�v�>t.y�q��]v��'B{�΃�!��1�>�]�N�R� �si�6����438ۮP��+���We�ח��=w8;&�� 7ddgh_:��������Vq-�vn�dB�w�8鴥KK��~�s����v�Dba�a_����#l�q;��`�>��*揖��؀����R3�cn-�X��lV4���0���D`��qX�??�$c�_>D��Sчxf� }�c�ԕ(���i���W�$�|�l"�
<�_�񼛍ҙ�����n�����K(�S���ŭ�#�\����h�W����� ��E�#��p1~v�J��|Ί��'�U�R�x�<eSKo޺�(�KK �J��� �<��B�Tm�[�]Ϡ�e*��?���>�a�������BKY�����K�X]��	5m^A=md|)�ߵV���1+䭵+���O�"�X��J�3�n>�c@���x|�����X;�*��&f��Jg�DJt+�<"7&: �=\��0b���G�!aC�^��Ҷ�Sx����Q�؃�4�}�m���ku�H���ۛVjEmm6�����rx舯a��� ��Ve1����`�_�,U��Uc�՝�dH���!!1gԦ�'C@�۔���z��o0�)GCg�9k�r
�������L`�T���&< ��.�Ia-�/:����Z���hT3�F
@춀;��sd�]���`��g��{�o��>�٨�E��s��ԑ}����Q�q	�����\�v����;�u$��G%�a��7�ȶ�6���U�ٷP����=�m�H��dƔ���Mn\���j':�K3��(��w(q_�X�h!S9x�bzr����{32M�ɲL�˗ں6|��a��/���%6R�\a�քsXUԯ��V�Q����$%|2�q��)�����eek�Qe��Ƶ�SL�w,Ũ�N��C8K���~!��&n�ig�_y��-c�j�(C�P����摌�k��,RфC~P"�危 �px�|B��7\���=�j6�h+��Ja�U�U&R�1�T���tў�*aQ�@�B߃�`��=(�L�o��)m�]J�O����G1N�lf�L�gdm��G'p�ԕy}�|#��^Dͮ�QQ҆�Ј����N��B]���3���&Q�l^-�¾
k@?�V�('�1&IC~����?�R����\+���ř�7(@ϭ&���X8M�ے7?^fL?)&8�9ޱ��MX I׵������ȕ�	���)\�I�.<��W�Ty��_Q��}
�'�=W���W |?�M�v`v���p�R_�<�B�9�\zj�̯����S1z���_�'�.(�3��my<��iε��I++اS�a\0ʭ3�诠�H�L�	S�*�/�j�"��Yt�@v�˨��MQ��4}�h�'$��*��������đ�Y!��ܜ�0��PK��d�^�-U�W�oV��η�����u�����h�k��$Ѹ_ݙ7�e��P��V#W�JBp�*i|I�9I�h���tҍ� ���隣���檜��^/k4e4����z�B���!2�2$�l��-���Uy��$�"�����:_�!M�#?�M���A*�%@F<���s0��ʪ�$immv�Ա��~bYM���4���E�(O<$��=U�-N�̝���`���8E����"�bܥM0�[����A�*`[�����D�Π��+g̃_~j����r��D�B	0�όE��p~L�¦�]l�d�;S�B]��c�A�]=��^�?e=��W�RdJU�����(2��R˚�}U�,�,�;�� ���9��-�F���D�a��!�$�kb]��:l�I�/����t�1��/�C��Т�kuO6�"Iu�O�1z��E�=B����}�ŀm�k1ňv�	Xʬ|i�)1�V#����W��tF<�%��>Y�?z��9����x����'���ݧ]�t��g9�8���9~��o�3~l�{:���LP4��C���}wMd���J���FQT��{n�c%�E)�=b���,TMx������%o�s�$�d�-�0V�y�аwb>��쏁��x� 8�T�R���a3��3���N��=�.�c��	�nB�+�w�؂�
�K�S�x��v�O��^�s9i�0D(ʍ�~t�Q�ˤ+��~Ucp�=��>�k�~!i����;ziqg��*k�e�k�zn���P|6[��D��*��-;VNN�M��(��#�A�Q�:O%���ΚG�AI�g�o�KG�9�,�	��v�8���� T�Zk�7+��W	�[����Y��y����NF6��8��'b�*G�6� R�e�I�	��_^�k�ED���x�b"Y����S�.�H8e���|찚M�AK<7����	2�~��*��;��uR��@;4�
�����_�����*8{����˟�LkY*��|��Ȃ���q�w$��>��j��%�����I��q���X�O�w�_F�܉6ˋ�fg���"�2�Q��[TN��U���Ү��=���y �6yx.�Ͱ1~��<�~Ohb6؆Fx�:� �Ԑ�h��[x�B�,ϱUF�{)�Y��ɏ�v>u�S*��)��C�Z�tF��t8�H���ȇ�S��Z���*�
���M���-2���������4p_��8�KGphBYa�N�B��t],PJH(Et�9���	-pek�ݺ�֪9�� ?�� �y��Opa��8�	޿z@z��0P�P��[�N��}�i��s�.���!�C��0�/4�{561(�y�;1pm�u�I�.ٻ�_ V���IA���کwT_@ 6$9��ٽE������a��qmU��HJj��pC;e���x�.ٺ����/�/k��R~!8յԫE��T�:/�"fv:�|e�� #�U�F|�;��~d
�r�bJ|�c�$�
`i��/v�l���ć~��I�c%�ʝ>v��VC.M8o��9��Uo��k�8m}�uʲ+ &U��)y�TA�R0x<A��7���s��a[�8w��?�#��ֵ~�����8P]�l�Tk�:��c���^{9窝:B�@;<��e��I��^�:�)��ǉ��T�!��s"�hnC9�`�lBO�
�F|�hZQ+8�qc+֧t!Q��Ir9��S���(��ywXjŎ$e�wP�zp��~��([��\*�t�u���+�SD���Y�ߣ{�n����ٕ�`A�q����	\�em�$�<�ۇJ��p5ِ�4*g��
��ҾA����y86ՠ���V<v�6��n=��g����S+P�a�\?'m�ࡠ�����dȹh����}ܱB����bA��W4ZU���"�6vb�eUf�sv��%�g�"zJœ�n�����I�-#\΋hm6-VB;�91���ֆ�	�::�y6j-�c��Z��^������HK���/0�����G(��V�g=R��LO�[ ��G��]�'b�#�y�L�/��ZY4-p�Q��d,[��dtǋ�`Pߴ"�f
`��J��\�&hW�ݮx&�$���$���m��̄����h����[��/�75�!����F��31We?�=�e
D�g^�mm�̫V�d��'�/����Y��L�|T>���i�'H�z�n�NO�%�sI��A���g�G�y,)��n�(ʶ4�0?� ����vLl�=��*�/�.�d�����]�8�D�vh�
Q$}�ʦ�>e�����@��y_d�f��?2*_q����⒟)[����p�A�,�I�LW��:W�ю��+�ĺ�9�7C+�w��7^�:z��.G���
/�K����3ݝ"��<D8Z�c�@��w>�L{������|��P���RX����Ĥ!����H2qBcM惣��88�����j��
���Ԝi�,�sVZ��M�Y�@l��W$�N�6�>��z�Gia�Z���-̳��9/CJ��+	������~�;�����s_[H�i�ƴ_dk�SL4��_�al�ISY����uj4m�]��H��=�̢(j`%-JJ�����M%L\���W�P�Oߍҹ�6�K��k�_5Ud�J�)#M�I�FFH��a�c ��T-��	��|�A,m�ϼ6{����:MGNg�e6 �
(����h�����\��ݠ6"���ۤ�rl�P�����,Su��#��ͨ Ů�6�~�HO�֫��ܧ���X��)"w[=+�͕C�^��i�)kDހ�\ɒ))6M��禇�>~B�7+��^���z����f���	�0�sb�M�&���1�[�w9�T¢Ȓa�@��an��Q�&���]�Ӭi��M���`r��Ω�O>d"YW3٧8�"�1�n�� ��S�Z|,M,���y���8���(R�2]R8"j�Y��%�P���֧2F�s�NE��fK�������J��1�Ri����i���Xt%�h�$�f�hae�j��M���R^�.3�#F(>u-J)��{6�a��\Νm`��o�}+5�I4K%q�4�p��:;>�K�䫈Z5�{H��M1��K�s-T�'P�Zf(����%�1�47�5^}p˅j��(�B����Vxv���~+���\C��!k2�g;ܪ6��C.��V]6�!�*�1�iG2K���,p-��S,�t�,�X���2��íW:P������5ĺ�=�V�.��U���l��H0���V�����Yw����ey��<��>��-�HC�l��|'����ۜʱyz"Ytӏsc�v�8*�1�G��� �,�D8�9���N��ҩEA��1IG�����N'��Y'Y�ֿ`�7�����p��%��Ϲ��ɋD����n9Ԁ���=���4�m�.}����M���熐�B��6�L�T[�T�Bs8Y������i�J@.��K<��3�W�>�G�-��ߏa4/�'1�ͩF|�Фk֌�W�*h)��4�`
���C"�I�BC0d�3y�M<���tv�n��>�w�Ū�R�_�q��c�0vE����ӫ����
�S�]%*�WA#(Y��.�~�v�Nb=�G��p�̉���n�d'�N��(##���O�u�(7��ֶ���[�W-�BΪ����Ee8)O�>�wW�U(0B3����J��>_�Ꜥ�sނ4��߉G-�����5�p�'�8k���Fl>6m�iRCi��l8 �'3*�>�Ce(N3��^fq�HE���Z�mu��e�
���ţ�PSD�e7��Q8���_'�MI��F��Q,�}�J�����Y6���7�:(C�Ĥ�E��3�����'=�ʨ['0��4M(!��y$iqPdTY�����Pd�M�̹�=�}n�|˃(]-EI32��9&_Wy;�����gt���뇎����=���b��-��n�����S=�&�"��1/��ﮭ<b�z�FeW���(o��_�)2�h��5g��ä� �-7��f@��!��!x�;ݞ�+�G"���F�wG��h���X��LCG!Q��57U-��]���e�8WA�4BC�����h��&�Mٓ�������yRVS��w}����a��Z*�j�vuHj,��ɍ'��f�yV�V�W���j�<X:#�db�j��i���7�~�"�KM9(.����'��ZA/.]��}>�}�*����L�!�O@ �:�H����c�i��v#� �����}`c$��TK��#k�A���hrG���0J�Z�%y��)ck���	���/�D潸���k�05M�����(ӻ�H�]$0T�����<B��@��ݯ{�l�WǨ]��W�?��-����NEUFPt7�jeb���|��0�pb܁N\V�"�)��>M鲘��am��_c,$L�H�=��3F�Q�#�S�Mtz�	�D�F�1�_i��ee��(Fw2+@����	Q���l�!�YG��$ ��FQ!8Dȯ��T��4��G�����>*IﾭDP���G�L���ؤ�����A���P������ÌkI��i61T��ڏ��\9yԥj.�Y`�I(a �X�l��_g��؀�-VA��i���
�*A�{>�B�*�&����<�@9��\�⁶g�����U|E�^��2�xd�|����4�<H9�]˵i�W�>L���v�9h`7$�W����m�����o�����+lx\�8���U0���|Yc���߳�'L7Es���?:BD_�r|5+�P��k�ȭ�	8#��.q� ��=�V�-�Pa������J]��[�FEB�\?Y�0�.��K�S,�Y�W@��m�L2�"�D{x�5͝���>ԟf^!q�)X��0�斂k5��w\y��7|������X���Ě�O7Y�M领Z�]Zg����s��(y��խx�zb:\[�Z���K9	�;0��;�q.���t��pO����y"���JiOؗ:W��0)"��ӵȦ�E��Vtځ��)bz�/�����ۦ�yů�l��J�����~�"�X����؆H�턴����Mc��3s9���6�/��f$�����pR�������Xx��I����
��12�w6VQ��;?���܌���KR����M��,�/Ր��)�C������\��U�q�Eks�46�7UL���$Q�?�:�_W�]�+�h��רA�t�to$��@z�4^���}S�:4cd.v /w�֯���J���.L?�Tnߔ ��J�`RV4�3#|�.U����Z���3���Ȉ���S;��C� ֏2�"��+��5'�3)ǉ�ԍJ�1���>���P�,?6�7�5ʨG�?,� @����*��k:zL�-�g��D#���Cl�l*c�q�E8[f�(E�'*N�^G�a�o��Y�:T^?&�cY�/������٧��Q �o\W�O������@�c�K]0��b㈥����M�R�i��L�=�ӠyK�j��XN6F�S���H8\�����9�į,ho���k�|�Vo�a܁�T���L��r����@����x9.p�N���GiR���:+����=�i;�u���
7z�/���D:�k��6�SxT����ͻuT���?� N� ��סrU�=U��ԏEګ7&Qu@f�H<�Y;��b�ߡk	�D���7H{����'4)S�F(h�6����oK܉�f(�M��\�oR3���W�%�f&_���Ψj;Ҏ�N�V絝�=r�6XI�Z�����o�~�e���E]�n�WXOඨ�ٕ{�����aڴ�,'�n�!x{��D�P��M��mc�Z�#	AY|Gd�A���/�0DV[�<�-2��<d`^T0�����M�w���ٹ�Ύ\���o��&d�\���:�Ʈ-�ym�'�N�SP��Z����������(=���»Om�ј����4���"���D�	W������m��KЋ��f�E��~Ɯ�Y�����?�թ��W�`���DW,1�̶���䊋0n�zv�w4Gͯ��'�����q#����G�c>�)6^sL$q�AU��lѢ(��2��>RL�nx���ɘ�8S�'�Yeͼ|JM9�� ���J�4�un���������=򫫆��X��t��4}w�{ѥv�^?��(I����.jx�ʌ���*�����rX��+d�㔽���t�:�цĭL2\މ��Cv���p��s�!K��R�C8�zgF$
�Gcﺫ�fٜV��TR;m�U(�|����Z�n�ޡ����b���;���jy̾���HW7�n��y�
�����)m�B��ۗ��g0x<k<����!�����Qɬ �ˬ�A�!�޵���A :'�������Y"c�ZOP�&5r��b����2��r7(�	�`�i]��Ӝ
�i�NsZDO�X�1Wsw�ݰ�m�����Q��	���E4������ap!)���^_��
k�w��u{z�����4�/3�(�9Y�q��_�U$ol���6tU�2���d������/��?ԋ�f�<�v�t�g�ʔ⣜Er����!�b0?��A�m���4��.�h(��̦@��۞������F�J��͚��W����a. �i�������Qۣ���3����'A�|\(^2٫(fm�ͮ~�������e�hf�+'J��vEs� L� �%p�o~���>)Y4��v���Tϴ-�]FrK�w!CI<j��Аy�G/?�o�R=1#T���!�c:�"�3���f��<1�y�3a���R��ظ�ނ����ɢ�l�X�������ȗ�8F�Y�
�1�4�:�e��ƈP�>Y�Յ9����)���	�;���ҭA��;��g���-��+=�j89�)�^���eT3�:l2*�_e�R�gq���M��P܊YF�u%4��.ޗ�~�c��	Z?4õ��n=�8���hAȠ��àD�qV��,���H03�ycnQ�XOd
��qg_��(Z�� h�҃d+=�lN΢L�H���.��ߘW�[`�42&`̒��D�����	�MW�]��}��O����#��u��#cc�KUv�wM,F�,9��N��!�&�3^v���yBߦh8�N!S�����1 }Ş
��F�!N�3'�D�%%1r�I�kT�%�C�X����Q��o;�ߧ̤(�Csh�d�=�߭���%�A�锃�M���Ε$��<�{�K���R\N�]��ށA���U�6	NÅ5Y~{ ���Z��(��K��;Ӑgf�CΉ��4� �>2O�M�{?����ȭ���iS�4"w���D��_�3=�V��:>�7Vs	�/��+yu0�ل<�ӟ��|�+M��[�?cZAH���Vo.b�`e��˛U�"ճ���\TG[��MRA���8��WQf�V11{C+��z|�2܋J.�@��I�s�T��}ͯ1�����}���L"v9:S��
��[�a�(��k��)�ǔԼ(��mmF,
����">�#-(����qFK�Ln���@�����H�L�0&�U�6�A�g�ܪB*�����s�D�kR\�u�y�c/agJ;�^@'n�2k�S�Q'}�B�:�\:��44��T��������:O����PfI}��Ru�n)�9���t�ӵ��(zP�W
�$a`�υ��*���(�/҅�yv~RAoqm�A�L�Ж1�?����We3�,�tz�l;0����Ns���ix��ҍ/�MJ�J ��$(��r�&�Ӛ4�?��fm�EPk ��'�ȕ��BL� m��/���
j���c2������,��m^��q�r�o��!��)�h��A���\oL��w��r�����*��`�-�qnbB�{�-C'T�(�&r���q�/�d©��B��_>�}�˟�}�p-���-#XO6�J���V��ɬY�V���"�=��,���#�+n���F
��^��^xE฾��EC��Ĥ��i�:�XCrҌ�xmW��Tt	�T����o6����9�콅k~��e/#˥��wX�
�@'�[��飩���9:�	����������a�t,�2|����q�9M�[~>-YSM���}��fՇ�)�F�_�u.K��l/��W͹�S_H*|�y�����mb:�<���yI������?wdu�#[���xy1'n�D�	0�p���I~�%��i���Eg�������ԅzq���u���A=����+!��i&/���U2'c"�:jGvr;��e�Q�|G���4��FR���X��8+�;��Ŗ����l�w�p;U���/§���N��r+�дa J���I�@�O4~�cKK��GѺ��	��_J3�W��svZ{�O˿?Y Y4o�;�Y�f8�������h�Q����F��C�����J]+�A!�>.88��@c�-k����Ui�U�0I��'����9)��ށ6z�h���K��.!
�D�9��x"DH=���zh�>q�+��J)�tp�{��Y�\�z���"�}�k��A*��F}��K)�뾏ߙ�i*��(R���z��Z˧p���f��C��Z/P��x<8� 
�����/�躒@�o��N���)���)�Y�Yز�+I��������<H@��<q9����q翐��(v��,
Va�̷�%.��M������ N;}��3^�4��������s��F����9���sI0��vQ�9Sl9Y��2-hb?IwD�2�J�3Zv\т�۠�wV�5��j�C¾�&rSyM��Γ_C8Ya��t��)i��^�Oq�#n�v�o��5#�r�=
���z�G��MD��~��`L�)EgfU���&<��;�F]�s	�V�p�TAH�o<$!e���_�i����q�(9�r����dhE�T�l��	4{�8K=%�����E絹�.�0��f�����6C���fe��5z�����cX�FE]�\A�>�~���ȒlՍߗg�.:���.�����7��mg�=t��^v���������7�=F�/+��2=M1;�Ǧ���A��O��Y,��o&H�V�:��]�;��N]�SVW��%�V)�  ڝ)<`��Ա&��Y��M�ݲK�|$@��^��)�`��ڈ!Z�a1�TCf���V������[�Y��7r������#���,  F��GG�'�-q��P�m�ܟp���	Im��d������]u����!B'7֠�?\�a���ա��k~\~D���\���ُ;u������s�+��_�ɭe32�B�<t��#���b��EcS����o�R���,����%�����Wz(%�0����6q{^�v��샸;�-j�p�Kh\�խ,�`/��qԢ5��%�ɽ��=br��a�c�s�ZX8},U�L1��Ļ�-nj{��hFC�x��B7v~�L�0)mmz2��r������	_'L��ߩW�9^ՃP����� �+�Q��0[E��%Om8�!ޜZJe�uwr�zH�`"P�{����|s5+��,���Rqa	�뙙�� \J�/��.P��я�#�^�� ש�SZ�S�q�h�� [
,d�v�u0{�1�n�и����͛��[�~�g�DhZ�AGD؛���UF���;�p=>X��Q+Ɉ�R�����b	�X�z��!��C�ڂ��ӸE�+�)f�*�kQh�QX���A��.�w���Ɂ��=X�:w��n�:�8X����H�uǵ��w�s,(����Bk��5k#_R�;kC�/��Y ���c�P�[r$!�4Iң����o��L�������p�[NPuE��C���ؚ��24Uj�	9DP�CbK{A�=�?=�f~����D"��C+J* S��_���A\�j���x?�9_��ai�2qO|���̰Fv�����=6ᆊ����\��}�H�9������_)�,	x�e��a��B���;6吓��]�����Pb����R�����0S�=]8�TN_}pj�cA�ΑJ\߉�_�W[��>ˆ_�$
����P�-|T�*��"?~_)VH���n��?��D���sX����U|P�ǂEɭ�l���6ܵ�z'��$�3s��w�IV砟Z�Kk��`_�������Ì�p��8W�#�3��W�	�/�Էp��Eu�{�ͧ~s��p�=Ȉ暵�:�t�5(�	�Q����p��e�|]���I�e�er�4�>�+$�Kb|��~k����J�� �M,��hx3b����:En_�hy�ԋ>����bQC�!�.�n�m����9:wD�'�L�T�0��^`�x�]�E��e�R(��;�A�Q��������HѺI�T�f�]Ɉ8�7<㜑	�A���Ҏ�\;ڡs�/H[��tH�t�c4x	"#?�ۮ"���L�^�� �`c�-H�����4:ϰn��^��y,�x���P��Mi҇ ��v_���28�X�k�f�n��0�*����MVQ�3�%�qB�EFPP�"]�a�x��ٱ���w=Q6�����{��-��7��D�C�\�~����K`v�nW<�Kc/z�\�}��5�c$6L�;1�d��@I�����;�\x("��s����?���ٴ�P��9���aQRL^*�ڜ�ur��t	���	%�>)P$yb�>��x\��|,ѝj��V��N�^C�T�p�v�(_�}"�ӤU��ח���{��s��}&~G<|c�\Zjob����v@�k�J��
 �/�;�c��WN�W���'+EH�hk�����4�0�����wQ�A�K�Ԡ6�s�5=M�8��ڱfS��x�ɻ�yHd� R�߬`��R��"�~Yڐ�/,�)֔�.��D�ĳ�jr/�V(�%o�"�9M�T�_S!���}���UiL3�db��'���AB���\̘5rHf���l_0��e�߰�z���e�|�r7�~)m�[��*�*�`r	1(�cŖ�ʂ��x<͊z�u9�H|����fEc����b��&CC���φ�tQR��i9�`Ch�����곬3���w5C���س�!t�;)�ry�)����1�eP8��=�/K��$�h��LM�̊��ey[��Ķ�{��{�f��%�Y���Vg���9^����ih�)�q�`^� ���14�Yk�
؛Nŷ��"����(׶m͏������}`�0�nXk����\�����MV^Z�z1��{�	:BF� q�Q�ьT���Z�a�5�˄�$
�J� -��'i����5��Y����0/��wRg����ؾ�hj�C��h��1o�u�ܲA-+\<-^�ӊ�ߔR��C������#�P>yyx!K���"`�Lr�-F?�O*s)��V�Gٯ&��!j7�e�a޸b��(@��� q�`>�D�ȅ���mba}��B�MK#Ԗ��e�fbB����,&X��Q��UJ��2��"k�\H�,c�(5s`�P�/&��e�ᤰ�.U����ʼ��`�D#�N�P�Tu�[��ߚ�0�P�fL��b=U��^��]5F?y����<�Qim˪�4x���ɠ)v=�,T@6���wMoW;T�` v)�(�Ϥ�d�(�23���`�r`�H����Տ@_ֿDi���"2��0þr����9�' l���Fc��Q<�<}O���^9	ɟ�qi��h�-�GևF���������%*3�c�.�)�8�n�9[e9�i�:�o��ya��4�W>�(~W����BT![���J}r)���PfS����VP�g:�mfMy�Ѥ�LK��C�jH�&l�?��*�V ���ȁ���c,�te�[�x�����5| �p���د�` hE���c@��x��dx��6��}��c`�_Y^i(E)��rt���ֈ�7�@��^� #\�U6t�1k�[\�KLi/�ś�pː���.=��s�HM��I�t]U��q�3�z����$�8�XT`菉��D�9O���SY���D�H�:;�K��Ѧ����q���l���щ7��hd�}�TP)���,c��u�,���)��U���Z�W��p�·��w�a�[ �ǎl�(��k�GRT�.iFR��1����:�Q��Ira(5	f�R��e�pE5,X��7��y��(��0Op dyjR�fF�_	w2��si�F6���@vX����q����?�2N���#/�lL/пQ���-@��f�~��x��5cd0�QE�A&D[oj�"��QB`U������e��xW&��)���n^T�Y��l���6�R�q��^I��`�p�K��	D��'���qNs Էu����U'5���yƳT�ǵ�����G�r�|3`��dR0��z�d	�R�I�+9N�Jqx+�G�q�T�V�UIƫj��B\0#��FU^���Y��D�P�ND��'�"h�?�R��V69����@F"��>�.�ɣ4���%j�JRW'x�0
U�V�M�WaW+)q�L�j�m�:��
�),]^6���2�W�j�F�!�g��bGڅ֍Z��՛Ѿ�L�zm�R�;�[�LB@�orkz&�؄�4���}l����0޾pp�3��~b�t�&�5�y̗`��%�(��mWv{�#X�u�Ϭ��fj�<p�,rc�76�4��zxMR��@S3���K�(��t������Gz��Jq������7q\����H�s�@��9��Ŏ��a@����t �C]?��SK�?�# }�}��EVU�����"�s���˴s�F���RIq�-#$l	^�ʏL�95L:W��|��C�X��u:�
��רb����6��e��g��s4ǧ����m��a62j�Öz��
�s��'�2�O�R��ݪv:��jT�zp<�d#pClI[u�ʌY����fA:JHk������E���5S��A�j4���}E���p��k�
z��Z��~���������i�i�Y�:�߂�\�Jr��j�^�s�sd�I.C��3I��Dtac!L�������E�Qy��w2���*o�L�;#7���D�r2�X���={���kV'�����&H��D�i�c��[ܼ��+D+� ��e���i�е	g@aA\������.�����*>�@B�G�D�f	&3Z�#9����S�����h�#Ǘݗ$�qA�E���ܜ����1�f�J:3~�eD�#�D��M�Szg�3Y�	��6��|kk+��r���,�>D�YoW$]Q�vr�S��9]CÉQi�S��@[�+��)g�#�<�IL�p� �N_>/(��u��z�9WE�X��'cx9Ǘ�qߑ���1?)_<�@y��JB�_z(w�؈��@[1S��8�Z����z�R���*9����?s7�5L���\�{�2L�*1��=������<Ie�}ʝ��g��b\�R�&A1t�����]��&8@},�|�U9��= �����­����q�r��$b�$��<����R�-3wP�\$W2�[b�~���9����^��Q��2 ��B�����e��%}v��	n�-!=@v��
6��]@�^ �@��<\�3ً�׸!J��}���;��s�2�����4#<��4���[������)��1�
d���*|�C���7��-ލ�N����j�ǚzx�F����=b�کĚ�(n���FJ4y����Za�����#w��t������K�m�����M9��-!�Z6�!�+�XMs��bM�<�`���a�J캁����k~��oj*��"b�@�.E�@���+��J#�n!U�9g;�n��V��+��yio���-�|��KUD1'4�>_8/��$�4���)~?.�Վ�u��4�=Fpq��9 �}>�/R �h�q�ӟ��񭧿S�����W�Τ?578�r�Ù�<��NT?ߔ?.��Umfv	�Fj�rN�J�Rl�4��	��VDf��Ub�Ӧ���wV0��#�bQ8\n�%��-����\b��!��i���C}����x��'�H�F�0��ư7�5BY�~O����o�]A�������vz�/Ĉ���'�6�u�������z����feر��<%"���,�NZ%@)���}��gs��Eq��{��ٺ~��cE�`�a��]��&LSV6v���9�և��+�ͽ��{�օ1j���c	4&���4�<A��N3c�&ۂA%1H���K	U9���x��*�Aٷ&��?��`��S�¼*��@��R ��|���ˮlҵ����d���� ��L�RA��<�f[�Bv���a������TOr���!~X���2��K������=��[T��6h�@�5ތ!Z��Xo�T۩�	A7�W�p�n���ِ?�����5��6�*-���J�m(M̎���.�[��JJlRq#�6˳Bz�N)��D�!����|�w,�A��� �6��2NL��]yY=���{w$u��u�eC��<3U��ZM?�ƵY%ߗ�G<J��S}��{�R`�d�6�[�e��� ñk�H��U}�;���]���0,�����ӡ<�b��tӠ�à���W1g�� X��T��uvT&�_h��?�R<��m�R���"@Nu�D�{�8��������.�C�`a3E�oJvC������(]���x��)�"sȾRwQ��m9L�k ���+����یO`��{��Bfó�Ņ�(�<���k���>(�^��u1�W>J�A����L�M�u�GT�M�m�0�^U91T�Q>���L���~	J��� ����E��|Hx1����Y�Z�m7i��]���Gz\�o�=�����W�����$���8�;u�3�%�Z5�V1E���Bg�e��Gw+�7[��eF�T��!Ȓ�Gzxi�Խ[�����l�G��=]�w3�k�~92��>�WΥ
�v�O28߅s������ {y1�1Õ���.�N�	�"5ޚ^J��{9�c�򭤠 ��&�~#^M��%s#��bT#'���>���qM�zGL�}$�g���@�.�E�5|k�6K�kl:����'v�r-"	�I`5î��(_�������}���]��{�;Q6�R���5�|���fs�lwK��	�K�D�L�D<�p�VmS�Xa�a���$0@����\�7�6G�h�
R�SUO#}�NK�[eLÿD� �^ߠ�Z���� �W�J�F�9��h~L��Y;WK�{�U8 o�d�5Q�q.�,B��mo�/�ԽI	��pǮ,j�:!��]<1[mo{T�c������ғ���"S�Bݭܭ�Qnh
ER��^�/	�ʾ�;�RT���d��O���G�[�gY�ֹp�Π�@��bh�Bn��b�����l\�e�JEZ6-� 9�K��.^'�R��A��͡�:�U#P��J�R��54^`�L��#��#^sx�Y
�qU�#�̺*��=2�NI1���S�%�PR�ڎޑ��U����7��E�����$�_}.��)5�����\��ܩ���9Q�-]��-��E�����ڎS6urŎ�a6k�; �+�����Fݎ¬�S���z"H�C����VxS5����mJ�����L��̤ޔ�U�+���������k�I�G�,@I�ҝ˕�!)!a�夗�W����>$0�g|�r��3 �%��]��Pk��mڴNs/;�����s{��$�2Z��dI��HAVs�>k�b��p<<v�-�ĉ�Jv��"�f�&d3�]!��ed��C�B2����jȟ=�I�t&p��+��g�fU4��!O��^��Pls��G /R��p��^��8�?�۪Q��-`j'��G��އu�
�+Jh���E���t����|�!��\%���쥧�Bu=&^�RJA+3K_��|V0��f�Gb�|������zO������T;g+�Gg;����Ԏel��^ەS!,����,�f�	��#�ܙ�m٦XE�f�_�P,�i���v�R�M r8n� �ko^�B�V�<�d"�K��5*c3��ás8�Cf���]�u���}P���J���~*|Eo[[�=�[�I��uhҌ?lst����B^z�_���Q���2d-��u��"�x�h�<1��E�e�D��r��q�("�+�X��5��jY��@T)�͘W�1��"@��ѻ��#�y$8˖�ؠ����|�h���'|��<� g�q��`r���Hk�`� ߴ�'Ŗ���5��0E�6mA.�̴6ۉ�KlXY�zƆ���b,W�Xއ�<!��M>�i��N
�����Y�`������ @l�<$����"�i�{*�����J�(&�z��5 ��Y��b���8��BŲ���@?8e�F�f;`�����$lĚ62|d�����&7�Y����4@��,^Ţ�(�$��C�A�0��I�Ŝ�B�E_b�0��[l�.>�"�B�SԴ zN�7�ֺ@l�΅1���Q.,�%��d����Mx��N��Xr��ȴ��I��a~��&���w�h���Y}a�?��D8�����`Y�W|n�RFr�MU��	�~��)��r����+��}if�<��"�{ܥ����b��J�q?���G-%��E (��.%�%+� a���T=X�Н�^�xvoR���&���U�_���V1���w]�C3Z@�퀳����?�d#��)CMb�8�:H��:�NF���/\A����瑚j-�a�����&���-������s����_�DۉL0�p:2�dm��bL&�%	9�ƪ�+�2.0�O9��y�x���$�B�1cZ1hP?m������V4"1L�<��qn'e���{|.�WQ>���ĺ;��d��h������������!��QuT	2�.�O��x�]�9uq���}�p�Кun]��))R�Kf,շ�����&�5����Q��v�@�,����h`�F�7m�����;G�v����@�_o}�� �����m!�?lM>2d7�-2"���=�]�ԍ���M��E�x�dt(��-Q��*ԓ?!�?��C��[f�\v$�{ȵ���}�z>)�v�RWqm��i�>�cV�ͻ������JޝS��N6��H&�9T�:[�`�G��������;��g \��R4��%�{���NM���u����8S�v3�X=����h㑜;X�I��G�Ngw�����|A $�T��Y"�_9T.}A%'D�Tn,��@�j��:��\Q�ķ���a�W(��W���$O@K<8�C9.����g��j	�r)u�9�3�}��sR��y�� /�#�ޥ����n�m_��ͯ0�s��V�������W2v��Ä�B�Ց�t7+S���^�kU��Em��s��9�S���,��j�Qo��6Q'v����D���{^ͬ��+P}}L%ET�τ�s�STn������1��9���l�8#Ķa�#S�p١�P_~@�D�)� qL�:y�=|%����.{�:J�_�X8!����NEX� Kֻ0E@���{�[.�$�p n��Kٌh���0)�"�m:Q���eɑ rd�(c�S���.�Ӗ����^��;K�$��޳��FMʏ��k��[SYp�C)G��+����\�zz���z�Ls֤��mru�t$�>��Un{��f�Q� ����t���R�z���%;ȇ��:6}|���aJ�M�,���1��#�{�6 ��}��[~�$ga''h�a�R�����BB9 ��M�|�,I� �о�يH4��g�u�W���s)���"C�ڨK��e�0Vv+S�-P(x0�F�1ə��䤎J�L-�����cY�/���Lɘ���X�m���P�1���kF���"�O{���E���=�k�X�'�.s�8ae� ���%;�bکR��I������p��A��V�=�D�\�?J�l�0׽A�Ε��24��2����iG	n��~d㱩��kU�KϦ�1oX��z^�����#-��^�V�{y�~_���I��H���2^\�s�sk��t �kQ��P��*��ȋ�Z/�A�	� \������z<i� !:��=,)RA���$��#h�� ���C��dI|e�=��Lr6ѹŬ� ��{�\5V%+8�O�*{�G��|��Z*��Q�4��n�7)����'�U��N��uss�~蜣L��5��v�y�f&o0���0��"��0��q��5.����c	u�$�{��މJ;���9�E\�D�aƊ�r�l@29�*�<� ��oa��f�=n�
��:Ĥ�/�/�@Ӄ�|-"�<r���D�Y=��2�JGi�&�Ŧ��]�͐K��u�F�\�}�O��ڦ7Z=^�������A���Ҵi<�?F�?�	�<iV:IZ��F*��Q�|o<�_� �~y�2��1j{|J�!���{N%�Yn�M���X�6��6W.�e�DWD�s���/�0�=c���l�98&)��Α^�-`��CK�0���ZkX�"�#���&<9rs����ݒ1�郡5�Z�E/(&^\���ͳ�	�x��T��hD��:�'%��:�k "�y��}P�t�Ee]<d �;�M m�d�����O��Q;n9 j�2��r�2�̼=���O��l	Z1E�� �;���r����  ��-6L1����/Z��ŨRZ!���X���8��!'7�%I���~<۪�o��"��%g�¤=�%F�CmA$d����s�W����׍'R�ܾ<<���[��,w�(��"�����ڒ���a�S(�;2	s�P�'xSȥo����*����BR*��t�:��x�1	��Z�vfG��^ �3��� �U'h?�m�.<�ǉ�	��̮�d ���n}!���ws+�*8}|���%e5��T�����t$�='�yz�7�1��u�e��-�����~ᶶT���噟�C����������h�3v����vD|�ۢͪ5YYC!��p�!#��;� �ārsg������*�e�dov�7�]���6�6)-��A_13���#�x!��s���J�j���]6|���5����@I���m�i[��-��<��-{-5�X~��Iq�ί��ֺ�_F>e�
;< i�
��ֹ$Hj�ױ���"���Aǲ�C���C�َ��EX��6q���1T�����GY*BVX�
0,���ԢY�2Y�K�uq���ڕb�>Wid���Ӝo%��+���n���3a:�vc�xs�Y�m�:~���z��%�r�*����֒������3�8f�©w�onh���=���h�TY^��S�)sȖ�����aefs�F�>����uk�c#n��kU;y-�d��f�X��7���A�Wz��֗�ŬjO�`f�\,���r✸� �N�=�hB�޺�NH�N��)���eƖ�o��gdfq,rI��r�{V�#7��G�'�M~�uz�uI�I��<�f��k���c�4;����%N,�C�;�O�D�[1�4m���SШT���g�A�Ɖ4��]+Q�=,|&b�:d�.S����V�!�o��m[@�YH�d͂B��U�Iُ-����W	"ّK���@�*R� ��j����l}>J\�ng��Get�ϵ >މA�HM	�0���Z�MbPfiC^��?��o^�̋xp8�����X:5cQ�nް��+��6q��gm����� �*��JX����|}�C�A� 66�DN�?���k�o����'���,�:�2��MUN����5���j�1+J�@6�	U�t��	�z:6�O�%J���R�V#e����G��䚾��1�5z͒A3��"6�jG�/�T}4[˪nm�d@��O����Q/��5/�CtI�����V,׀0g��Gc�ȗ$�:;c�a��e�_CJ<�<W.ݢ"��v،o�ˎDjT�X8�ʳ���mZ�����a:P�+�@�f��a�qI��S*�~�s[HS%Y%�#}�N��3�n�����iz������x�U6u9���)��W��<�w�_<��&������
"��+C�~~�,���3v�!L< ���;E��]����눹Ƀ<��D�Q����)U��U�"�����1��4�+>�pS�e $O��aKR�𴈄9�ļ��e�$)�k�<C����D�˸
d��u?�O�g�_��(R����؍QNa�#Eo��bAkJ��wZ��NY�3�h4�/�_$c1���r�a���e� � A�C�`�E��wb�J�eh�i�,��]Q�kk����T�'J_c5����͹jx+��`�]��Ü��m{
�VV�/�5���A��Qˢ
n���i9w�&��ef��d��%�]�2�D�,��y��������(��3H��%(֢ 9:|��#bY�X����2����n6s��'ݝ[�)�2){Yj��=���&����*J��X&o8�ߠ�y\ w*)�v�~Sb T��O��|1���[��}N�a�qP��*yC��I����ͯNo� ew[/�7=�z��!�[��9ɠP&�)��6����oA�q��i�xB'{��l���,>��}�P���뻿a̵1!�lSK-5&NHD�+�Z�z���v��;��&�<c�M�C���	PaqMuԌk�t�Y���������&!����+��c��em4o�hmh�XӞ����]��U�L���s�:�=cX?2��V����ZtE����@�~�w���
��_�xj U��'ͧ&�� 0����lv8z�<r�s���`��F�N��;��uC�X�:9��	��A��I�YI������'��2���%�F՘;��́k��>"@64�Ə�Ȣ)f���_
�zݏ&��9�=��O�F,�=����@�ƶ��!�g|Z�����Vi�y{��$H�π����x��M�(�ͮ�l�H�+���_$$�Ϊ�����bѺ�'��y�\�������7����p�����U�ːh�Uoe��Z��0�מ�+���m���iY�"QV|�c�~�.8�P�NHPVJ{����p�b([��=9nU|79��D�a�v���?�*�M񲶟���5�}]( q�K~u����$4�a���7�[X7�g�an��m�����L�~{�!p�'�&qto��<J.b�'���@S����3]��/ð��SE/�=�TtO����	�k��	�oA����,���I�'-�S�P���U�2�0�q�f4]N֗P��w{z�T���d$������+��i�M���[�����t������(�u�~$BM�w��BO�"������,����b�W�5l�_�b�5�m��6i�-�C=;rj� ׺(�Y�B�I@E�o��$��X�C?h��.�>���ʖ���������pn((9Wk$�{l=oi"������#�Y��7���i~c-I&\�,hD������=��T�'�K���3��ɷ���@�9���~J,��B��~�w�Ԅ�#�m��_�����.��@8��@)�\����H��������0��x�u<}���Kj� �Wd1vW�12J�TK��:(ؓ�m_�I�����*��(�0��#q�o,9^�\@Hϱ�o�K��~�ͼp��,�F��K��]DU��mly�Fv����<�e�,:�ꡠG���t��6Ҥ��lW���ΖtPvI��*;�,m:�]ދE��>cո�DMdv�e�e� _=����H���b���9�5!�ƌ���Ao8��!7 ��x5.�r�����TBo��'X��K$�ݷ�M���	/�$����W�3����e�Z�8v�M���F�c����:���(��`�ݓ7V��}��'�qʝ(ؔ�y]�M�ރ%����0���ܮ������p��؇���]�Ь;E���H��s�A-��g�����m�Ec�M�ׂq'4�Q៘����&v��u��"Bp0�Y�y���"���;��ӓ�uTD�o��3#����(��L ��Ɵc( L�v�tK��g�[_�[�>�A�o��o��ȯYI��@u��]�TH$$�s�� �[�+U�lTcz��6s2H�u�^�n��if3��a����Ǆ7�FX�f��^�����{���~Z�ƻ�xzϝF��m�'�y4�w��V�<�h�<$�([}J�f+'4$$4�A{��'�p٭�?����:W#??0m]�V�xz�᯸'yO-y�h�HX���rb^RhZ[���	83#=�m���z�o+��:֓��:_���5��d��GO�c7ǚh|���ТB���-Q)~\Լ�y᱁s��Y2���	+#��OQ	;}Kt�EO��e㻜���snݹס����I|�ڣ�a=S�wz�-��G��M ���ZbLf���E��FMm����b�zm��yE�u��׹>["�s��j�yE�,p��ѿ�>4��x��DN�a,�M�pׄ(�B����q�^(�e�S7���͞�#Ao?.�	ƺ^9wX��nN2�1���+�ֳ)IB]�!�,��n��t�
�1���p�g��n�U�#�h�P7d��Ȣˎ}��e ��EӴp�D b�˿E�b��;j� XzX&B۷���M��<C<zЈ�^@�D��gf*�?�N�;�G���o�&OB.D����y �q�Ț���E;M��~�n�������PGA>$��{���.@	mJm���?	�Td:�a�w?���k�������H&�*����>���h�ՉsP�y�7�79��PӬH��j���g��v���N̟��ٿ�X
�--s�|S��B�Լ�@�8�}� ��%R�2��BC�8C����0� u�`M٠�{w�q�w=�#X|�jST�(ڸ]�p����h�/��w[�SG�$c���k��W(6�;�á���J����Q�C��rK(��f���b���оP����BŚET�y����OL2〆�?F�Aw��z�G��t7�iV�M��RX����I���r������r"�����m��ա5/�����/�Zn3LF�����hD ���BdU�8ab�+.tH���.=V��	uZgMLbdh__��u�ٓ#a雒��RTO1b��2[\�۸�݁*f)�]�&0�0c�~k|�f�k(l,�򃧫wf��Դ�JV�I}L�'(�Û0��J�#�Q޳�r������_DJ)�G_��4�S��Ap�݊��5L�������l.�(Mp���Q\�_X�Ťľ��:�����]R�E�a��JS���<��Àg���M��l�`.=�a���pŋ �u�7�hl��'a����-�W�23�h����̀�ZX[�k����U�;
�)��������)���m�R�o1�.&䞻o�Xi��ʫC-9ᑨA?X�n�l���g����[��N�^��O���!��c�R��d�C k��?F6�7B�݂�i(&Э�~mh_��JхG&@R�Z�j�@�V��f��w��Vi]�ݶ����Vqܦ@�|��0FQ�,�!��&B)�#AB�T�3��/n��a�|G�*+lҁN�nrjd8�gꆪ����r�[���C��0��C��0��1�d�,nht'Y����S�����7�$�`
�X��/�)��x67�#�Į��������J�Gl$\ ���S��-��jB`�/M��*J��퐟�&M�faH1��z��i�M������bk�R>�@���8�C�$�`�M����]�%��+x��.F��h��Ѣ���BQ�W�\y\w2�Y�T��+�f�xnǛ*O�D��'st�ƐNw����oPj@�r�-�9�p��O��ݍ�0��eY���\���Bo�ё��\�da��)���5�8X&�n��?ԝ=c��v������8��on[�d��va}l���1K��|�_���*���op��bn��L34CB�az�qr%bii�@`�]N��{ 	T�k��C��]�ߏe6���tzϫ�n�ktA�t�j#���WO�HcNɯ�?B��8>:gX�2A��*���;$Gu/�pcM����e�� d@�E�w� ��1#c������]);��5��z)o)�H){2"�[F#7�M&�^���(��.��g{A�^X��3��iD���ˁ�#���@z_����^s/���X�TD��f.�}Q��`c�B	v�ei�4� �ޫ_�	���=͝��΍�
.�~�r�G��,i���r�ܸ�@��c&C���>����+�݁�>z�D!n1C�z�-���vR����'��[-��],�ـcl�$F뎾9e�y�V��3����>�6��F�op�8�!�Z�����5���Ò2@����|<>�AƐ����yC�H" �@�&�<���K�)���Ʃ��Zx�L�2>ޗ����ltnʫ�E��5�p\�#�}$"�ԵQ �3��W�QZ��!�r_/D�Zq+[��<@.��7}���s/�)���S�~ac��{I��HR�gpz�!�UU|�Vs$5J����Uݓ¥z'� ���%�uם9��`�ն^�}���#j9��wq٫�V��j�;M��n�v	p&{�`�=����-O��[]t�%� ���;���\��ڐ���{�������g����Ǽ�kmܐ�sq�d薑�/X��p�yh2x����� ��Ȝ���f/)+L����g��a�?��?�r0ڶ9���;>M݂��wpS:g���(3�w�{��L��r"�r��.���?���p̶��%��^�u�)����5�[S��%�X����u��)x!��C��)q�>����{7���e��	���^4�E'�P�>�78�1���>[��K��W�QK��u������W)�"���M�ȳ̯�:C�0G��Z=�,��/n��\Z�h�z)Jp����f��ǿ��� ���;},�Ӕ�v3
���oc�� "�X���Qr�7>~+�4�2|�#�����ʕ�_���+=KxKO�0��nh1��j����FT�����
� ����%Nk�D�#w.O����&s��D�ņ)ʙ�Ќ��}��� ���6���>������ZD�Xgő�m�KG�d��ń��B�t�OE��1�EC8!�D���P����G3L&�:���qr�!��}Ʊj`�@�˟��W6��u�� �����}�n���Ϻ��r[&�D�B7�����/<xw��,���%�;�ԣ�'�٠�r���O�]���qO�s_�mp8��S�y�Ny�ȿ��9��aH̾�K=��lE#C����ٌ�-a��<v,�W1b\aݙQ��4��}�v ���{UG�!�Oɹ��9Ѡ�e�N�����Q��
���e�Yu%ƈ��i ��T.�7����j�ڧ=zᳶ�*�6�N��`�nPa(�Z��U�2s,�$e�˶��͒��H��di�'�ƅ�O�,�I�%���tl5�0��G��(�>�v����m"�$v	JZ����|;1}e~T��C8
p:�~"�д A�R;�-��S9]%H�)YK8�}�ن��� ��| �ТV0�kRp��o���̭��ț=i��bH��lUDԧ}Ͻ4d\:X�L��Ilc���r�*�D�B�,�*�+ʵuM0���v�b��vB^��s1�UC��1/����1ԙn$��y2������q�?� V*d�P�k }�B�i������u~�>Z��������s|D�3cى���J��ٿ|wPQ]�L��D�ѿT;;���_+�UU䬊���������{�Ȟ��0�T7���By!Z�r��%i�p\&�� ��Z���L�7k���c���LJ:)���6%�@zʊCI�'��2 L�]�֒L֤%�XNKf�|z-AxZ�Rf��9��G���)�DNrj9#g���6�DF�]���UAv&�rDJ��W��=!!�4��ch ( ېT�	�%,��(�>J�β7*��7�4D#��M�QtI�������ے�W�Y����[�T�U�v�3ƪ���c�&��v�F+ �J;���!��!�����s�U
hL�*�#�U�ww�_�t��0@� X ��nR"PG5���;��ARA3l+ˈ�i({�.��BK�^� ����s���2x�A�m�}�q\��p��Ȇ6@�bn�n�~�[�Kk������yɸ�Z�F*��	����_s0�O�d�r�qEߎ���|I����X�Js����o<OH9�	4��(N
��@~SP�i��3M�U2A�c��n�3�#ܶ�UM3BB/� 8a��_�������Kp������5�l�801H�AjM��;��ީ�'��t}�DR�6�)�vo����f��}��ԋ$GNM\����B�Ό{j�8�ћ#a�2n�;~�3?���o���}���ؕ�Px&U"ʤ7���E?�<���0Қ`��z��M�1]������n%ٽ��g��|���z���ɡ��6�R�4*Ms;�����v�����w.��q�J]��)����嚣ǰxK�1���D��.� YS����<���]]q�׍L��h�q�y��~=����fs�~|����#�����c�1�VX�ʑ�Vֽ�O\�3\Yj�s>n�Ū�w*�S�%��v\���S�ipu	]�v��;+(�G�0[$G���Byb�I��Ih��� �i흄-zbå͖�[T��W��U{-�2�v`]�Ne�|Bm�ݪ�D=�lp��������>�ӵ!|}5�o�1��ɗ�Y�)D~�+��P0�Rb���JӶ$9��s�{*���e6G������a�U��?T.�L2��+�=Ƚbdp�c��<j�G�14j�6o��s1��;{Ǐ���;�Qe����¡�R�I��pnG�����n�}$W*a�zK���/�`�<Ol�xgr�v��޳d�}ܕ�~�>�?�v:V:�T�p����I��;BЖ�kUYw4_j'71P�Q~ӛ�Ÿ[��L��8�����]ǎ+�[^p�}�B.A^��_���B�;P��?7X�lp즭/'A])I�n����N�.H%�����+;k\o���GW�ʶ��t��������O)F��8�>1�k�:c(��`��"���.k)A
M2�� ��g-�a"��*Ux��Aq)O	M5�~5Kx�l�/��Y<�a�y�N	��
j���'�JN�k���.É���}-)��~c��	_�����$����q��ȱ����m�t�R�����p#w8�F���伨��u��Hj�F�U�#m�3/�.��7�\J9Tf��J����͢'B����F7����}Ù{	sûp0K6�1Yl��;z8���>�����<!/��B���-�î(k2O����_������U�al�z��6��,r�z>�����:�z� %gʇFۿFF�4�SNTqC����bNN����Y�w���  �@�0±W#�A��&�{_�,2S��v�u�R��N[Sܬ��L�L.���jVV�j4���Ή��1��HF|'���P��A��%��@f����!׫�Gφi���͸��2���z��ە�M��-��F�����ҥ��,W�%6Z~�F[���w��ѧ�lv�]���(�<��խ�6��.�-�c_qD.p�
�J�HH�he�	a���b �r+��R;��NZ��fT`A3;��M>�P���W�u�4�BE�u8js|&��i3by��_|���k?^̎�]eH��#��=�1��ȸTM��E����&&{��* �P���T�����b��]�̾z�k+{*j���(P;^���z�o �T�V�V�N�B�%\�T�&4s/hK|�S��o0Q��F���6XN�V?s����-��:ha^�Y�@6ه�ǃK9)�\Qq�&�\ix2�A�F[�*Pv}p�f�߀-�l�ݖ���
3�wϗ��^]�ܶ��Q���[�� m�����Q=VjJ3�-m̺p� #�7	�x��m�C�-:�	�e\S�7�ɐ����"�:F������JO0P^lX�
���IF
����5
'n�Z#+i�޾)�B+�|����]��S��K?���Fuj��ٞ01����L7lj��d�9��ٻ)����k~�!�1r�k��RE����b�2��[dC6���gU������>��μW#C�bы�34���-\�錃��	|� ɶ4���WCh�yؑk�V�y��*
'�<ط�]/<8r�A�h,�مK!//�a�>����4N�H+%-Cx�!X�,�H^���D�����]��%5|:��H}�H������w�A�.ܲ�J��t]�X��,1Aݺ���.Ha�.)�rq�_T���x w53S����/���I�(������("�����M�6��_�������Uc�/�N�+�����x����T/��a�Py�~&#��g�D�d�B$��R}\����d?f��P3�o�I��#}-�w�/���ty��0VG1Z�7U5�¿/)�[�7Ş�_�J��h찔Uֆ�Zؘ���Y�W!'y�XV2��6f��|7��a��	La	����n�>85"H���Т�w>�����8��������7�ub&�2�tC(j�Y���A��%���6xlM5�!�R��Z'ei⿂�@��	�q��rFq���Nv������K�l�ڧ��� �t�qu�����,3f͠e������x=�� V,�C��۹�Z]���4G��J�z�Ŋ-�M�@f	���X��� ��3�6�����=4H�,B�<�&��"��|�:��F8��*��|��e�����+���xO�tc�{�>��??���#±lEXl,3S��\���|7�����A����E�ű��'����/tzڢ�'
���(S�[����[�{��KY�s�*����ۜ1Y(�}�HO��̯�BfO��gs����/c[��!�4+��h{�5���
\�L�9�n(�_in uħ��%d���eN|i��f���iH���FU���es̎�}�_p<��48rxO��Æ���f
N9*��&J���YC5��[�qm���}�|`l�Ƀ֠r�a����6cI�"�@�������CN���F����}��lŊ�鸴�Y[�2Lc�B����7���B�u���aS����KO�!쐛�#S�V�4�+��c�����!�s6JMH`�P��J;j#��Ǳ�r�B�������$c��P��:�^{\^<�+�چ΀$����f���5���y4���Yr�Bi>����JI`K�*�֢l3�AX]Fz	v��{����A���ON0Ϸ�_*/-��.�y���h�x�
��x���y��0���V}h����VN��|�;Ȯ��Xp����i���#��>n��CP#��7 3 P�qn2Z��D��4G�G��u����p��k�0CH�.����gQ��� �r�ux��d�d@�$b�qA�������]�E��fL�=s˱%9�#ȭ����L���;N�y�"�����ܓ������4���'�ē���s{���O`�(s�R�L�s2�@	{j2�6H^�G//W�	E>��*/�9R���)f(�9�a L;������uh�{1�nwA~���S����BR.i3:�ŀ(R��-"T�X�3��-�"*�u�(�̦�l��w4�ym{24*ƅ�>x�B6hխ۝��m��\��+#cZE�Yl�O�6�)n��I�0u]�az�9M��D�?JX���,:�>q���0ܚ�bw*C���
be��E�Fli����YEss;�P�k�ܶ��5��J�����LX���IU�Yᢷ���gB�4D��j�����#Ո��օ?τ^v���Q�9��ٗZ�1��J�F��Z���B�
��zr������U&�jŬA��8���&?bh�_���/�����'�N0w�L�K��+��֋qO�����T�{�7���e�aO{Ne+��v��p��Q<�A�2��A4�Y��j4�iD�k��$+�c{,E��_�W�0�8C��H�;�e�a��� җҢ撣|��"����^HA3�kE�݇q��n�~�@z＠�G'P�R\���&k:����.�\dKy�Ѐ��m�����lL��ܗY���X�KBusW�� �e�!�2�7�k����}Ld�0�E��Wx����q+�/aJ���m��kmUh�SZ�=�wK�,���=�N��y���i�SA����S� ����I��!dDq��4��nB\�%�8��R@��+o��]��,"��io.ϲ��]��һvԧ���Лu 9���i�F">��~S���t�܎5w#h�.��/�q^:���.(����;	X�;?䋥�\A��v���H��Ut�re�~�i��W����MΔ9�s�~���&��&��|���{��bM���2B�D�L�������y����^p���ʌXBL5%B�+������ޡw6������� $Y��Φ��όdns7x�1*#ô�ͥ1�g������9�"Z�-�1��Z슣AF� �a�?�E,T�v_kDn8s���ޥ��	��L��t��,�h�Ȟ�����B~�6eT���g�΃��h�^��r�%�.�|;�(U�3�����]�r�M;r�f�{��BإÇ]�w`uj�G$Vg��j\PӃ+�g1,B�S�>F
i����������K�}Q 3���[�W���Çv�������b���q��]X诞����]9��B�5�)"s�R�}_M��	)�
'F�pM������A%V���~w�4�=_3�h�7ц�w�y�F�̖� f� ����z���E�𸵨�1�_���).��d�+[�b�d�n	hL���$�Ә6By�*�֒(([����is����$8t'
���nW�G�B$��8R6+��L��U����-Wʏ�K?z�'�:Zj��J�&}���ߝ �hJ����!�c���2�l�:�ie ,B�S%ޕe�}c�E2;vK��.J55) ��RF��|�o?f�i���ඩb-mZ^wBՈ8��s�b8ezd�G;:ا1��$����+z�z�����@�c.ׅ���{4a�	����� ��n!���-.���c�7�=Ry���˹T�<8�<R�-�e���@�~
!�xm�V˅Ľ&_ ��� ��<���mv��dǹ�;Ji$Џ�
�n�ڢ%.�hW����&�H0^���1�B�@nE���p��^J�� )LՁX����O�i�[J�<OSFtw�����-�R�j����-x�JU+^���_�g���|x�E��� �v��5'Z�%�12��}#dn���\�`/����/�L2 ��OT�J���2&�~dN�^.��@i9���Ű ̭�ݽ����߁檶�
@>T��c�ꈚQ52jT�{�t�EV
D��
�G�u�1vfez�_[%����ɮqH�y��^cGLݒ�v]�����WD:����oO���b;����xC�q���Zj��j���O��6RC_���`@K����tu�	u��$����ibU��p�)ә�]�(��ws��ʖ�����?��^K�
�f]���x�G9�B��6.�)&��q�����2���`���l���7������ t5��`�B�+�A��	(�!A�����E��E��ݿz�M�9����8������T��'��+��d�,�i�b�ظ� zݼ���`�}�I�}����z�cz�g�|��V�O0�M"� a�A,y�ZXfPl�lV�������J���_Q��/M�'�Sq�Ṣ�U?�k�u���5�σ�[��>�6ٴI"�)Tb�^c�д�O������?)jq>�J+E~��c�7U��5[
��uE�[�_:C߾�G��)����e: )[�V�R���94 �F�2�Eʂ��`�a�.7�;���~�M'�;�H�c�E��-�r^�S����; �^�CJ�wG4Q^@�>������Q�D����x����)Ľ��`�[���go��ƹ�`+/./4�`��Q���ܭ�QQvl>�K�#�W*/����'�� ���/A�ص.��pw���lj�g���;�f�6ڨ-��5��B*4����~��$}=�PM�2]��¹�G&pZ^8���gỤ�E�0��I4��?�ab�/���)��uߤ���zh9��~4Zf�k�W�	G����Aw���b�:��Q'啬y��mr99�"5�o3\s*����.��
��`dr�y�a&"�C91Wu�|}��§cDAjZ�%?�=��*��T�\+��|�\��G�Lտ�-޽��jd�xA��h�l�i
�T�Z�e�6G�>�O���F������ au��Hļ$&G-|&���;r��5��,9�+j���g�P"W%���U�a�dM'���?��ՙ\�ٷ~��,a�R���u]�%vu/1~����:�;Q8�/6�}7����ZL��i��e�Uu�|+T��G���wMІ��R�ⱶ�Ն�(�ǭ��Y�²Sz���J,�Q�t.U\%�Ǐ�ACB�^)�'��;m!C�1�E�lў2+4��k}���A	�J��ʶ�p�梯�ꮼ���g��l�j7�m�i=���k�Ĵ�+7
���$�a=�`1k��~�i�}���<��/������_�D�$��'P���"�r��`���	��4�s�~����>h��G�7��(��D��=�tH/�sO��~Ę�x�1|ޥ���Q!���E�*\�/d��De�
l���]�*g������B����z�h74��*̍���.G�Hkr��v�J�k�(�`�~�Bp=�
x�}��j2�w�P,۰��l��<�t��U��q�=N:BU\�\<�>�?�.��b\oZ*ON/3(Qc
�2,] I� ��X����6��[{+�FQ�G��}�����?<@K���X�������v�F��8�Z	k`=������j�Շ?Q	Kx4F�v�^�n��{ �p��'�͗�:�Q#��%޼��!����T2�(�^Ẋ��I�p�tz����Ő��p��{�9��5!�3l"?&�E:�����Lv��Տ�T���� J(g�{��&�%T�~��o������6e�o��&�@��<�-B���Bz��^<�?��r�a�j�L
��}ö�g����:��ջ}��&
�����IX��bP��}���1D�$�;�_���3bS 0�����3�o�l:Y_�2H
���A�b�~ME����mK�`�� �
m`�y3���x_��nq���
������Z1�?�
4�q����%;�����JiJ�֌�����/B��n��]p#�q^�W=?��+�t�ե$�T��KO�Գ4��8�p��,���x;����'�˅��&�H��L�j +h�دO�D\�H	d{1VDH~����㱙<�`!t*���'�x]6�4�Q0ct�[�"��Y��[���<�rr�`��7g`��q����Q�`�\�x��j��n_I�~w��D�;�n~����=��V�@���\�i���neUnD{>���s�T�����:(z�`���)vA36rh90oD���dXMƠ(���-/h%C�>T��u���;ݒ RԼ="ˇ�#��5-C�qvk����2�@�K�*�H;߽�EIѣ�4kN�B ߸7Y9����֌�^:���q���?~�q	���2#�&���Ҵ��[�T���s�w
�b-�%{;�.83���ߢ!�l�B��bQ��<��צq��Ӈ@����j]p�SUi��S�ͨ௞��	�g!�\�v{��|"X�!�~I�����Fj~�w�k��T/�A�ٓ�76[������R�6��|�~l�+�`�P 
���cz���J�Р����p��C?���8�f���Yڞ�y+�!��s�uj.����æ/�/�Z�-�L���	��}'X�:�j�yW3���I�{6s�>o���� 0�IM8f儡���,��k�>�tRBum�$�Ðp��$gt�% `�/�l:�u�+q��J��]�E\�&_G�O�fqDx8l<���ZX�8�����JT���y
���X4����xI����]ĘV5��2�A����+/ͯ�4�M���W��wՂ��K����j��';7/�:�uX�h�6�h�+���ø�0\6H�U(/�Ѽ�?����:���a{��!l�����=�6{�"���l�*l$�5˥A0��I�W����30x�S���#a���7*��_#!vwQ�O{�M&Nm�'j8Sc�p�]���A�.�y��QV����C�vt�t���u�"�i}����J�9pe�H��;6:+��&�r3�Al�>��������=�G�Il�Db
��=�ݧ�?$���5��c��(���'���?����������'�
�����p=�)o^�bҠnb��9C�	"�ǔ���;,N��}'���?��ss��x����Ն�0А���I}�&7u�Tlj��I���V`�-��w�N�6�O#�5K�Ѧş��Ld���"Ω�#���!
ӲA��d"��!UI�떯(�d��4x5�g��g9%@���V�9�J�E/s���b�3�#8n�y�?�0���E)�)�	w���8?-þE�a�‶�=V��As���8j����Oq�������:26�f` ��,v��y�I.B�}�-�@�t�l�,�0K�B�M��hVy����|W'MФ��Bv�+X^����-'�+�n���B���]u�q�q�]L�������@`�;I�P3x
��W�4�C��L��!��:%v3k�𖪺��C���s����e��٩ڟ���o�3*��83��iem�[g�/�"����pͽ�Q�A�T��[雝Yb	�fès�����u�R������S0��{�!y��Wj����MT�O�U@PL�3�m-�<C@��`��,���;(l��Ͱ���f�
��,i�|��7;����/��(Wd�N���f�W�DY`��n㽣�$��~e�9�����&��b�k�-�F�a�`�ݨ��?�T4_ݬ���!8�/]Mi8�%�;�+R�UС^��u����.�zww<"�D�M���r-UZ�U���&��^,	�Y�TĄ�r���dA+����G�	i61�������c�M[z�=5�Az2X�r�0��4��o�{���7oyO��,2�	�F���D�\�[�	�-#�z�֮��C��nq.L>u�G\��b+ט�o�n�����ݫ-t��0��-@���<��Yh��^�`ͥ`�*@Ѕ���#'b����=u���GZ���{k��'P�u �M�٩)�F��X-��?8�?���GO���=M{Â�y(t�� ��+$�_Պ��x	�%[0S�)�&yXS/�մ>v���\��
?oe)��)�iaP�(ץ[rG��T��E��V����(�AQqQ�2�`���/���7Qeb_��&Ny%�l�V�� �p*F��CED!	��8�HF8��5�5a{%V���ϥ)���D�~��@KW�,���G熑"�F�5ԩ*[��5�	^���ºV�����L~�\��Ӂ��4��y�tb�S}S\�۝��+�\��E������AJc�e���ca�}�䊿o�X�q@n�4Ƹ|�T�kK�^4���Q��i�?�b��.���;��6�zW�.��CN�����+�f��Q��5��k�ss�Bj�����v�E�� �'qX�[!�%p�2g��p&�����&�-�K�V����R3���ް��+N#���7�D���?1@7���Vg�"��Q?�$�Z�$_�(��x��v�K�-q�1�~A�*4	�P�~��у*-��*V�<O�����<I�KO�AT�y�#�2-�
��"D�}h��RҎ�~#��6X�3�/�*�`k�*���2�x��L�p'�yY2��t$�0W.!K�C�w//��}�y=����jx�2Y�}�Đ���W�Bu
rxΫ>"���H ��Ye��`'����F.v�P�6�����*��
�<�"��p��;�A3|�'�|�H�B��t��<�M��s݁!��d� ������VT==<���2�gM�Z>��*��9Awo�=��bj�!4CmD�(�Y���?g4͟�ϻa�mK�"�<u��K1X�toe����H/�lthZ��j�?d�mV)8�E�6q�(6�%���"c'2iU��A�殾��W����W�&�1>�����$o���LB��8��:+�����˦����A}<18ҿ�o�n�I��=wo'؆�R.B�U�`��b��B��.���me!CaSJ�*qE;}|p��d�7�.2�������RG�u��[VO�m<b�}'g������МXI�$2p�T9z����~s���)[����3�^��;��p
?fPy����\ˀ�$�Ø7"���[6�Z�u:��e֯�?�W~+�,iG�QP��
��D|��W4�^?Ny6A�$O��+1/���d����.5��߉Ao�,:��ʬ&�.�u˲����d������F�3����������1��s>�[��W�2E�G�NusѤ�8Iy^�-�qg����iq��TG%/(n���'�x�U*ſ$,
���Q��s���=��`d��k�;f��]O��,���5ġ��Mo�R�2WVR��P��� ��]�l蔫f7��p�K��g ��.�� =!�Y�x䬴Ž�;��0t���vbhM7��8���|<��6A:�ۆ�s65�v,���WcS����������95,�qB��a��Bl�%a0��q{�y��)��:~! ������GE
y��L@��hT����QM���K�Sq3�f`��1�#�%�oÄ��x{��1�s�)�y�rq������+�!E3|�Uf]���TF���mܙ��:Y&9'G� @���<��)�*	�K�y��Ø��)�䌗1�4_0��E�J�l��>�<���g��VSP:hX��o�# �wT~|7�+�N�h�8h\�����Z��W��E!�˻WD#Ԙ*fE��fq���-��M��C-s���2cf����	D5����u��7�wAL�X�t�1J�*��jf��`;S�=�:���.����������s��^>W^l�xQ�J��!´Ym}���Ufo�>�d�Þ�I2�Ķ�ס=RAn�����Fad)ڳ ���s�b)���9��mY=������j���[���*�e���0���3��nH�5HB�<�<H����$�İqy��}o0'#�=÷��2F���H����t�BΦHt�nR������� ��l��A���AO�$����%ϐ��@t��{ơ�� �oH)i ���0e/��A�yv���Æ:��t�3����aBއ�u�h�,��`�Ƕ���Pes���~F�,��dv�_N�Fa	ޛyP=����v��5�,8�O^t��\7��視��GO��P��γ�E�G;��QA�%%���� �L�a��2���u'p+�M�OwF	����6H�/���QE���OV�����Ƕ�_����r]A�w��7�1�^�@[~�ۇ��p}h0_;�SѭG>����6��cėr0]�R%-��%g��йeCNK���Lg����QSv�eB��뽿x��r
P�+��~x��IKR$��Q3�K�&f��>�3�ROHN��>=N�gq�N;.Z%ց(Y�=�+�*�M��sR�J����`'ρ�'�/W��-AD����;ى�@����JG�dN��S8��۱���MT�'Zi%G)�;<{d���X�!O-�d��U3S(>�%
����B̰+�^�k����{�x*L�������i2y��n5��ݎ��u���*�cm]��*'W�K�!�OB��[�a���K��"VP�n��@w��@�g�{t�U��}-�895�e���
Ce��E:n �_ rx�1 ���7d���^�|Y����h���+���b�_J�P'kv4�d)#D��z�0�ڜPg$oj.�"��q�R�O�A�bKެ�̮ʣ��9��YC`F��:�4��
vK������Y��9���}DK�׫�l[��*l`B(��ҠfX#�7�W�\\���r�N�8��P�B���r@��΋rނV����Jb@����don�J�Q��.��[�~ď��'b� �:yf�S�/�H��Bo�Q;�|�]r��ʿ����_�D΢�m.ߜ{G�8{��a �|�y	�{�ڒ	Z����ϻ�]e�uk�6�X�w�n�������S$\���sd@�V�-�x`�{�Y�E�c�WສS�%�Z��jR9�FvdV0��&�@����m�K��-��iZS�V��>���IO��WӠ
�Iwg����t�_.%wH6�#���?�'��^o�}��q%��	��5Pb�QN6�v�ڢ�2 v��Wɫ�y���yr�ڇ~�
�v M�G�Ҭߪ��w��=��T��{N�w=��}ef�Nf�Y,��;�0j-�����.�*9!1<,I*,`E"=��l�h�H	xt�����2�s1��M�OvX9%A��B�V�蟗��ʏ\u;S����S�h������f]��d\�	��_*��WD'�������C탮_iϘ���Bg��.~�X&t[\��&��uc+�s+��h��I��WӦ6�x����(E�c��@��8����ƪ⌥x����+��E�[:v�H��l��NV��YQz�l��{�sC��)�%�,C��@���B �Q!�	&�6O�7Uq`cu�U^�a�=�{�$E�%+�9����đ��z�,�u*"c��We ����)@�;$a�3N������\�K3�a��.��`+F7�eҮ��g�p��0dr�g*f6QƜ-�2�QŴ������Oy� ��]n
*G��Ac�w��YMx"AT{*��[#򑯦���Igٜ���9=�uR��G�!'�{�	93$<�7�#���s��K�~��;���6W�U�* y�L�0IMqBCp�H6���������(s�/�?�Uk7�����U��1N�,���Aإ ��O��f�1���#�BLAk�8��5TR!�u�\"��XJ�hQ�<� �Y`;G�
C%�����9���$�p<V���:��7�9~,�&���0��h�K�W2�t�n��+5��A���4I ��MZ�-3�nm��{��|�]��a�+����'�Kq5�8��{ON_��"�Ps�\��i�,��g��eR�c�W!5<���٘�q�q�>����M#|;�%?��n)�����'��H�5<"��;�]�+&J%c��ݺ�7Z��yL�{�+�H�&�& 6�㣋��}ޒ��t�`�"ǹ�s+���]�>��9�nw��-��mYp,�݌��Ŏ�,���P�r��$���"���7�@رmdOzC`�����m!}�Q�J�L��{v�B|or]E?K#ޣ87�8�E[����L� �1�c�g���td{]䙝�o���� �ª7�{'0κ6����q�[�7q�8�	K�g�i8O��o�>gh�uk��{�MYcp{ƒ�P& �&e^�0zJx��OU�2"]=-2o
�]`w����U��W&C%U<f!�o����|r{2B�Ǫ��?�::�E�)�k��-͖��0���
������gG�4~�D�n���|G�������˪�:=�V�x��H´)�K|24���)`��:.�mk�@�~[L#���wNQ��v]�n#&'N�˽[�߸B����<�	F��G�`����5�8P��?�C�՚F��ϒ���?�z�LPf����5����V>�N�;��_�d�����<С��\�g/#7I7�[J��|X�[a?�{5Ҭ�4�2xm��%�N�9������g轊	:iךT��uY�	V3�Y鍞��p>:�4#���}e�V��(��n,D�'D�y)L�����T�i^�b)!�	-T��S�v�:�^��T�t���̩���7E�q����33�r��Ґ[����fl5@�6�G��$��R+m)���y5oG�N���n���]R9	�����.Q^�@�v8�����B�)9L���U�b����wg���kB����I7�-͗��%����-��8ͅ#X#܊���;�]S��=r[\��j��v#^��E�Wi�"O\^k9��vG����E��u�6�-P��SLׯn��:���Q:� �b��]�a]����s!"�i�oK���t�,ń�9�e�5��j�g���Y��yi��9@�2���`�vt�i���93�@�A�kQǑ��zK!ZQ6�#�W���Lk�>�nVu��e&i��8�:
�����0�@�����pG,�sD�������H���_�5�MF����.:�����^����~y�!�B�+2/GB���>�,��{Q�̆ޕL��;���ӟݗ?��1Y }0��Y��K	b`��"G�F��篣����h�'��y�.)���5�~�E?�r�a�'~��bY7
n2��v�2S�)��b���1
���I��b����<�>|ˡ���<������,mm`��$�ݫֹ���
�L�p��¸u��Pm)�X��_��\���N���Gvݟ"*��|	����kE	}'y����􉁶Us����D�C";	��K<��JV��G6�i7n�i*J/}�t����eʂ��ᱲn_G�Ǵ[Q@�v՚=..+�ya��8*�)2��Z�N	.��r�ق_�Gs��	��K���� X�]XbL|�kB:��p-HimT�+�Swڼ����"w%1*{�[@^Y�	�:�������Պ�s�J$�Po��G�R�l����2�O�>1~�wN��l@�sB�r�7nm�P�?���꓏���9f#������3���|���&��D�@��+�!+�w#[r�~���Tq_�pvk�)�֮[T磣��9���У��L$l1��űݎ�+L�@=�o���E5�k�����o����Xo<,�p�G�k�o��}�E�o���gxG����DF�Vʲļ�(h|
-�"�'�R���$M�����_�ٖ�4�5|}M���R~V��/��2�\^�����u�fg�� d�T���/ߝ���L7ߛ�yE|g�+�t�%�yW%^A\�-�ʨ�(�nw��������%f���h6�(P�r��<��@U]tVn�1Om��Ԕ�辵���	͈9k�C���P�w�؂�S��v n��lb��ν��IS�#�NY��
���&G�M�ꊦ����V߾*����T>��g��y�08I��v�@�JJ���� {�q���0�a�T��^A����\G�� ���x�^W̝�S�Yn����!}�)���dc���h�k��m�5t/�Q���J��~NFρ$���u��:�`,��eoV[�ZXX*�A���VuW��b,9�Ø}+ǿ��J�x_�_�&�9���O�����E�꺬N�=�K��E1)ŷ]
HYP>?<�C�v6"'Y�m��T�����
@�����3��)�z�$r���|H�l�2ð�����Z��������}����-��*�㬡��Cb�	Ŗ��4�G��./��/#$��p��jSd��q�DX��Vk��>Q3
%��X:a���]e�����X\gG�E�[W���.&�{ܠ�̖��
*W�q�0�2JVYjP7j�"!�`�LB��8Eťq.-�ϱ�RR+�Ju��e`�	�R�h.�:}���ϊ)Cf0W���@�a�_��8��6X�,y5YX�|+c�nI����KC�T�
Q$�Tۜ�ѵ|8�X�����Nuʍg��9�z%�6�S��ײg��3�M竾H��ad4�=;�I�r�m"=�ˣ+J�Z������� :��L��|\�楖��dP��9�F�h5/_�ܟ�Qd�����&'\�RL��Ʊ�3�b�_���g�|���u��C�� �Ǡ 0�h;�6��-�)��Xy�GA�?�S��7�����8'S�����u��]���]*p���.Rӫ���i�I�6$[����?7r[�Sf� �Q�h��NaC�w�{2�]0�yiӪ�p/�r8���=.�c)+��	�Ж78ҩkL@1�q�#���d3��+�]�U���F]���u��1��}�cj�ѓ�ps�b�`;h	���!��B=3���հ��i~VW�2e� -Џ4,�f,4;`o^�0��Ե�kz����#�W}?1̷C
g���m�I�*��I�-�~4�%3�)||f�5�5X�u��a� /C~�b�^�2"�.��0�Fˡ����"�zw�gt6Z�>L	cS7?�Pժ�i��t�i�c����f�*_伥��k����������{mn���L��E�J������Y^�,��g��@]ށeK�����U �c<��Ae�����IaB���wn��u�*tN�	fl�����L���-^unXч���"��p�Z�|]�ߦ^��,�}���px����*K�N�Wc�&=\�;�
�8%���PO��۽V�����b�[����8q ����D�.Z�$��N�>�b����1u�BƼ�[ͶV�ֻI�[���t¿0����t��&�k��z�\�f��*&�b��ĊTRқ�$���� ڈ<^����w�DX�sФ���p��5X�,��N�57�|��lP��`d(�v!�GT��%7J�M�~��N<=�%�oD�:����Q|�I�s�6d⥘c�Lկc��Z�'��j�U�5kT�?g(��x��r*c�����g���e���0��F|�d<��L���_�V�t����y[�V����q���'G?��ZMbBtv]�&�Zp�dW����Z��x�]�+��I7"���q����>�8� txwSe��Q�CXܨ�
����H٦�[�k���s氫���5>��L-n14�?iy��4S"0� M�p�VLҜp`Լ���U�>:[�����a�	�;VKI�@e��y��NPr���g4�u�G���:P6u�	N�j��t���(��J���E���)��.~��OpeJ~Dk� g����4�f7^�%��L�Zo���s�:#l��
B1���MY�����������#{/}��f^���D�3��c���Fxg'�:ȯ��ZJxy�5�Fo���=LA��*���@N��Z����A�x��~` ���:������~��+��=���X��=&hy�Z�
�$QN�JdH8�h������]��O���c*�r/N�nzb��hN?��r��c̫�	>
�Vo9���c��Y��2ܡsQv�;S�����eaV�~�Yit�X�k���w�h��+��Á��i�VjXW9��G )���S6��w=����f�1�t�%��-�s�Pkp��-�H�2�T5l:	�����꽹�0|X�&���f�iF��?e��!e;1"�[�����*yO*<`[�力B�����Q����9z������YᏎq��bi�(��<A�M0�|�����~Mm�Ka����̨rx�/�g-c�ț&"��m�.�,�X$}�n�"Y�ocLF�ɰ"�Cqj����zijN(F���h�I>{�6	s`%�JA�V�1��%m����7@x!h�0����:�����;�����J߀�)S��@��4Y$�u�Y�$:���
�umx���Au����G	4�^s�i�Q�l��"�al��wQ*�A�w͉A��*�8��E�H�	XRM�
K{���wH��w�.�=`��?�m��N\����i� ����p-na;��s��_��
$�
�����7��������sx�V�ͷ�
�k^~%l\-0E����s� 		�zƄ"�Qċ$����˲��-�>��f�<G�b	�&)<����þ��-����R@��p45���~ͶV^�;zO�;@��xnb|����M�$����3|F>`�soD���M�g/�y���h����oq!�F��A���+PF3AR�8؊֪�6h$���;��_d:�z�X��٘�n=��6�!s��Hr����Z�8��#���cs��.����,��OȫM��$\�6K$��\H���5b!�QM�?�h!����$)�ˆ��#c[�L�ҙ�*�v�z���[Oy�!>��H�Q�TN\o	zh�{���K��������Ӹ=�g�c�`8�r�zbm���=G? SD�x\�"����S������k�p�+Y�����Ҥ���
Q�������{�<�s8�,PG5
�Aڱ��G�G��H[���S�f��m�V����x�,¸	��Z�^,e-���C��N�B���k��o q����pC\��&�k	�E4��JRD��ƥu5���}no~��htae�Y���۷���H��N,(�n�nsA�f�%ɮ�a=K�~��W�dfmaȯ�g��D}�G��ת�Xf&,������qZ�x\��TZ�2$�w51w{㞓ӛ?10�T�J:��jԧ�.�,I���@�2�+L��uEX�f.F$�t�t�@e�,� �K��A����$�X��gi79�ye!6���u|��ϻ����#�^cu�!�.0/R�,r�QaL��:�N"Ǒ=,�1�BDC��Xߖ�C�s#�>v��qG����R��rαl���-
I�ۖ�#h�JY,��K*�=0�2C(������;�n���� B��`T��h�����prHu���������<��V���$%�5Y�4�V�L���5�x�,���G
�j�D�i���4�1��ut�� #\����'�w�)�CW�o�*�>-9�ZZ�J &�<�����+�pՠ[�|�U�$�s�ì���R �� ,4 ��a��{��і���c��J��	')n�97�>������YmX+�]�R�z��lj�&6X�KQ|OZ�Ѭ�Mx~e���=zN$"�	�e�+p$؃r�Օ���N��V�n�f��;	��|�$/~��E�`-���e���j7�*�*Ŕ��)Jc��1��%�خ�3q�
�P]�)U���mo4sS�`������?Q �=gn+���)2��+�sB����dV0�S_U�mK���rYMٕZ��d��Ob��i�����l&Yt��%�f�~e�0Q�PN6���[���ĩ���4!W'D��*�䦉�$��|���W���$�8��3G�R�g��n�axE��g�h/�
.�s��D}G���E	����7}���Y�A4�j&�S7^{����e&��b��q{B5��q�y�s^{�-�n䚑�%?��o�!�J��͈Xr��iy��:)�Ex�5�^V�=3���ۘ��q�&nb�~��i8m����
 [���Gyo�G,�4�>ٝ|�H#��g�l�X�� 7��n2���rVӕ���|�xY�o�`*:w.�w�)��|N㊢8V��3����K�̧7�_�^oC������3��x3�>/i[�Y�ϐ��eiS��(�w��.��Gӯ�"�W8&6o�,���n�cT%7T� �B&��x��i6!��#�G���j�.E�P��l+������d���{!]�����p���eO~Tr�]�L52$��ԕ��F��|\ښ�uG������r���LQ}���f�8�ɑm!���/t�`�B� \��j�!5�I6�{wF�A�2'z��r�o���n�q�s^.���#2�f۠1���j���.�zƴ.�]=�x_���ն`�V��9��eU��l���Q)�T��*�
Ճ(KH� ���R�-V�V&9���H)�gDb6�U�B�%���kS�95/Q��	����mo ̰��2;��8<�Zœ�j������ި��S�Lx"��ՇG>�K�MT���ͼ�vns�5����\�^�f2� ��ǐ������Lx��}xr�/�y*���Q�9�M�T1��מߏ�C��8xqV����g�/��/�f��!�������*�T���I�T�t�N`�����i�$��[#�@�`�\��� ��@v:�7B����eӎ�3��VG��,�usv�x��������}?Hg���Yń�l�<+6?$�p�1o��I�2.�c�-��X/&j�Zê���`A���c��vl���1��G�֔�V���S�#[>�� >.������J=�N���UWrl&�E����H���j�j�ȶ�咴�,'a�I�
@6�Q�oȧ�1���ipZ/��5����8�����I�Ǧ��cb$�r��!�9�?}]��)>���b��=14}IQ=f��m��� U<F����D�<�bT|4J*��4?�젹s��f�yr�:l�"f}Z�R�_��6�dh�й������Oś�
���E��OH(�	%F~kĆN�|��X����w&T����F�h3{Y�d���۝@M4�44�#����=j��y7��F�iޝ�:2�����vm&�z��A��c��ݑA�<�����劓�N��$d��WI�`������:��h-��2�Tk_[��H-�n*�F^�q�Z���f��b����Fj��ϲz`_ڎ���kU��*fWu��~�ӇɃE�:�r��I�����h��~y��:��������:K���(pg���{sy
�.QY,�&�{#{���N8��me	�ڥM\𒰴p���BM����1����G�蟕�����f��BcI&sC�n�[XQ2v�l��~J����3��BMT�Ҡ�Q!z��{Ep-.M���AAE��#���w7Ьe+*\���Q2�������9�H���0��g5���z�G>�{#4Td�2��X�mR���&������Bj�2Հ�����6�ۑ�Ur��T�US�~��'1�P⇕ʶ�[Sg���ܳ�♜"$bY�Tl���ȩi��2�N��n�vC���^�v���oLƑW�������rI_�PĜ7�#��aa%�>�{VP���04�L7Oq�<�����[U�7����o@,�uaa��(t{�e��C)v�+�tK�$߮�q��z�GxXhQB��BO��5z�1���K����05��X�nx�oޝ}-VМ?�D~ᰗ]597�.{.t��Ԩ�и�6i�z
-����Lx\(���J�VC:�o�)�7�1E7ɵQ�'�;�������>a�z���Ht��d��>�(���!���>>�v�%�v[�� ��ͧ�^��<^��?4��.�|�v�&	�!��oF���{�xA�\I���Z�.F�$���Ǔ�'�1����d0�׾�k���C2Ӵ�T�<��t(�~XA�m��7��v
6�n��#Ώ]Ŕ[�y��f�]b���g^�ԭ>������ʻ���$�	ZP��h�,p�2a�N b�1)5[	�KBet�]6Bw����c��߻�|�d�e��3(�{+�P�(�����	K��.�g;¹x���rl	P˩ǝ鸛z�HBh@�$GDD�l�������dW�r���w��o���DL��X��qcA�h/V�����F>	f��v����U�^`r��F�]���GyuY���OKw..5��+�"�nc����O���ȪWr�%�\�Y�"�'�!�`�����Su58�"�I����*�S_�����KϪ���+�� ��:�O"�
][��0װ*��A��Z��4Ұ��[q\a���{�J5����O���gT��5]��Oש����j$+���7��Yi�%i��Be) ���
�­P����]:\g�N�G��w
 �N�恛�iM�Y�E�T`�eҺ�Z��D؉`��~������b��lhr]q>s�����Ɍ�z�H�^�r�����u�����QQW=���'��Y-1|�2c���`��&����|㩣�Q��#���1bY`�%"o��Ҡ`bM�H>��Ai����<��SIbVѕ����صj!m|;��@fyx�F.�CIV�pP�.��?F����aW�:��<��}�����~��)�-QK|C�#�_�O�3ם?T�5���k���s�����bY�� $�������]���';��.%���a�����
9 F����RI� �X��ɗ������Q�2�l6����)�gi2r{�f-����&:���g���2�@�q�}�Fشr�B��uͷ��GX,T��Ҷ*ܧ���>-U#�����tv��Mj)0�����BV� KZ��C�g�Dc7�����?����^�Nԍ�k3n�^���_�QZf}gk��ݒֲ`:�u1�)�ɣ+�>�S���bcF��S����޹�A�`�1�?����\�0&��~���g����%�X���T��թ��ide� ��bU&k6���݉o��� �fX^0%����6,�PtC2�`���M�rM��W<�-dzS���66�'���a
�͹6���K�Ė��V�C/����p*(g܋�3�P�����5(�ᒪ�����A�3��1!��J�{��)oF0h�6i�����9.KG�.�?�!@E_�Pm�42ۧT�*�<�T��71z[���W��F����dIC��� _��i���IK����ɦg�$i���
)!��?`ؓ��������f�q+g�&���������x���]��PA�%kh�۸%�j�l�1*O�HSԘ��l
ե�'��YC̩�+�$'�������������ݞ؅b�~۟H1g�E�(N� ��2������BSC��C�j>����?u��s3eB�b_Me}����
yk�MJM�F��ʓ�ԡ�9�I	է7�?�kI�L �����9���&hpV*h��ϣR�U-�5����H�md.%s�����L]�i�;�c}���T�q*Y>����?�9�'hVJ�� �l{񜉢�\�C��^D��t ���ݩIW���$��2u�#V�HPo��0sxt����G�>�XV��c���;���l��.�49J�Mw����{3�Tl'���$�#51�X1�n�ǁM�y��1��o^����5;���bc4�k+Ph�r-�,�J3ɝo�v�� �&7���R��4m�B��&�m�T�Dߙi`��{����=�`!$.��O«-�i�|��B��څ�Ʌ;	�ɷ�Ѽq������U����n ��&��6�G�4�����`�ii�[	�T4��Q�K�ϯ��󖲌�>���ѽQG)�;\}�H S	��/�-KĿYQ�s]�[&zD�3�g�6%��Ǽ�_Ar��u�0�7��J�qg�����$`����>�)�����lU��ёW|e�IV`�n�U"gW�H&R��0�:����qلٮ�`�|�S�U��/'E�zmF�b�˰�{�Gm��|����G��� ҄(}�j��8O�7�j�˫9�a�YrS.+K�j"��W��+����b��f���(�F����?	3P��2g&?`6���_�ۢO�V����<ɻ��WK�?#���Rl�k=y5��ޗ(������\����U�%h;I�WAN8�G1jm���fI�fNl�'/�px6)!_.e߭O;w���{���U�_X#��k�n̈���9 -ާf������h㿝vc���xҳf��Q5��i���o  ^M��������l�ss�_vhP�Y�?y��k�G�7YU>��Q;^EO��70�{?�[��A���=v�LW����R{h2g�+X�P({��[�;�[�}���KЇ�!�H�`�V�R*'d����4��O�[R�b��
��4��4p�����'���kOX�M�^_���Y
T�;���@גO	�a��)���O�;����Z�;�߉q�e+k���49��̓�������V��X{9%׹����s���RIu���Q��K�Ʋw��|�:�FXn��W=	tU�;�d�9��z\������9����<q0bO���_�9�J�a@����kY�����#N��OFjs��p�7�$
�>�W��-̑w����-Rn��j�6&Z
��M0˭��؝^��iyt$y��l����e� �k�v%k�<=�i�3��&��0���`t��!���6*.��
9��� ��ޥu��Q��w�9e
�%�%M��m��wN#�󸖻2k�T��®��M&�>?�Gkˣ����6����,u�r�/�0ׇ��c�TH����2w��3����GY�W#���>���ƌp&�� �K�*���C}�([�wd��*�1����D��{|�_:MM�[������@�ȟ�Skbf���_�r{�bHlE���~|��.-}�%�Pi,�p��E�K�T��0����r4��b���n����Iu�p�WDP�|
���b�Q�i�p=49�J�,݁yT��
�v�.�g�}M�wj�A����u�]%p�>���u���Bf(�16�<@���9�`8�c�l��]�m�mln��=E�M�{�`���q]����H@Bf�+=��V��YcZo3x�R�[����I���3�Y�}���aۭ� 9so"��)��=!aө�Z�(kבiv��
��pCi��wH����'�ՄFt
r�Bu�{l��<R���c�&���-���J`��%-��FD��q���+e����u�Ő����+=y�������wD�fx��a�d]s����$���3������_-���ՇEnC���?'nA�5qjh�[��ʧBW�_ƠL#���h�ZfK{�m�[���Y�i|�i� Lޯ�>�u5�Z�����ӪT&�mqhH_�)���¿L} �T�t��>ծ	j�}
��Y�}kۓ�>�%Se��H�8R�����ћ�a����l��]1�9Z�إ��J]R��XJ�xD�8Y��}Qy�L��gݷ�L�p/=�kA]1��!�ܯ��b�Z�PG#�Xt��5�2k4�oy������A/1+Ў�׃�S3)�ڢ�)���=�A�������U��6棿9�V�i��2����#\K�o���8f���Ή��.RzT�[�+���G�Y���Xg�ȿ���$�k$�V��v�J�&�!�eH�)Z�7W�C�Cͧ՗&��-7��ꫴ���5 GE��.��$'���	`G��������-h+��Zձ��Q�~�L�!d=o�*��jg���^:H�Lr��R���I�~wc�ʌ0eY�[�K�f0jh��Pt��Հ�����ywf���U�qg����/��!C]PKO䴣�Q�c�u������Q�`0��v����
���@�� \��P��-� E�EԌ�VX?TƔ��-�9��9�[�����RZ��ꧠ*�O_O���!@U�)��Ky�Q����hDϼ�Jt7Ҏ�d��3-&7�Z+%_��:�L��;_P���Z����ں�l�,bΔmՇ	`k�5pc�#�n�+TE�*�[ z��&*��A��ß6t�b�d�_�߽���-��JF$���'Ѝ��v�ܛ�h�� ��ډ?�\JT�w�5��ߒ��y��˓*��	������Vh$��^MX~Z��b�V��s�0p��V�n�7��d=��f�]�C� i�)!;��k3�IӦ�3b/J�ceӑ��`m>3"�|�Lbib4��I]�@ġ9Xy�i��k)��c�Ry4�}�?ȓǩӡ�}Z�Ĭ���v�p:G�Q�	E��:��5�X�i��'z~�����3�>�c5�)�R_$��;ysD���hert�����1��y�蒟j~b��d���Cﺇ#G�1�j�
)��i�Z���s��b��u���� n�� �~*�	2{ý�x���5���Y4���i�� ��!g	�"�"8uZc�Ce�06s �#�K:}���7V��j��)�'��|fm&e�$��o�-�Ô!���J�\��T5�z�<#rsd���Ԇ^=Kl�x�h��]	���n��s^CЇq:��$*��l�� �k#��s0��L�Q����qY�0e�_�#�T�L�1}3�⭆_����I�5ɔ{�犬ҙ\�T�=>��4ق\�b�`v�&=����;����cM��F�s���3u^���:���T1��yAj|P���h�V������[:h���u�`73#ŧ��s� �
2s�qsT ���uRs�~0�~o���g7�,<��e��zX��N�oTLr��O�VQ��i<n�E����#��3ugk� ɱv=�o���v3x����ᦛ�mD{����a ��r�������%���]��gB�j�;~eP$��&��K��o{�q�)U����koU`��(��a�ß�пˊX��qN_a���nboqqd�{�#paZ0�bu���Bu.������{y���@YV���v�f�FY�s�#k�wp�/x��E���K!��	��9�ŝ�t�mk.��p 65�МdXת��	h�\����̪���E�E�Y��0�8V�Anz�K�ɗ���zY�ٱ�41��k��1�/ZPl����v��U��zw��X��t��]��-��S2>R��|5�>�놏��-�ZB��1ά�m�ʝJ�]�,E�vS�����B ����oH��OH�WF-!�r�V^��f�{�<���ŗ�^+`Ю��s�8�wد�*j��_�?��<�vQ9��F���N0��G��Cû�
[ȥE0n�s��� ��PZQ�}����p�q��l���y��}�	�ZP*�-��	(gи��X���M�Ʋ|�n{�flc��S����t��j�s.���)���{�16]PTad�2r+�q %,�2c�̐7
��2H^8�?��c�|kH0�.��-�h���.��VYgU3.��g�Y�.�vXwο���A8��dq���+��,�?����PO��ǔ�|&�F%W�!�L0�*����e�APk�I����!�]����-�03�z���+XvO�tk���3�KU�>ʉ�ʤp.�a��k_�� ���Qs�	�H����?�=Ҕ��'�04a�hBi�2�=B bs����TR�����-����Tu*0u�̯`��$���5���ǐ"�Ça0�o�.�KyG�cZ��QI�L�j5���a,����L�������-G'�ћ�k�Dö��뛼�K�}�%�Z�툫�̡GyMGo�+�U���@�
�'��I��69��Z�\������ r�2)���˿�J��TL��5�f�&�۬ IF.��3������,�!h����Q�k$i{H��Zݍu�O 3�V�4�#(��'�Q=2�f�tUK#�6b�8�k�HP�a��֓FE���q��~�_�o_���ⴱO���<���L�1/�p�<���@9�]��"�����Q<�P׎r)���p.ӽ�`i02��sI���ǊSa^��7.��ų�Cn;ڭ����ќ�
v��:��V������Hs�^�V]'	�UJ3�C�-K�xՙM�`a��M�2�鷥1C7�(&^�h��2��X��
S��e
�qm�4ztC�Ab�ՑF�_���VQC���:��֥Z�/O�z���w�H-�s���٧jD�Ͳ���l�}�<V�t���-܃1�l-��K;�XN�<��'�߭Ox�'��Z�I��O�, �δQ�Č_CV=��7���f�K���2=>�`�۴ؑ�����w�s^�hAt},>����B.X�lwKa��u$�F�?H�x0�㌋cx�9�]b��� �r�1��"B��̤��86R5Gu�I��c	;[�.�L�Ǽ�����
]�v-"{8-�U�j�I>d�m}n5-�\_�)z"�<��$X��0�}���#�9�m�h��&���D=j�/�5?�ƌ��Ie��ԓ���	���uo�վO����<Mr��ExG�[�0fMn���8��CO����i�p��t�O�r�Օ��F�\��έ��/��U��x�s�h�/~�X���@$ ��v{ʆ�*i�c�v!�W�=Aح�A�5�n#�]��@��~��6�[��6���~���dժ�+!U����0�b�t+�/�1O]��=%#��2Jg�P�:S�-�#�t�B���6� w����p�d}�a�IA�# �H��CT�)b�.=!r��޻�K��T�nm5����U7\ ��,+Kq�ހ-Tj}�e��<Qu��;T���'cg��
^��\HM��
�4�0ևV~w[/��C�$Ǌx׊�"��~����7�&tW���W7��6�Tz�s�E	bM
܅	���l�WV����f F�6~ӕ�����-� �(P2�B�����~���q
�k�RŬ+�:9�o<x#֊Aut	���Ө� ��b�I.e]�sp\#�1�$��7|��k3��)�<�i"��?仉+�z?�.�>�P��2��O�h���b᭹5&9�I}�y⠅���P��bca�i�QpZ������r)�Q�[DP�2��^��X�T�6n�/W� ����OJ{{~��n
S�Sƭtς	8aX������|��дi��T�.k�[���ĩq����zv� �>�Fe�ѽ|S~r�S�+�V��h(X$�9�]bT�W��_5QW�n*��|�.{Q_���jq��cG-���Jl\��,L�j��n�G���߇C<�E��z�Y�n03���-�yTn���|��l0�v�R�d�F�,*o���G.���8S���,������;�X��T���3f�V7�AB�3�L�&��<99���YN�e� Z1V��BBu�\�`�~��Z@���Ǹ�L��Q��IK!��b"�7�b��K
t�$���s�K�T���}��JRp�z�2c�6���8 h�2� J�l�3�*	h���ݟyx�jN%7D�#�OܸJ�+��g�s[��S7�俊��~�ٝ��1
��th)"�t�j^�1��^�Jz}�´�'`1�6�hm���M6~G~E��j��6;��KŻ���$;�m�l�(��Yg�;��?����i�"��C������v1�1�U��D�{��t'g�)�OƱ��^�ힼꝝgD���"�3Y��~��B�<�2�@A�^�|��% �����W��L�)�(�'�̭��4[�����0+��Ypԉb��W�@�/p�����L}~�'�*E2,n�t�n �sb��T�"���+�߷���SM¿����Q�X�ԭ�0`$��5���� ���5�v���5/�(�(M��\#�w�.�bRB%>��J�@~��w\�]�c��*ۆM���'.��fF�r��Z �U�g�_َA��/�S>���Q�W�`�t\�(G���/B��>;��G8��$��[��	�Uΐq������<�C���N`����Q/����9�R�ܰ؏��=x\N�j�a�w�]�B�]�gΎ��ٶ��# ;wz��@��\U��svM��i�~E����x��Q���*�ȉ;�[��x���1�0�U��Ui|/��Oy����g&�~�,M%Gk�ЇV�î�HGR&�7	EN�=k;��I��	:D��Y�g%��[*aZ�5��x��9p6�E�fC�����і��D�a@�ӡ�֢���á�rG���1���&)A?NS
�bR���n*��*���MVwm�B�������w���H$Q������@u�°LA���KZ�p��$�T���L�� ~�<�ʔD�������u�}%S1��n���|�-����-4�7v��1��־�)�y�~0ţD�j&B��S�F���Է	��2���.�,�OP��;H�<x�a
������H2�i_I���Z����f�|���qO�%���2w�}M��~M�ǧ3�܌�z(w��m�����l� ���"\$�&�銰�;��<�=�_�{Pb��YV�:m�~xY�T�4~�.(G��j��V.U³B\D�$qt�yI����� �\���𞲑,�la�d3��
s-���m�����>���i���G��� ^��G;�����G��`
��r�|ϦE�::��XU"�C�=������Q�sGs&7����Β#�#S<��IMr_�#�<BZᒆ���J�����֋�����Ɣa�[�29Đ�DW/K{}KC����w�e�ې8��\�Ɵ�Ȗ\��=M��d�
�r�f:MLf���Ϝ��u4/ԋ��͡9����.;΃V�&0KFc�~�a�N�5���n��AIv�B>�h��R+Yy�]k�XE'X�CG!�JǼ�}�n��xۏ��]���U�����G�*�%�AU�.r/�;UܔF��P��a��O���"c�+���-[��N������=0�K꼑�
A��6l�kYL��аU��_sh�h��t��I�R��	3�8��w�-:h˳tA<�&|�Cd��=z��zE�Ro�JV`�E��}B�1*n�	]-.���x�B��>N�ڢ�<���=����.�b ��.�h�7;cI�G��}�X?'op����PsjC�C���		+��y.�'���Ù���|����'���7�%]����Hk�`��'Md�n�D��6,��+,.߳+�:��q�bhNw�b J�(#-���艐��8���hE���TD��f�!�s`.KuW:~�n�!x�!t��iV��Y��W�g�AK�nmh$�B&ʺ�w���Zh}�Qb7���Tw�l,�@F������K<���f0iO��֐YF�-"�9�쥐&�����!ʬ���X�H`�V��U�n!){�'��	����z�ngv�cm���h�}���ȘSQȐu��g�#�0X�s�?O��"�|�ɷ��A7r�"VE���G�Dhh
��B0��_�@��D���WI��*�=�[I���ҷ�F~G������g*�þSj܂Z�?����ߗ���L��F�ę�T~;���z("����-�_3Q�����Tx��u������?�;,H?� #?���*��*P���Ӥ�[Z���Q�C�y{#�L7UP(\2�m�aԃ-¹\B+�:T�N����T:v8��+��+�N�dY!t���Aj��?��2��P�E���+��d֤�O;�1Ԧ��V��oGp�d����X��}����d�H[��j�I K�r&sUQ)��D���u<ss����w/QT�L�N���֞�ځ�C�a�_�a��p\֙�� ��� ��#(L�Ń�\an�׸��%�H�A����:��>�w�$k�Hf��_�z�D��|�~]� �[��⦏��nY0������Q��0f��i����Hs��&�6���4�>�/Z	�2M��V���A=�X�Z�e*�*W�<��?}Q ���\JK^���` C����9D�f)[E3����������QG�x|�
���Ƹ$�d�h�@��R���c���V ���kT���aj2�
��5�]i�r캠��E;m��=�AB�qVa�/�~��?�G���]B����?�eՍ.����� \�;�o2N��3�M��Ã�с�A0|$J3V�1[(ƯB�
p��R+� o<&)<ɇz
n������o=ws�Á���� ���7���nD3d8��7=�~���a�0=�8��R���:;�|zm���`����9�a���Z㤜
4In�� �8`9��C̨@��0��h.��r%v��R�W���9j��=�oUm���h���� lL��TׂK�ߒ��\�C`����'��]m�w��YY95��E��&m��8���`a}\wO5���ZQGz�\���\�G�˕��l1c�����H\
��� ��0���ƽU]+��������4m�Q�g��T�?�2�F}*L�hӂ����k�p�>��UҰ��DQ���C����U����q���wb	>*�(��B> �'�+��lߌ��lZ3=���|�����H�,-���_�E�Ò��+eHb��O���;�qJ��àW�d��= ���wB�a�aW�6�ZU�/z��C�M~c�`�ld�n�lIk���,v�H
3�j�(X�B���0�43/5�:M�(v�����b��~<	��zG�����Kγ�90(��.xaF:�f7�Y�j��2te;չ�r���u��,w�u�r�rA�i�&B�Ԝ��ѴI���<���b���"�h��	��Qy&�@e� ���_��'o���vq~�z_
�������տ|T��̘��iāae;�X��n�rP��U���y�A	�5Zh���}ei��L!e݈D���+N���}��m�H�@��H�:H?�`�r^��X ?{��6�N�LV�{k��M0���erbYprC��Q1���Y[�r��Sg�dߪ�Z1'n�rh��H`6���^`f��;4��F��9��v����f��CS���m������VIg}��=�mAħ�ĭ�O��@V�$�m+<!j#�4,��䛏�dx���N��oby�����STː�����E��o��������c��1ҟ�����6����4S��T6�$o1��_�⺳�����Ȓ�`i�GI@�;�yu�rT�/��00N1u�[ICuO�s˝�6�;��QQ��3Nƴ���	���8溉��Y� ʬ��E�u/Eo����QF�"2܀$�db�ݷNME*\+�}ܥ�m�M��*�Ei� ���~��ϔ�Q�|�V����U͸a%�*���N.eڲ�n8���ە}�=�J��B.��h�0�L"��x �/�r�ۯy��?B'��x�;3��j�N&�&n�(�Z:xX7���*���c6F��[�c�~G��EoBz���V�����^{��,X]/V�����X��pb}	�9���oQ;@N�x��!ќ+wq_����W���NTF�{YW2�I�4O" y�Xy�+8Ri����%�Ð���u~m��B���n`חz���N�'$k�/��<)���Of��O�ˈ*z]�8�� x���_e(�K_�1	M��zc������2���59^M�[�<��d�����+��eLG14����: ݔ��	��h�����x��7�o����n$Ia����-�?������!�Qjbg��b��x�!�t���릢����p]�M�TS��>W�`|���e#�ȭ��;�Ȍ�-��(Yo��%���n����<�P��zQ�u��	�S��e��,|�ř��SXo)J|�0�.(�
��@I�A������Թ�/>u�ÿ������#��OIc1�]{�Ͱ�{��"���~fR]gs�
RU���
fӺ1���2}�U�$َ���>�f����`�ye��Td�oR��'~���N��3�lWE[RD�3������{1�i�9��Ե<��cd\)}���Ռ��%��n�߿�������mp��ӂ%��'K��E�Ȓ�ڤL&x;�B�����|V�XbW�%�:�&�ZF�q�W�+�~`Bڠ>MP��1mM`��8����pT�G�$~�Z��谦����&q]�}�r۳�W���D�8���%Rn��4��>D�m��9NŔɴ�9�2̙a4�<$e���1)m=B��7I< gS�G��fg�}ޕT��M������xgn���_H��}�@��y1S�΃�=�7m���K�6o����.ഺ���R��Eh�#���n^@tmH������v���Ms\���*�c�{$�
=��꥘�t�s���.#�延����Q�鈞D�N��0M,5+B��~�H�=�&���*e����ޑ��/�/܇�������w����q%#t��e�I�{����>Y���B5��w�u�W�j�kbt�џ;kX�Kdv��ZT�*ޏ���"�S��%��3�v���$O2oL\$M6�<����-�,Us(��D�]:4Z"�i�C�3���v0l��-=��쥼4�&+�y���J��t�^�k3�-0}�:X�d�E,�U��Z���zU���d��J���ն��.VM��x�9�ceV;����y5�8�5{6'l���r���%~�����\�b���� ��j�����'1я��r��Fr�4щ�pj�gX20�$�l��>�T�{T����{�mh�v-F�qT����dM���pnB6��T�!-�GC�dǓbs�=�j<hڿ��]�Ժ2~�݋�9-�V����}��/��*oo0FY�|��*�ޑ`������ၦԩ��4���E0q<�����+G�YS�
#�(z��g'B�!�4�@\Yf0*[8QBzKMx�I9��*��.�ߦٲ�fO��Q�B9[Sk�����~m�J�$vea��)s��M�V::�O�l�����n�=)
�<z�#'
x&~��� �:���c6{)�-��ݙ���dLͤu2v��x���̢Y�O� �)���F�oִ������7����ϵ9ֺ��f-+Ң��h�_|���z�������<�P�khm�1�n����e���\�q��S�b�0�0�!l���l�j�z�$?9��,s-���=yC���O�S������w��H
W�-��m�7�m��2�݋H�`�/�;�O�S~�۟Dĉ�Az�����f��ͺ����+�i�ӽ�D~b=ަ�0w͔=�����%[t�p|w��`���>�%��
�a���d�$[���yn�Y�6�	������\T�D瑮�=�mxN� ^�MY�7S����ی�[,�A�k,.�U'b�^�S���(��@j��o��jf㑹���ئ<����U�*rD.�7���L����<@���[<T8�5�F
������)�����>_�2���O=���MA��^m5�	�݋;��=�rd�w*Fr�VT�I�dxp"�Q��Ԕ^!?+�/�ߢY�H1�o_PwԠ{�#2 @B��$�E���_MZ�N��&t��iV�|�w����3�0;��� W5���mi]�~��x�
��ՠ�x�ҧ(T�!ܱ~���=%a!�v���np!W�J�Б�X+�b��������.��H!=�òA�}��JGIrn���2������p2O�����_aĭ��ϲ �$�I�9��M��x�����Kɣ�wQ��G�jV�$��P2��b�l
f��]#�G:����rKTcΛ�g��yՕ�E�Є�9�G�n�"e|�J\#,�2zqn<
��]�>� �<y�(�<,b��ސms9�y��^��{��y�O;'���o��v�{�"��T�0�8�n�jIj�Ңƙ���!I��5�GC���b(�%[���X#4��[XL2�^�q��+bo�� D�<xr\��X �{
dvŢe��.�A6�WS]�b�#�0c��h��D ��0�}s>��@o]&Љ�/�����A�Hƈ�ҏV�/��.�V�rQ����]8�Ƴ�ۂ�!��ؑ��q�"�>�"����3^|���;^%q���@LW{L��FzZB���Gf.�#�SVo
���@ �� ��N�C��$8��k;� d�X�"֝旇�:Ml\��>�vxO��dX3�B-���p�}4�0����'��.�z�F x��c�Խ-t 8��h��nBB,:�PJ��0�����) 	����xa�O ����G������*�0�y3�h1�|���L7���B��~�W� 5���P�8Q����>q����������~�q ʹ������q�"�T"�N�'S!���Ѐ��9�-?��n���Rg�X�	��T{�(��I� $�i���G5ψ�?��V�
��~�><DY|#-l���#:���m�:1�o���v���HQ��sz�~�|(W��6i�åJ���	QM��띄\���?a��"�H�1���*��M��0��Rc��ʀr8�/8m�YY��ȟö&�o��kk�H���������f7�$�&����3�WZ'+��L�QWF�b/�[��1�«�_��������s�~qmR*��V*��h��;��x資��x�)�<kx��V[׀�K����Q���,,��ie�Tg�ʼ�-<0�Fٖ�3�u��>";=���!��cL�XPl�} '!�BZ���Eڣl���b��,j�����b2b2|�jV�`<�1�&v6z���O���3���P|d0�O�%ݔ��u���њ��q=�Y��D��яfc�jrRH��n�Kn��+��B�6'�P��@K=ɢ?N��������ͅ �N9h�3���4�*�8|/?`VTB�}8�~�\}��ﺚy�		��A�x���@�ͬ�4��@�ф�Ry1?"u��~�|����˃�[�G�4���	�M"���xn����7����/A_%��Zvȶ�'��]���ꁫ�*V����W]7�(���P���D�Ž����љ��؊���!{�!���2}ۗG�Ư��@ᾃ�Y�t�*K�<�h�ò<�~�1E뎯��T�P0�N�)1~D��K1�Є�KG����6"�"���>�M4}G@p#"���x�&���+��BƄF�����22G'��⋘�c��P���� {��u���^�g�KJ��~�YY�P0 �&B����m&|�h�w������CFD�D�����w��-t�({9���C�J���;�ư�|�=�4�ă!����ۧ]��F�듖P8��l���cS�(������K���d�v�z�.�M�*����ܧ���*#���s���*��w�-lJ�5��= ������)�Sg[�<�i����AV����(ɘ���8A�3m��zE���ֲu�z���u��P��do.@%j�B�5n�-s��YD{f�W�/H%
޽�o���`�9C�?�	B�M�K���p,ߣjD�إA7�QW4���
>�����&��҇�Q��ܯB��,�,��Dm?��*�>�HJ�#��i��NɯmB�Eh�R���R�{]"Dو����k()AX	-�&3Mu������c=��RG}�`���0�Ѩ�v
dC#��7�%��YI|�
D���XI.a-Ǚ����Gu�:��H~�;��N��"�+ȴ ���W�fm�c2�5����
�roO0hD;˺����>��{�v��ʪ(�n"u�`A.��e�٪���!�8y�H�@I��'V9��� m�;Nc��I���8��f.'dg�а�5�f�π����FVsm=]6�>�t��]3 ��� �6�|:����ätq�4H>���dk9|��Al:6i������A�ّL��xO̯;wP�	9ʶd�r�#�-�=��"8�4���� �ʠx	�B�0k�����$-x�D��6�ؼf06�|1��E���}�����Y3�Z�E��օm+
�G���3���)Z��� \Y�3 ۀ�o=,�M����$�SK�3����M(ڸ�1�G4��w��kp�{WrA��B�
�y� �|gW��)��Cj/A�x8�a?� �lr�{��瓡o�jh&����i�I!h'{���б��UA^��!z*��'��}�E���� ��l�l'��r�����D9`))e#��g%Ab5��N������	���\m����~�wْ���}�cn+����>6����*Aa˓�KM�{B|�/fԌ�>�x9!\�6Pw�܅ Y�~R���cO��,�ⴅ�y���:��G���]��k�%�JӪ�������ҁԢ�75*us��t~�y�'��g�l#.�Y��Z��Z�)��l�Zs��*aV
��WÞ���J��2�H	������5���z�Ρ	����'�d� )��`&E\Fk��L'	Шے���_�@�*ʅ�@���@Ȑ��������.��oO{������)`��C����j0:,Ԕ����Ec�����ۢ�
d�'���H���Z��Ŕ(��Hcͬ#Ԋ�C��*
ч�p�o>�%�-��/�?��|�/�������]�4%�]K�L <	�*#���e�����X*�9�];��=�q~��B4q�W�K�Hʞ��/��hY�Q,��p6Yߊ�������"J!}��#t����!�E6�Q>���$�i��.H?5�d���&��j4"~[�`=��n�Y����~!.ڠuͭ�bݻ�G��$�&�Pmd@��%���(�|g�SU�d����8�"�.�PyaiB��6�kZ��)]z�����U������_��E�y�"]���9h;��� q@��U�>*�8�e�3���K�R��Ov��Ж���l'�������>�#T�6��d�h�9=���6m�rR���d�>H�ĤFMrY���Q*|ꊱ�U8�{蒑�G+�A�I�ܑnS!P0�8^(�Wk�;_���YHU���~���0��:¦�^�SN��w8Tx��[��ӎj�O����x�h�T�=�2h�W�@Y+&��
������frRi�n��9�����O��"�d��E����O]%99���WTR2{�4�r�[o��8��#�S܏P��:Ľt{l-��D�'o��ni����=Ɔ���A�l��٬��:��N����2&W�������I3/��I�rvXf]������Y�����7�F�v�B�3z�MGp"O]�hQ�a y3���"YK�0���qCV���ZK�>� ����" ��D'U܅W߳�kp�JQE
�V���A�WH RQe�- �{E4$+��iPc[�2еTk�z��IO
B�"����$��
'��,x�Xj��YDZW�r~�������A�T<,J�`�� �%��o��?�o��(*�&m�X]>�В�fL��5#Xʡ� 1Fw�TOUv��� A�6`3��]O&F�Gc����o����Qk����L]8���p�����d"��9�)�D�l59�ZI�p=��Ȱ��g1�w����'�#�b��^�#{�71�B��ZeȄ�
��ްE������>s��t�����U	C�ّ��߹߇�n�C���Bu+E���Os�H���m="��%³ֲm��U��n[� ������*䉮�J�G-�>۟��A<��[���(��H��/��m�B�z���w����W'}�tC�5��+El�gՑU��G�@d�?rH./ב�~ƛL�����"���{to �{y��={���`(\�m��8��z�v���7��?a����̾�E��?cp�u"H��I�R�䙎�[�A@V�W�p�n0%N[��)&�U�Q�y�t�U;	p_?�=V/�:v�u�5��
'�1��52���*����ne2�92��7$��OT�H5m�ij<���v�n�>�i�
��J93�����M���KPã82�h������� �¤'�g��qxV0��n�U���^���?���^��aҚ� ��T��ff�6x��+:���,!���h׾Q"�5�)�pJ
G�]\B��MO-���wQDL��[��!Cr��
/*�$A3���y\�"*�*"!�hC��Y��l�v0�����Cu���^y�>����{^>��)F]N�V�Ѭl�b� �	H�zB�J�hZ#M���,�'𹮁���A�R��1;)�f4;�S�I%Y8�}�o�c�>C�� ��~2�9�bةS�^���kf*s��F>�*J�?�Oش�/�����}Z�@�d�߳�śS������u���s���n�+���(��1+�b���x�UW�s����:�1%2N���D%����B�)v����d��8^�&QDD�)7G��r���h�K�BJ�"/S��L���b�&H���K�t�nm�_��	}޲��Ֆ��n�SHr�Z
3����F�c��B�H /�`w�u�߃I)�|̲���p���t��1�E�*)���K̡��Ͼ�s�4�=ِ��������<
������Պ��*i�+��Oe�y�g��}�\���%�����0��X�3�
�3({ȱV�7�	���l�o7�&I�(kL����`%{Q�9[z/�eKZoE��ԍ������X�jyN��n9�Z��-�)�|F��K{5��q,����6����n�[5��z��N���E�+GZ(�����1���v�0�?R��K��|��SErGҊ��sdk�x������Hj�d�j�0��В +j�ƀH`ڱ�ӪR&Zy�n�G�Y4  S�ģ��S����sH�X�Ԇ/w�j��6�ODٸ2.�O;I��L�~l��X２af�C��:A��c�1��9�N�āj0�	Š>���^q�LQQ3Sy�5��$��o*��N�s�:}a���ܺ��<C�����:��;�+���T_��W�w����_���ܵm�#F_m"@v����_ΌiI���l2a��N��Z�F��_�k��ꨟ��3�`Ů��]��A�K�h�E�,�و��F7βȵ����9^/1ɞK�~�K}���)Oͭ+���|wx��f�f�~�᪱�hB}��,l.,)���V�e}(h�@b���xY�f���ư�%=�9w\_I����"c%���)gLK��s{��È�X�W}����v;����-��lB7~ie�uC|��ռ�J۷31E��!9�Oz6���ˑ�&J���+����@��Z՛}�L7�4o�,�{Dn;��M�����@v�e��c(Y%2���Vk��m+'�Q��FMJͧ��/Ӛv�\Pad0W��)=�!��DH��v��$L�`���"�T��QUP�a��f��~�-pU�B(E��+"=S�|�5$�9���q�/�#�_S�h�ٰ70�������P.,�S�1f&,h�&,оFG�=�rB�E+5�0���F�,�R����{�Z:�:9fu�{��Q��녨�C#��@�� ��K�pI�> YMH�0��:�$���3������=� c�t\�?�^h�N�E*���)A���m��K�G~fJ�W=|^���DO�:ِ|[߁��]��-rQ4.~_��H�����=�ōHM}؋���x[w[|{�h׺��ʕ�Dؼ'
��o4�ѵ�����t���`p �#+̎��ͼ������s�0`�w��]^iKҍЭRQ�e�J�� $5s�V�ޣFN�%ϩ���]LoY�#:J��Ey��b-(�E�Gw��f��^�;��~[D�]=�d���Wn�<(%D���/d�Z��6h�8�r��.A�mt��/QD��,GEށ�%�� u�r�@�M����X���\�R�l�0''��;���c+A�'�<&����ګf!Z�9Ȕ)�#4�u�-$L�ɢܺ�Fw}6P6��k����p�x|D�NlnM.�+�'b�bTLp�F���J{*q��')o�KO�mc	��!�\�-]M���U0a2Wd:�ThTY���ŊCb歪8n��*d���br���L����^�Th��[�x�bZ�~Al��V�<�\ ��D�]K^�	y�Μ�BΈ�1���I��MR@!Y���6�m��c��_af3�f��H<����{ �����w��ys@̀Z,!��M�b��%Y3�U��g�	*R
��P>��b�~ uNH��M ~p����������x��·���t�����-�#�XFO��$�\!j@1���B!��s[�i��U�`��1�u������f{��{k6�O���	0��C���G�%?��Q�SjR6���1��KG���L-�p�"�s)�`Q$��Q�ٹ�q�M�Z�Ka�+%�+6i(M�3I����V�,�ԉI�I���KD�?��'A;f�����������ք����b�ų�����(o�ڻJ$���Hq���	��-H&)�����!�R���:�T��R�ϴ��y���)"�E����J�
��z_�=���Y��8l�t[z����P^v���D�<O;�r�^3�! V�R5��*:�k�Vʬ�k��c(K�*�o�U�EQ�B�C��(�1O��0w��?$�KY-�H�;��v�ʈ�0��?cf�[�(�a�p���!Y����;/�q�v �m����r.'gC�Np�M� {�@=^ 8��th1���p^;��n[�U��!��cu���~��&~�?@�ˡK��l����Ec�a_�Z��KD%P����;3���-پ)��/�%TR$���{@/˰;рě23g�/��񰧊j΋\~��r(ݍNIG�	�����u~ʪS��i�/�I��(d�.�)ǰ�^0oG�V���dD��hІ~~_�?���D�����P�N����]��*N�u�q=��(�{��͂���l�eg"k�y���� �[k����x`mK��4�n�y�F𪹆���j�]���n$�7�e+��4Y�bQ�vk[�G+����-Rn(@��)*]�h��:OΆڭ�b3�!^L��.���raI���PHK�
�������Ӛ�z$�S�14�~�A�����_�~JjPy*� �w�]�Ouv��;搨!�I�g�|p�$�+���b֔Njn���C��H�4ַ���F/��b���)K�3Ǉ!髲����~%q�-��o�wY[|{���e0���i�ܖ�9Q�>w�3u��f�g�\y����8�3��`�#\n��8�����"CB7׍�}��w�p��g.Weu�A{'I��'����$0������ ��,��ߌ~���aPk6��w!R��#�1.���)�n]�j9mF�T�ek*���A�!��Kp��QA�J��IUx3��1�FW���v*��u��"��F�C/q��H���_c�Q,���{e����<� ֍���p���U������}j�RA�X�����|�'l�3��g����S���b��ymY�����I��N��uQ�{�Jj����y-��M�2��Í���K��NDG����]r��;j�Ձ�ˊ��z��U�m����
P����x���|�9cu��<��ϋ�%���d�}�q)�?Y���4�g�@'٦@��H��k*�����%\�+9G��;/�^i�:�/����g\�7�<g�N�+����md���ʢX�!���!/.�5��azZs�]`��'l�J���Em�e�Y���VB��U΄I����q�����_M�C��F���ͼ�I?�����դ��@G��[CL�x]���~��B�,��<E���Kc@y de����x����.xܢ�8@;/�ғeԟ=��0����Ytm��
�SUh���VV�:��[;�:G�ÖWEJ��JyئaZS @f��W.�Z�!pڪ�
-c� בC!�d�٠ll['���*W��;��-�Gl��(�p���3Zֲ�O� ��7@IjD�R^IQ �j�m7�; �`'�	�2oh��	�C㲖Lv����J �2g��sn����Y�Z�/���x�f����錹F֪�z�Ǿ&3���� �=ӒF3���[L2dӗ�v���ض��I�/��Ic��.'����d	\[+�J=l�{/��>?�PW8-��[�<O�."�D7�}3�R8������E�E�9*�Mx�4���{�)M�����$tT���9wiAq��M�`��$���vS�Dn����S.�(ξ�ecX���!�	'M�ǖ�Z����$n�9R�L`_����=��T�G����|/���6�F�8�8�)2��>zI��t��Y`&�X��j�C��e"��#&�kt�X�4���e3Rf�c���4�����Ͱ�W���<�w�U�����U����~m��D^@N��`���ѿL�	��Ѻ����P�y3����"�̮���m6eC� 8=B?M��B�E��3z3��q� ��p�b�cai�#k��75}���g�����K�
�fqZgZ�!0G\8mUh|`]ghG��h��&2��gf��)����6�,�N�P�
e���Mob�pp`C+�q�7��wQcة�'�ӽKN/T�5���An�:Ͳ�e���l�¸m��}I��%b�!õ[ƒ\�!�qBڮ�n\����ev9��hj�Hލ��+��P�<��]Y�%�F�_�(V���c�fȫ�c.�(��Z�����.?3|�x*G%O*8��d:;i�!~�8<c�;;��U&���GN�,�^(	��+�*�H�2���a�cV�M���d���Q|��GK�K;FػǸ��ny\.C�|�aQ�ڤ��5Q��ݪr}Y��I~���'-����3�3zb���D�t�s5�D#K�$���y׿�������՟��p������x��s��b4��#����u��M��]��eL�X�;���@q�Y��z�*"��܎LI`X�s�;��}��U�'`��{=�2~Ѷ/f�O�TF�E���u�
��ٟ�iȳyxn�f<JeX^��T��/P�6B��c��hJz+'4l�CZ�F�8�[r� �ʿp���HH�Iހsy�/x��*���"���7����.	a�2�U��75ç�b��ƍ��d'��g6k.\Z����IB�������l�0���2�)[�>��9qp��/L����t����͠�]ׄӱ3?�o�ˁll.�ۜ{���X��L;@��W��ߞs9E���,��Hku�]f��P�2<�	nY�������¤����P汌;�H+L3E���*��'��y[*O�k���d�qYǪ�Y����O�R����Ah�mC����ȼ�Y��\e�k��|_��ꥬ�Y�3h�Lȯ"q�GLZ�����=��۾Yu�����Q:ܻjF{jN/��q"K�4f/�=�!���6(���v�����8�S�{ojLb����8˗i).4�Cl`��R�ʙ�M�Oߩ
���E,�S��v�L8�/���f��4ͦlV���4A�t���t�~�]tN�ڛᒴ�{�.�ۈ�_�ac1H�	"�Zi��M�4�s�`�@ݸ���#h��4�H���J����(X��*�7	 �Z5e;�+��t�,�s1�[��ت
?��/ͅK��0�{r�ǳphU�V�	=�t7�U����?��Hp�,�<���pHH$�lك)��;�H���[{�'\ꪌ�W�4p�ַ��6��I%��������EWU%
)�W�}8�� F02�WC{(�v�?�D}`a7�Ձ@�^eO�r�IǨ5��(V״�m���j���Q.o���<Y�s-��M>`)����C�;}�0N!D��һ�_zP�"SQ��7a��!o�6�w���Y��dA�&Z(��C�
gpF�k�<Y�����;�*�F��vһ�ʼ?D��i_���
�RK� ��8 $��X9��J����ݍ�gmL �a:c����CG�p+E�T���Y��ۙL{ ��<e�T�N���lɟ&��g���RHz��	���v�5��p<:������`�fʆT�{�'\��ϫ�c���[:��'��˃ψ�QF5�q�g�s�l�k�^�C�-���;�$coD�gU�9�_��(y��n���ZZ�I��-� si���!���Xzq�G� �sm_�,g��R����7�sj�ۮB��?�W	�UE�,���ʤ^Q*W�t�$�O�� ��;ǿ�
�|8�/?Ĥ��-M;a/�b��є �}�0�Yȟ\h���AX 3�Ar1|s�}Y~R�a�;g�9�
Ҕ׹�K�������A�lm��W>�t��ڡ����Yʔ7^�r��6��U�qi���2d!1Ղ9f��|La��l����4!~��$Q�HYS?s�l��]R���S�y�+�6��-�4Q�YKK�mڭ��o�����ӟ�ۛ0$����T�l!��~��{7����0�>�*�2�5Ȼ5����r�d�	B��Bp�0���Ίf*{�#�*�z���#���&\P�T]��uŇ�pvo��x�ϐ�I��k��8<:���ƺx�M2޸=��/�6P�:���2�/
pO����bfI�=7O��;�{���;W��a��P8�)���ڲ-Cb+�@¿��%6��2 _����9���G��e�,�����B튒��Ч|�7ϩ�����V�[ ����{�W�?P1ue~�3�1֦� �:7ѿ������r�ۉ�5�w�6��Z�, x� ���X��;J��.�0k.T�v�9�aG��u�� �����˦+8,��~���͉�e�Nn����6եmck�1t�Y��t�6Q�M$��lA�P�������(��x�[��!␘����	���W��u���CX0���b��}Mˊb㵇�a�9�LT/���0G�����k��'R�Կ����T����[�V�NX6��r?�vD5jJ�b�����I(v�YH��p(��&
8{~pE�Q��4s��G�<�Wm�0mV(�b:aw��`&rKN2�����kk���ѦC=Hۄ��J�\�{Y��93s.�[�&�0Ϫx[Ps�Ƥ����WI�@`s��p4���g �ꈙ�`I޺~Se�����*����dDH8&CE� V𬴖��i�k]�&"��E?ZU�k=L�zf����ʋ1d��!���^�}Ԥ&�
���{�NJ���)F�ͮ &�2b<���2�����,��I*O畷�͆�T4� ��@+�%���FxP4]f1�����)�KD8_^o?���������9l(�O���W��l�/Ո�}w�ځѻx�w�q©��#����t���G<`���C0��$�%��o����ЯG�O=y\�B�s%]&���}���aRk���@���(|�-)y��nOs_j_�B	�8$�v�/�H��17P�ωН��g�Eӌ�"�D[r�[Քpx"�F���#�מ�|V:$:b���M�\�2����0
a����Ԗ��;�E�+��[T�	�g���\	�v�,jUZ;�g�Y�6���w0l����fqw��R5�x�"�~�^�k�#i�/���J

�[ȑ�h�%�C�m�ɅL<�r�pY+<�8��$��;z� �B�d2�&�':[Q�9I$G�!������^��;\Ҕ&G�W蔛����L+#��u�
1�n램z�j����ݪ�.k^�T?���׆�gy�X��7���cF���jN����쇨�Bv��	�r�߾��D-�N�R��Y��:�.� 'غ��>�`U!|z�%����;,qE�[*l�s�F��~��D�T�c�/མ��)�r��c��;��n�!�LE�z��l�# �}�(M��$�&쯌�;!�<�M9V��Fˣ��,Qwk��ݰMTng�glӨ�&̽��.�
UΙ]6�3_w�[���_鷸�\;Zu`�Z>�f�+�[��$��>�:�����l������򫤊h�d���F���L��
�Vg���y����ot��g���3��+�B�;+�+T��Jd�OGOd�AsP�)���C��9��P��#�d?�M�я��e��V�_��-/�@��6�-�ā�I���C����/�S(���A=�h,��(39@k�����8&2twCɣ�����X�T���ݤe�fh�O1,HJ�獰�q?+�
�JO�F_Z�&�1+@��:�P����w��k�"��ϯ@[Y�҇z"e乻9E6���b��&��$���K��G�"υ�@]4!�d���mU2���ύu�)��0_L�����e�{n@i�3���5���#�)�QUWv�1&ET{�P]H�	�fX��{��3j��ї�\���=;��V��7��t��ȳ���^LQ	�NZ�@o�VǞv�՗�x�3�	_=�C;Zr2�q��5.>sg*:s��;�%3׀d��)h�Siȹe�%/.��7Ї�@%q�t��?��:����!7PH~�r�i*I*�Ź��*B�a��3\FV�a{g���T�ӝ��U�kk��T��|Yl�G�Yt���g8��b�I@�Ry�]�a��Aڤ>4*��5g�£��­s�E@���/�/�˘����N��Es���g�A�
��N$��z6���տ�H<z��`i_�c����>L�RN��ᔮ�W��T��c�i���vEo}@�7k�r�$�Ư�����$���c�RKƲ{^#�	z4sWx��2�S0y�yU=4�����,� �Ǭ�;���6�hme003�u
��h.e|;�i��#�ʙ��hP\�yn�ʻ� 1+�K	}�E)6�>v��Me����\��YWK�.�刄2Hc+]���-����J��R����	o���Li�Y���-����X)t�v��,(ȬQ��i9և/d��������;*%��+
���ZR�
H�����g	7L��A��*�DF��g -rե�&_`�CA5;�]0�C5}U�p-~$�|P�Y�A��؍2�^��R���:�w�jiw���MxL���N����Bj���C������%�^ٞ��e}�i80k�m�������g0�pƽ���1Em?�$��4�C����H�!Y�)�WZ�;	AZ������K���Uc9�O	�o#�(G�(�/���/\3cK�.�DM�<���/x�a R[�mհ�{�a�cRF�E���]^#�)���;w��U:�ٷ��¢!�EۉU����b�~x-B���{g�ÿO��bz����7�/���������ZSط�
���A�X����ʗ�8(��Z�r�.�(ݗb����M�޽M�D�S	q����%v����uqj���}���a�	�ۥ��W�%��� �V�v#��+��_Pa�����&��4�2�Q�n���O�lֽ��R�*���W����42��,hG)��)O����鄢.,ҳ5�;'Oe��ۊ�Ë�0��=A�Q�tt'�5y�H�-@����;�u�h�}��1�����<;6
�{�T86}.���A|���I�OB����Xi�>T#��a�֝Yg4n^�Rٸī$6��Iu
�ԇ�u�RD���.�9)(KY�0K�\��
�A�)s������Y�*]����=����ӄ}8��!{u�w������8l�z�����hNf�T2���|2����Ս��H��p��C.�"� M)�n�*��u�n���͉��Q1g��M�3����Q��2������H�8�Ir��\ν��q���2�&�UUqv�����!�^E�(�<�z{��=�i�Zn2�b|r��a�=�29��`J.
�(�T��rW ZilP�%�R�i2o���v����ӊ_k=�57%*41��G�+�籑D����}t�4�%=Ip�:� �rJ�y�1���p��>-���۰4��*���	>:�t���/�%�������pB۰h��u�ed�i蛒'�X���+��B� ,N�@g933�A7��z�>�� �8�ډ�@���"xt���8nX'�y�K���/�l�8��ȃo�T�l��X�L*����w��5�^���'���̓HW�lo��8�ͽy��C��'eo}�	��AY���y	��N;��5f��<���t�5ց�%�\���>����u�����gS3?��V\�
����#�T����L��̍!o��Krc�,k�f�SN:���Tw�`����K����Is�6]))�����\����ʔ�������>s�fq~G�E%>љSIQ����G�Ŵ�~㛐;*�o��G�.�1�/����y�6��eV�PYJ�A���qjO_A�4/���ksh��c����j�Y�Wm��������E^��]����=�m���(���A/>�f|߄�OM�_&y�r��,rJi�j��e��_c���<�9��z#HA4$��>�v���xS�.�w$�Ub�1��[����M��d�42����
�Ԑ�_pm.��
��Ec@S_��#S�|��dS@z��h���?�x_�=�H7�X�̰����Yw���<v�o�K/by��Y�=�?�1͡5�:?r�x&�X�@TD�;��e�s�iQ:!k����eA`�c��Ǆϝoծ�����Ji��a턶T��6�p5W�G�p��IHȩ��������7mBq���c*��$�uL�z`�����@�P����S+?�Sּo�@�|�=G�:�%s�͗�����b��/ ��a�E/#�Id�nz�aW��Q�����ׁFM��i��2��G؋����_�;^�@�hк
A��,����[Ӝ8}3b��I�*p�0���.��y=�)�P����o�qH��8^XY�"\~M�^�����"����u5�_���C�F�Ip��סrTZOI�2�~��>�â�ߠi2�AsY�����Í,ߧȆ�E�2��T&�ʖ/�7�n�%���ۏ���,�C�ڗ=�d�갍	m�� ~�=|�\E�hG0���iHxˢ^`]�3ۥ��|)��s�'��B烓��3)93�=0�ޣet�޿x��gc���:AY:���9����U- �ùF%�X�,5~N��A��n�4�w0�ޗ��WId|S,T90x�.��W�itl�����`����b�)GL,y��;����=w�M�'8�z���l6$�AY�V��TzīX	�H�4�;�#r��;����Z��:0(�@M\���N�k���,;^�����㖏M\�ȉ�D�R����
�)5H��]��ư�h��N]�,^�t�d�ʔF@�<D�ݛ�;n@�H������m{�qmf�&y{�b�jQAJ��,�x v��1cx�Ƹ?I\Z��/Y���oR��[܌s�`��A���HG>�\��o7.������Vm*��0�|z���H�:G�4!����x�����֢�K,�3����!B����[���y�Gzy.�Ş�]�}���{��À�}��Á¹�4Uӫ6D�	vlf��~e��f��h��&M˝�-H��J�U1,xI�m�rQ5#� 2���h����=R�m��
&"7~XC�3��<��Ӯ9	0u<j��;9# �u��@&�7<g>�P	4���Υ�b�!Wz}���<m)�M���8*<`'KP��s�ޖd|��ѷ.¹�qj����Q� �Ʋ.y�($��8jܨڟ��ey���M�ږ[��RTq���p&)nm�O[æ��٭��x3q�7���������zs�SƏ�;�������g�����J+bQ�K�֓\��q�kL��M}$�� �B���Q��= ��j�c1}H�
���z�{Ȕi�o9˖ݿ���Ѐ��7��u99�}�j�����6�2(��0���;@5��f�_Ö���]�e\�8;�9B��:J;y����������
��HK�_�Z
��u�r�Au������kMO=�����O�Z�q�ەE��Mz3[� �|Y�*�ؐ�F�ҿ[b�������:p�o�i���Jn{����U�ޜ����qXcS�.��>h��-��ve@�B����7Ѕ`U1E���('%B�Z�WE�x$��:�9����6��ޛęv��_��B;�嵀P��f<Q�U�K���#y!�iIfGZ�1ށCѠj|�����,��ʫ�����, ��
[�5�x�o����ʋ���&�7�p��-�I�+zX^T��kC��n�s�I*�o��[�e�s�T�u"I��0n��"���.�B�Oo�RF�9��/��u8�첖7�x��>
AG-��K��nJ�U�qTk���m���$��C
�j��k��O���Ӎ�����?A?����-|���7�g퍭8��N�n^\�nQcN���t(���������7h�����8�9xR2W�Я�Y��fH�ݭ)��lY�s"�����X�'��69��1D���g�%X��W�U&��m��;P��L,������3P�^s���9��ǖ7�A
q�����dO&o�M�b`����F�}z��h_�"�s��9���	��/�������b����Q�w���#�����h���/AG�2�#�'�c�Ə�j���P���ގ3��,-Y��~�o�	�z���2|Y�7�+�nD$MTŷ�q�YC��T��7]�"R*q�%0�!�B�E��o�.ڐL{��tK2�� I�S��p`�d\��+�k1r���{m��l$�*��v��ei�&�Ǭ�'�$g1��(��lzX�(A�"U�e�H�s��:�8 #ė���7�����^ˏ�jn4�v,�C�@ڟe�Kh��M�-�9p��,�C!N�?�r����+�Ug��n�P�i��]~�%\l~N��ԣ�Ռ~�����:k���ۣǗ�V�g5��7q�h;+�yA��nec4T�^p<:5@��W���)��/�Gr"�1�f�r���KNeo�@@�;,�i�T|`�?�؊�`[�$�6+&�J#L5DlDA�?�Y�f'�r��R H��
���f����j�8��	�]�;0��ʌ3�	qd�1eBS�9��T_����_zV�(�%g%�����0^f5Z^w�R���i�~0��&���`�jČ�ޠ����T[����.ֆ���~��zi�X�K��ɓ'`���J��ݏ-̥E�*c�Ii`��O$���aTf~g��:�_�e�q�[D���:Df�Y�
�$�O���&y$�z�3LS���gB,C)��R�Kb�Os�Ma<"z1��Q���r��)B����`8���ތ�ڬ@ �������[�=<c��>���-����ne����aY�7�?�����\[�AE��<LV1g�^Ԫ|A��H��U�SԈ],�ɓ�FXP��`ϟ:j���V�2�՗��2Oن� ��;"����k��	TTߜE ]���ɭ����݅x��b���6t̯O[\͏���q��ک�F��˞�����	��ʜ������7?#c-X�����J�-d���>��7�R�ű��m]Ԏ�mX�Nǵ������Dt���X$�d���m�ɡ�h��YH�9�?�Y��f�\��ic��!�-���&�?�|$��<���to<G�we콒�SO�U���AN����`qn2uw[�ϝ�W�!�'��H0��eĚC)s�©�^� ��͍�ײ����@c��48m-�g�w�R��.: ��1�흾�tD�A^w�k���uN��K�v:Q6}���q#�M����d��(<޺���eF*�+����2�|=v�u����=�#$~�B(ͷ�?�ӫ�LT�v�_O�����O��ϲ;�H19]��OL��=x�;<�)��7�>�C�k�S��|Æ*ި�k�0>��3Mm^�S�Լl�A�O�������T�-���G*��)����D�^HNR!k����8�Ůr����f,M=v�*yf��{�4�R��R꾶�L� l����`.�A��ʣ�n�w�<�&�r
�(�IR�hF� CE܃��$���3E��)����^�3v�W��)�G��,E�1:��������a�?���!����9\�|���!���8s~��c @K���!����\* j���;3��QD�p'�qk��C~зi$:^Y���~6'<�}��\��zE\��=�׳�yPX�3���J �
��"*jz@1>��������@�������/�5Otv[}�٥�3'	����d9�ן�'��2�?6o[sfj��ӂV�l��߆�A��-�ZX1�u���7瞦�B���3�$��]���zY���vK���'G�3@����f)��B D� ���؂�p��h���1`�ߓ��TJ�d���	do�ιy����l�b筺�b��%c:�����a�!A#���#~�H$�[<r�I�=S+����?���{�:*U^�+�X<���;eb��3'��ba֜����ߏd�OLp1����S��I#c�{�6v{h$�r��cm��PFjRx8no7��Nn�`��u��?���Utؑl�ʹ���`��8
u���Ѿ����Ca��x�Y2�S'0�@M]�bX]X\n�\�o>�ж� F4�߸���8�(�i7G��?AQ��@�[�|b)�{�o��޴�a���r�}�L�OZ�.9:L/=�K�|	MA���H˽�H]I��u��g?��q���PT�] �՟����)��V���I�E�	�x�n/��x�c6`�n�:�_�^���$����cӼ�80O_ۘ����%����=���Kf����Y�@.����V��Z�EauQh�,������ùP��RI~3��g�;�J�[C^|~�nܘ��]����!����t���*4��C0�s��hBSq� �C?�7V��1C��9�:�W�U��A�J�[�mU#�ER ����<���Zm��W�}�>�	qM���SߒT`�Ӏ;�/�Y�JG%���&���j�1�z�ޙE�2�6�*{\�a	Z�o�űh#�����Ip������h�sS��񧧺Wk�U��9��V�F�c*�:�RJ���*U�ʤB�Y6;D�����3�d��:9$� ���#4��+j���n����R����G�Xtψ��b���'	v��|�"4BL��엣��aGQ�[�)�?��<�x��\1�����к�d\@���|[�����j�9���^N&AQ�!%lic_#�ݽ��
�fě+M1�e��o�~{O��[�qu=o\�bL����p��`]��M�>��1���C�g=�`J$��@ΩD�5>�KU��pLK����TѤt�}f�5Ż�\��;g����t3~����Ũ0�O1r��i\q��io*���N�G��d�Xڂk�'WY6��]�#�X�!NO���V�����F��g���2�~�-�������P$�Z�ʢ(g
.���1AUO�o��T
����C��}�)�ˤE(���+�G�@�0W�K�բ*N%Y�cOj �X&��,�H�.�S&���-"�w�:쇒3�zbsޮd����xi��gG#�������]ǅh��W~���I��&6����
9��C��\;;x�1B�m��jԏ>:gu7��C�9���X`�l��p� ��ńG�Dn�lπc`��+�h͖���
���3���	T��/���j8��b����Q��D ��SxPV��Ѿ�7������a�i�d��QݑjԘ�'��8nB���ڂ�{��l���E�dTU_����y)p�ڍ5��Az��C��ʎ��7&�辎f�,LaҔ�`?��p��Ls>C�j�T�{ 	��8�I�$}�!K������qC1�'�M��O/M~�;J���eWuH��|\3wS`.��T�m8�%9������}�1[������reA����ܲ6��C!a6'��`Z���'(��n6xKjN�z����	����;���rӝS�(�~���`'/�DNa�>放��e�4���;8�;i]��n0���M����y�&�q��T0��w��6C#�f_��&�-�y귺#���^��TG���J_	���w����9*<%���}`"�ǊYG�";7=�����#^j%}��DP�tXn��[w89�G�"� -�8{��j�v-��!@-���))f�L]�:R^���8gy�Vg0H8y�h�-�o�wɱZ\�:�����}�Wp�ƿ���n����]�v�*��٭K�8�ܫ�����'t�&1(f#fh�����������c���\��?X0���Kӏ��I�P�}�ҪGʃa�G���q�������C��!���/cG��Z�G2~��,w��s�__3MS�p|���"��t�����o�;�(�>!a�������D	��/���!�0�Ӡ��59��#�[�aA��0�^��+��{���Ȏ����)?/O�`a�`T�2Y(�N+!x�' �K�h+�_>�Z�-5p�����6��?�=�{�&$��g�3>�Z���@?4�晎[%�uz�=s�Yt�U�pI�7������2�=��l�W듡!�H`!���V?΅E��'Ϙ�2ޮ�{Q[�}��]�e�L��=��gR�5�i:��ή4�kW��j�)8n���ӡel��`��/��R��h�kĊp��6F��ٸ#�l�����{i�������< _�ٱ�:U�o�Q��Z'�K����
�&�_r��z�P�RD�4���g���Q���+� ���1C�6V�M�|o3�8ϷX@j�yI�t�]�eB0#��ƔeأIz��	c�Bd�Aa�ܓ$c�?>�a���������U�Wa�Q�P)m�x�bM����]n[#.׷��q�
�M�ܬ�ou�`���ՍDȍ��'����t�� CTT�;Y���1���EVw�#����+'��,u���J7JxӲ����ǒ�v�ʲ�zJ��:ǯ��w�Y��7��52[RD.�_"���-��F���f�'�N�JIR�;P=�@�����fYDh�f��L����6�aM�������羣���=4����Z���)"��fLy>^�)��J a��'u>z{��<���gZ���Ǘ��*#�`帱K[V��ԯ�JO=�����$���	y{ӞG��I���v"CC���߮Y\�$���{4C����f����*�ȨPM�M�z������K�S�����TV��3�o�~�cE�x+GI>��ߞ���~�G��Ge��ׯ��a{U��vŐɛ���J��4��G4x]��������M��=��S���墙^e�u��I����"&�e����@����v;����?;��2���|����:��	� r�%��*�������`�}R�;����hΉZ��d��t��s<ww�2�2�4D���R�6b�a&�Ro}�Q�4�����g��N� �=�i�	�-�l9'��ώ���C���#��BĴB���;���Ō�m dC�����3����E�cr���bF���A�8���~�*��0��."�A�E0��#�X*�Jv���ϲ�3��d�P�n��Y�k|eN^4ϢW\fuq'�u���L�cAYk��B�by�C�(Z\'�
p�7��]>.�f����|el��)�'�7Y�&!�h�S�c�)�Rfd���|\��Y��|1��-�_ڳ��6����UJ��r��|K�$��f,Ɓ����z��g�a�W�i�kq���@��������\��e�2N�@&J�yH��c�fe�z��?R���,8~�Ż��T~>�$W����6�6�����M<󋾻�-���d<�!^Ѳ���gw`�(!�2c��^4��mt+�)���}�"0�S�!�&�P ��V��I���s���匍�J��o�n�Y��*F�G��a'��a�*6�P(��6]�G�Bڭ���A��Mɾ��lPCb,�A֓x��l���g8r�����Q cc�(X�g�?7�c�e�s���k܃��hi�*>4�D����w�*�wc�;�.������q;���@Wa �k��� �'N��#׉	���y�S��U��x���sO.FJs�Wo���a�{ص�f�H�M�����w0����G\H\�������ԥ$�wbBE)u���'=$�@�2=�GR������&�$�j�z�yM�Y��9�<h)�U���l�����8ǀA���,"H�����$E@���9B\�p�\�5�Wt�O��{#��ݢ���5�����l���ը�<Ƭ���_��Ӎ}K�PV���yr�v"�w�^Q��	���>qn<X�4�OD�����r���[J�6����r�K��jH+M�ҡkA�y�C�`�~:K �w�{�ʐD�%���;��y+������������d���(�Er���m(�ol��쓳T�g�bȷel7q��YrU��*��=��Q�U����O/ܽ�\�rC�/ W`��^A��2SP��X�ڣ�/��*���Ybؾ�O�x-/�M�������#�h���x�7��
��R����X�,�\k�3��Iou/�-q�o&ۘ
#�������NFA҅�O�ѿp��Z�`��L��NY�Y0���t���b:������+�ʗR��=l��1�����K�������Z$�>՜�f�Sg��}�>�L��k���1L�5c��'yL�#=���jϣ��jd�E{G�\����p_N\��t���\F7е��Ӌ�a$]N2���I� 6G'���L$Efo���)Ӑ�n����|���52�-��������Bt����1m���7C���?�g!�#�kr���i +��w�dqEa��HOb� M��AsV�@�l��u|�mDۅ���U)����T��]ԅ�5L<��T�g�v	ʃ�<L��O5�^��nD�� C�a�Mp@�O�+!(s�2��K��#�Qvv�T3W� �7�#�q5�Y�p�
�E�V�B��0W���d���i	��Í?�G!���j�Ǜ´V	&s���>������,��_j���}��5���4��jYja[�42��e�tZ� �g\���,��"��Id^
��O	�
�|�1�.�lm��s��B��(��G�~�m��lq�&���Q��G��)�"K|L��V��`�J��_1DZ"���g $V
�YQ�]h*R|!p��[�J<xj��r�6_خ��@��}�̾Y�����a�����3�ցX����U�;���/������n�U��|,��&JyG��1�� ��K�	�Y��E�D  ��\��h�#�Y���ݦ� �M���i���M��s~J�E�Z!k��[Ϟ�H^r�; �v$Ѕ���7?���ݣn��k:D�$��tޖ���z��I\
M�RkK����^�2��ӧ F�{��o�(,%>����)�	V�.�I{�S�zBgTL!:�~F����-/�?Hщ;VD������Σ�W�N�'�%L�;����i�?f�E>�s�}^�D��s�w���`�6�nh�1�{a�E&
���m����=A�� Z:��|���h1]�?�B�(�-�2�y�T���C�A3��?!x��|vex��^�	��%.�7i�M�L��}7J�Dm8�熝�i�E����>��.Ңkd�0�`�H�	�^�N�k�i|�Oh�E�T� �~эw#����
~�5�sMTr|S�˳�GʜO̈́W��|����$t�չ��UiDwO�Ww�~5p���q�^��,��Ў�4�u0�c5�s	/��D�GtA��8���	0�MX+{�k�<;�\����PM�Ĳ�w��~�O�&��I'����H]�E�]�L�
�'.�����[U��lKl@����ؽ���1Y���O�19������� q/������\[�̨�rw�#e*�m�2��V�IK�33�ݽ��ف�䬀2)z b@(}�]h2;�����2o�"�(��?�߃D�Bڢie<���S�����7����l�}#ÿ�`��Njⰻ��]~6�������`���t��҈tQ�`�o$���v�_RQ���Nt�1��'����Ď��WO�q��=�	P�&�h��3�F�z��(�o���I�h�iL�'5�s`@�;��x�g�~<�����1*6�ʧ�OU,�ױ~�2�U���D�sw���l��X]��E��۬O��ݺ��G���r�e�*M[A9�Ο{U��ZK�u:|�ܦ�Z?(\�>�����ٵ���
�d��y`t�~���O�փ��wB�HB\�/	�z�Nw��%����lWڟ>n��+�۠�Hr}���q��LO��k�^���5��/����i�t�ʡw�PZ�T
��B���>��R�s�R�Pk�O�U<�==�M�v��HD�L�j�d�5d�
؏�/e8>r�L��h�$BeqD�n���ı�t�4����$��Lk�4�,��Z8�P�'.�N$���0��bH���{9�U>,Gg�n�N���Il_"��F#(b���8�m1$��9���|U/9��^�5���p���:��� �8<�5H0ҝ:)��ޑ �F�tOk�f�	�B}5���d�Ģ�;��F���A`An�V��)>���+m�o
��k���R7�����Bu&����p(C���V����A��׃5!w`%D��$uث�01t�nw�;��[���Xft�o�+h��ٮ�;!�2��js//e^�e�h;��d�����0>~�!��;�����:1�^=���+z��(��E��O��� 0ӓz��6@m)��?;������T���?��,r��q�4P�����FJy��Z���PA+�k����q���Ty��0��0�L5>m��Fa�+�V�>1��b��iK�����,�s
�ͽKN���	���:�S/�����#�/���1�������N��!��y��jD��kJ�q��~U~���y�T����	i:�d�r�1f���Z�s���_���G��([C4�AR�k�)�㔬٩���K�A�,~�7���0>h�c���T�b�@���KH}?R�'|
dtIs^���(Uz������' I���^�k�����E,��ⳳ�&�h\7���v�X3[*�%>,H�f6@�4�$2�IE�̚3���:��	������E?)u�j��)my�N*d��Ԣl�f��A�F�\
�Q-'��;n�G%~Α��Xϳ�AS�c�oo��;�ᎉ�{)<��TE��,��/={⹄����wˀ��<uS�E�+�.��'c
�R۝I��0fQ%��A�>�vnPEJ휕Ue�� �:M��Hf#D�N��B�ˣ�e@��v�P�_�A��N�z��у˩��ާ=��W����nQ8+z��ˎ�׼j>i�q�좆4�Ȁx�w�Z��)��C�!�����ϋx8���������oa\Z�"�)���#M`{Ȕ3նp;^pEPJ�&�B��&.w�,�^��r��dL8�����b'Ë/�}��<�$OeщkR���-���sx�hI�j}�(������.�l�J��MSr��/ p�Kl������jp?!���Z%6//���k#�Dx���gOў�Q�'&W��F&6�./*|��F�j��0�V�*�>�vتn�8�ׁ����7>����q��<�#1kc�\�Y ��#�K0��NJ�8�pZ	���(,��o���|�����ɳG��>�̂ ����Q����=�v�-�^l�^m���,�Ԃ�7�@��݄�y�T��g0���~�o$h��%�3m範"���u�6��̟
��i&.h����!+v���"{�_�>f��ۘ2�+��M�cd��(](h,����9��Gp���%�?�%�!u�v,�W
ǅ�3��>�y��٥r/(���ekz} u���q��6��,���l�����*����2%�J�6(��p�������2��hB����Ce��@�tY�m���NZ.��e�0r����Ə���
pzʅ�
H�r�/ΰE\.����������0�N%U�Ƥ�A��zn'��ժ�?*;(76j�:k���B�֯��D1wE{�>W���u��2 :lj�6�tǿ�(����k���B��J�|9^�)�>�^��,�����:H+o+U>���{8iؼ�<�+���q�=�*C/EY�D]Q�Hȓg�e(����
�;ᝑ��sk1և���l0X��M�=�X��<|��I-��	GD�8U�:�'�J���8�y�7�a��4G
r�x����[=T�Y�L/��s���ͽ{D�%Q��"���T���t�w}W��s�9��mC�iaꈎ�6�u4;;���p�F���˾795M��� 6*y]��N���[�!�-5ԓJ�v�s2?��]��Ez��ȳ�@3��G�ƥi��K���Th���:�m��c��'gЫ�O_�6���jJ@�D-�S.j{d��~~tħ>��;�]3 ��
���px�F<wQuߴ��̻~ (��^�����;9J�ة�H�!ڿ�r��ԙ��3z��1��>������y�АV2dhݍ�d���H��\����ō��Pڤ�#`�a�X8��?:���J,TP��W����Z����?Og1����AP���%`�O�ߧ�C���1��*�é�Vp��fr���qM\cz#e�w�ҍ9sP�Qs�Hi��1���+A�@Q�lK��l�2�R���`k[E��*}���0i��+�����o3u1�*{'�d�p�3M�r�2u&���Z�"�rt����$)�6�Q����dM�ߘ��';�0��xW�LhU�h�O"wŦY+"������K�(N�}�:�Vk�i5���_;�L5�DP=r���7�x຤�a�H8�R�}��A^�n�#�d],�������k{<����K:}��B�u��R�>�[�����
������f�p��@�˦��,�ENW00��?G�@X>qQ6��yK�(S� �,����k#�sw
	��fM�),�oU� ]���.��ˢ�=֛O EJ(/���L�,�!���,QG>cYU�Nr��u��<s���2��=	����S�&A�Dl�ϰ����hƃ�"j��a%��R%^����O'i5��ݴ� FP��-n=�J�}j�<�S	V�g��D���"f�1�(S�t��;a�g���7�KK}l�g�c�A��S�X�D�tY�_�%���(��@�Jydy5�������,ޞM�R2��ڞ
���
��O�հ�4D���V�R&ދ��]�]ݕ�
���,�f=`�Sn����_$�xY��Ʃ'��(Ff�dw�+����Q��'���H>�f#��(<}��7!�샶��g��?�_j�b\�������&�s�o��
���Q���Y8������{Q�{n8�z[�}���b�����5���Ž�"�R .����k%S����_�p�[�������~����Y���p�P%#7N�J/!~*��������1,�6��Q��$�8�R�>"�X�X��h+㗇6��Hm�?|FM䴭U��̻ꥱ/�����i�ݩ���[�F;"<_���A��@�#2��aT��4
d���#Ծgo����:�hMӫ9#f���y�2Ak���;�E���l�_S�����D�&7��X�.�^���t�k��;�����N� ���Ǐ�?S�P�4�}��
J$�wc���c�N[^A;�1��
 �uP�H�^s6 ��%i�p9O�ڎ������*:D��d#����� �������L ��5�+H�@v�PH�s� /��3ֈ��.rF_4���R�H�s'�eQ��pJ���1��d���ssM2�>�c�ި4~m�o�t�xV�t�(U��#�Wu�J~f�n��J��u��[Z2?nܟˣ�*�S4w
p��~Πy���ބ*��^�ia���ök7��<<zS��3���<��.fP3:8�c/���b���`��p�Me�R�Se(c�x%�{���v�b��P��j1Ug����Ϩ�U �$T��8硫t�"�n�]�
{�ـ*m��Aw��}1�E2���N��Ot��<�����U4���/{=N���׏gB�/�@�S��x �ڥ/��u�p%��8�n$T��0�X��(O�e�E�e��y�=sp�dKP]?s�p�Ⱦ��h��|��G�#���dv	mʢ4���$�)����H�e_7���ۂ��Q爗_p̷J��8�J�D���v�N~�����CI'=�|s�T�	O+����Zc�߭m91�9ĥ�B��%��D��N���U�Mz�mM���x�[?��6��� ��!·�Hp���a�����J�ైI�[��W������=/7̘m�nU[����l�𶖷є��瀗���Vȡ�����=Bbxj�Q��p5�x�._�$w�2���Z�3!���OQ���usQ�f��9��ŭ�N��zc�~]�شA��y��N=J���������"��R�/��%�O(֐�A5=�u�'|�ֺ��Иv��72R��Xzb┣�qL&����
gV����2��V�RoX`z�$����@ht�A�P�b0�3QU�o���9�W���P�l��_�A���`�Fv{��ʱ��Z�~���	��d�׹��"ר.�I5�f^������F�8�e �Z�������½��S�w��N�0���V�"�f����	�S���,� mK�!M�27�U��G$�J��ǭ��@O��Ssz�x~uU�ӺiÛ��Vb�f���0K��:5�%�~�Hse��i�����l{�q���+��Q��'���ׁn��,5�n�1�����ܖ����p>i,�n�XM���03�t���vL��oO�	�D�ԇ��`�f$ɓ�>(P����(7L�²v�ɢLW�oyƩ�[JCgB9�OZ���>��HN�g��l� �R��,<SsB�80&Q�Le���Z�M�<�>y�0ޥas�q�X X�f�)O>�B���.ʜ���Q4*�滧�E��=Ewď���X���d�,��<��_���I'��	��S��q����0ʿ��Fv��N&]����RQ�Sr�fɗ��C�ԙ� ����M�������+jsW�ʮ:Iٍ�H��/��U�[�"	��m|%�!�ec*��H�q/MCT��<��4C~�_i鱱�k��xP��(y�����J�4����J�ϴ���zL%.y��nI�@	����P�H_�me��I�o�����|�ސ����o��@F"��׀��S��ltQ�*�߷�\c�#�I�&V���\؟8�.kF���,X�t��������u��J؜�3
|Y��lC%D����~�п�{|S'D�����1A.wG]��0�bZ�椧V��:�e�R���P��ʑ����=�%kT�\����H�ƶ^��p�6{�����������|8��8E���Bj�s�tp������T��H(��vg*�Ф֎`r���tu�˼�VǪ�O��輳���P�R�w��(Hc%
QN�h�Vq����}�)��غ(��!ep4�%���׳�wJ]�0��|��p�30J����7$��RGo�PA^O����-)5�s�ۘ@�)�<�]�I)���5z?
[S���J����@���v?�(��'�8Eq��(֖9���k>r���#%�d���&�����RX�S��i�O�lW�����z���L��/��J4n�0�ſ��NV���b`��&*��߈�b�T�=:��C8ŀK���6s����uz=�OZ�L�5Vx�����i�1pn}�a[�w�>���A���@�h��e,ɝN�A|���H�`��#I���	X��㠁�'��0=���H���x5�]E��C���f�2|0�"e�D�x�Ҡ&�|R��T��i-�L� ��/cM�dA>)43���2��m+�l!"(J_T2z�s;�NjFg6~�yC����Ы�ݢm	,�h`��sޏ�#S��9H�T:����+~n�#�]^2��S<��k�[=jh馨���fE�R�-2�}Ic=?EMЁ�9��ș���aE,��B�DT���jtN$>ZMZ=��e�۔靶���Bx�cJ�i,��X�b�X���[�I$,��Q
��Y$�{��Ǚ8輿��kjY����Q�8���oA�A��j�6��Rug9�d��"*�L�㮥ڜx)7��:�oI"6� 
����6m<Afh5`�)،�s� ?������]Z4k�QH����v�zk �k�����*_P�|q��`#��0q;�!S/���hl�����ʼ�m�X�!��O�\�0��GVb�)��$<��	��;���+E;�ި�q�#O���&��� �0��"�^��=�����AX5�Z'k�Yd�N_w�'��j�3��q3��XJ��zH�<�@B�f���0�� =n���L��J	���O�Qm��'���ybΰ��Y��E�VO�@�{{�`��u�k;o ��'�9�?Ǘ�G�@j�b��w����[��K��?�uX�pT]2�HҶ���-=(R0��:��G��+=��ş��{(��T�`����x~A�p1o{+���*��y�^ɭV�A���%�-��"���p_��~�&�@f�C�wW��`��)x���ͅe��ړ����0ӈ�:��������e_q��X*��!��Ϊgք�L��e�5T\�d��0��J�|�d9?�v�I��v���E�c�ck�4U�<����j��j+LnGv�� ��T��d�*�4���eٷ3B��2���`{�F46?��㎢���u�/���<�����Q'�Òz��^���X#��(Y����l��ɉq/��h �A��R%����N{�c%Q��K�G_ �[�دVU��E ض�iO�4@3n�řQ�����:ĥ���)8d&��hhQ\��:7�E�cm���=y�����X���|�Q�P_Q�a?�(S���8�@H�Ҳ��J����	`z�^�4�n������j7	�xd>9I{�jK[�u�O2͊�1�d�!����Ys	��P�m��~���qӦu���o[֯��dB'=p޿�]� J�|]�Z�o2\��M��y�g��l8,W�k���^�3o�	�r�,ن/+�@n�gs١n�/��ǉ#r����Y�D�<���Z߿hgR`���}o������Mf/�GP���u`�U�\�&�:�k�GX�h�����z��#�)��r	+�W	��GP�(3�@x�����n[��u�8S����2�r�&�;^q� �{��OON��n"�Ftlm��K*3�t�΄Ԫf+�0��D �����xW��N��%|52͍�Z�T�-��� �>�a�Ǒ�RF�'~&�!� �-O����T� T����7M��&�\>��c�?�$�5u���ku�ZQx��0�Y�U�����",鯲
fY݁�gl��i���Y{:ʤ`�����'8�uB��R1����$	2p�QAA-��W&;�8\�]�X��I h��l�J<��*h� ,����g-�g�s�&��C5Zڷ�"�@3� �}|��u�y�*Y�>;Ӯ�;������o��d/#�F6a��թi꼧�P��L�%�o�V��܏�b��s�L��Z���[Y���z�@�&��Q��OIv<ŰKYj�6U���a��Q���_p�:�x�L�$D�Q"|�b^�/~����N��c��ys+���xX?m3�A�2�y���q5����ǣO.GZi����ໟ���>���M �q�2@0
2��dTkf��4��Uy��0J��}���T47)�ߗ��2��@�X��N��b*)4d���㘨&�uٴ�������נ�f����@�	���w����~Qm��w/��vmf��оS��v���⿵Cq��0��|[�����?$��"W� �2����{�
�iN����X���`���tF?.�'�`�B���@��x��U�J�F �W]�8Z��e����I5ږ-�Ѱl9�0��l�5*}b��Cs���i��%|<�W���3Пȏ��P&�%���BSm��r@��%*�kd�m���l�\hz�Z���p���>��~juC
���BD��^��4��NXx`��Q��i��7a]Or���fzQ�+��Ĵ�&�‡���=�^^Y£;���rw$���a�_t���8�j ��=ჭ�/�nf�BCN�bc�BL������&C����65����!��/r��D���ZjO���Qك�ݸeǔ�%x2:���9�݌}}N^�x�X`ɔ�w�YȨP׻���/��O��	�㵮�?v�k�#8H��g 5�y�">� rE8��:�&��5Қ?f��0s�O�����w�j�ّad��^e��ף������?b�M����@y�:Eާq��#�-;�W��^9��'�|2R�^9��ق�< 1�Q��fu$��б!W��3Z�S?{*/,u�RCR���xj���F��΋P���F�������grx
��vB�: �F��O�{�&i�w��m��-��/m�b�q�a��04����>�!���V&}h�ίA�DU�1ͦ�������x�C��Fܠ����'�퇰ÑS=b��'�QE�����E��>/"ml���:*o4d���%l�1���=|*���m�VT�~ؐbiجSP�r�RKhL���[��y���`S.T���0DAj�y�:�5��Cܕ,:�?��vv��!�|4�Z�cy,�Q����(@�Ay��G�u�uX� 󐹔"�Վ�bSw��.V��:�c��Ǒm��+��Bz�'��˄(���^����<t��C@�PR����6�'6Y��[�����c@,�h����պ��j��J>��١�����C]��"��<_�� G��%��*'����t�Zj��6�q�.(��P�š�M;�������"(7�x�O��A�V7��+����se���Oq�����u9�;uFN���Y�U�����XEdp�=���Cgh�{�jp�9|�A�,\=Lfa�ѐ��=�����;�Vѫ�0�`Ύ��G1��j�ِ@�h��TCDn�T:��D���1;���!5��P|a����	�R؃Sl��zm�Ab�,��=a�f&y������Nr�0��l���n
K��c󙨃Cn^.!���H^�^kN�gh+��y+��9�bϪ��⒤%"��`�]�{%T���+�S��Q7Sђn�ņ�P���l��Q��oh=ɤ�
G�J�!SN�ۼ� �����8�uc��So����>&c�dV�[�e�('i�Pn��
me�n�)�Sltܱ����������0��FiT�3��aEDV�{�DCfF	j�܀�Yk��5٬T��"����r�!��f��^�C��8������IQ���6�reh�C�dO�� hb06\�X�l}z��t�R��Il��U�@�l�����%?�򗇌����D�;-���m8~�޷~Yn���rd#C��;x��)*,#t��Æd޸��C?fOH���c��xJ�dG�����bI��}�x|Z÷�bP�zICʌ"�e� ��z5�|�Q�ڧ��] �Ďj@�6�~��B?�;;�4kqG���@S�k[&�ʨ�_���s�?�i�yT����jyR=��1흫9.�uM�,��YV��rOc����~ECVyQ��Q�]�����;����<�8�Q���=�qI>vo5k���7lHBި��Z��	��cua�y��������E� ��&�d1#M���t(�AX0�;�����\�Ha2����/Ăc���NJ	4ۜڙ�̤���-͟2ejw�r����&�CN\֠r{�kx��u|�W,��u���d�^2��V������9����]n�]t�◠hǻ�+��&]��|?�t2�K|b䢱[��oYs	Hu_3�_�L����(�6�}�Q��]�d�kpc5W����_��a^&&��&����7#����b�:YFn��`tp0w,Z�;�m�],L����!�v��Lsu�8�K�_�Z��s_`�O�eG2��߭šu^Z`篼U�h��QH��òm �>�fC���a�<?&��ՖE���v@�e�,T
P���Ȼ�
#��7�*<��s++����ɪ�������o������ɝ,�"�U0=g���� _
k/*�^ʦ[��C����!���L���@@�oU�5���WՊ�E'[�֬��@ފ�1�$��{5���Q�.�[r@�e7�m��`�f�L%"z���z��$���"�DN�{0�V!=�:n�����Ժ��_GF$���DБ�x���19��)a�V���&�S�|����رb��Ь�;�8�k�P�;8�WX��m��⽨
Q�{T1���R�b��0�C�3�X��d\8",��.$�D1=���­��`d��O�?|v�b��6wE�����F��d��HĞȘ��ƗPr46[N�����oV��]��^
M� �_0h�UY�)ٍ�+?-u]J�%º֋�\~^�� �J���q�A�nI�fhT:�L%AC��&�7�Q����ʆ�����޾��,}�&E��tz���l�C�e?1b�3BZ/nM.9�-�Z�ͻ�0�]�� D����j܃��-�h����4l��n��ć}c0t�BJӮ�s�f}=�9��S�S_�4��{޺��L�O�����6d��1Řv�)�t��ndK�Kj{-3�B���(��\�^�<�uA�	Q�#H��;گ$�ad���=�q��{UA���#G��HY�˻�l\o�} ��Dٙ6*��Sc��a
�Z_���y��*mf�4e+�/����{'�z�?*$�mO�we�Iw���S���G�j\��&A����2��u���� �Sn�d#XÍ��N���b#Ē�ɵ(<���7x<Z�f�P��� ���+w�q�G=���*6U��W�Ksm ,�?�� ��浈Xc��a���T8�"_I?��~�i�C9�c�[Dh���K�J�������M>�%;©�~��BX�� ���H���v[{Tt�g���������P�F��G����Eo�$��>+�����Ybs��M��n�&D��ߚY�R��f[�5�R�y��������=(p1UG:ȓ�n����X��N��ݡ����
��C�J�N\jtF�m]�X��j7PC��x�X�3�6�?����J�A���Ido!�O+�n ʨq���N+��8y���bw�����c��������+�sqfk�Q-� r\��G�7�׼p�a܀H��!>�\���]�̯o;���r�w\QU'�����3<g��8��a�'N�_���q&���
�m��� �]�p�� ��M?#�匞*&�$/���w8/�5<+���C˰aLa/��x5����{c�*Z9�Y����:��wS!��]Tt�5T������%�?�v���T;��M�K	j�j�c��֥I�M��C"Y�U&K�$��]�������y�V���Ux��G�8�4��Q�JG�!SwH����n���P�g�Wd�^�%a 9$z�Mj�C3�9J����TS�0�m����C��~#�j-��o��r�\��h�N6�A�� �l7*����7��/h�z��F�_j��l�������'9ݵ�]N��Z��u�dC�� S�V��(�T(�Fϱ���j)���l�KEm
�ֽͱ���M����Zpz�m��C'`5���K���}�9��6���q:y�V����2z��^c��T���B�-��3�r����a���\!3��^�R��(a��(�t��3�Ym+(s��U�v����Q����_�(��N�������Q�,ɷ}L�/�v=	���-էSQ�%'��d;�?.��
.`A���l�Bl?�`ǝn�+��[|���_��9��#:�F�+c�I��A�����0?Y��{
r���L�+�>����������^��V�0*t���a-,�*J���m9���&�(�aZ�$T��C��aa ��ډ0"������ﱍ��;l���4xY����id*�������H�\O���1�+�WTD:Q��ms��XК��_ο~�Z�t�F��d��(G�j���$�նiB=���|U6�?�e�9���B�E�Y�M��n���V��S�3�=@pg#1�s�u���q�#����� !�,p�OĤG�w� �l]����9|s���M'�H��h���7�L�h����bم0��n<��^��HiڞI$�`L��E-Eh���im�\F���&d��q��Õ��:	9Ђ��-�i�jL��sͯL*W�0�%�ԛ��aQ5���7���q��tJ~�1����t��sJ,�d~C���q���*ֵ������bN��i	�g"��f�B�	�@�o��>�e�Gk�ԺiNо:�e��c7�
vݺ���ar�Z~�RUZUA�~Z��/.����|od��}� ���C��N����-�SF��Q\MUiE�6C\9������Q�?9�P?{���9�w��ۏ��R��3������UBR��ݭO���.��I�����������KT`q�y���{U�|>��IT���S^x��0�s��{]6�Y�M�G"F��Z��z.���e��PA������f�����(�ưn#5K���p�E|�ldo��:��m��fӁ&�J�q����Zn�VY �J�k(Y���(���|�A�郞S�=&���r��\P2&V����B���0��d*N� 4Z�Kc3l��jq��)˕Փ��%����\v��T�C�d,*R�$^�-R���`�}���U�Dn���S!w�W{���{f���g0�RP���B���S^b5�z�Ǟ�s>�;Jj�z|���ۃZI�j��H;y���wT˹ כY����NQC'�p��<��g�Ob�{�P����H'������li�{$=�d�O>�S�F��/���a��G �hN�F95�+������Y�'�)Q�d����'���oL}H�x�������ז�|ֳE`j��^ x�C�o�A�M}�T�Ϊ)[tg�;�E��C�;������T.]��9�����)��x�d�63
�䠌� ��,���	25��kܓ��������XOhNߒ��a��Sy��2�C�"�x�D����Sb���G�(Cz�%x�i��:,��&�w��TH�"����L�pU%}~�y,��%�$g�`gQ�خ�u��w[�<�.�z�����n1��E4�4~]'���[.�*]�!)a�{=OC SO�+1d�CQ?�5�e�K�ȷ���7�O���)�J���T?2�P�T-�����q�g�, �"���lNwCT@/���B�x�������Ŏ6+�N�m_��O�G��i=%*�B��Z��w_^�H���'�M��ȋ��/O��ߌ;9�i}h����<`)S䗣�O"�?��$��4ћr�qLOH�D�.&�}$ewt�QQIg�"�>�~y�p�:~>���U�r�g2��x�5�w��R/d�L���D�TE�E�M3����yC 06�#�F��ZL>�Bqq��x-C<5�.��ߺ;�	X:0R��9��F\
��&�6��������� ;�i�b|�;���.��m*�͊��i%�:D���{*W��1m�c�#_�%y��9W:��U�~�glQ-[�Z���G�f�d��t�x�Y�EQ|b���C5�Tȉ�3��w��̏1�m������a���'|�����I&�_$�Y3<K���5g��){q�&�/iQ�tt-�P����Lz��Ta	��g��Ss=}׵{WF�u��gSv�@7	��h�z`+�;��y�h+���E�\�؈}E=�v�;e�_�4�k�_�c��o'7FU�˳*GD��2;U�ޑ�o�"S�J+I/��C��Q\�	�Y1�ĺIwS��"�nUk�{Ȉ�D��-I��2RI+)d��|9e��^O|��7.mJ� ؄�`ȁ��[��O*��7���ju>��p��|RF�"�k|�}竈�[�$Ȟ�ؤ��|�@��Ӱ�7��6x^��@W^7]��xsFY�R��Z*��ƕ����F�'Ֆ7�uW]3��PG �|�ν)F�#oU��Sp��1:�&h�oɇ�����a��/#p<�[��(�t�+���Ӈ��@x��I.��%���p��&��A�:ϡ߇<1j�5,���}���1����뾑-��n��rz�ά�u*�����	w����Эx�ؠT�����2hF��!9;�Q��'��`W�����C�7���U��ƔHA9�DF	�+Yw_���=d=�L���0wS�H����GYf|#'�n�o�S��Z8~�X/<qŶ�U�dѽ�)�)ٯ\�KB.Ŋ���eE'�=g$z�$�]3��T_�h���������PG/���Z�t_$�G� :^|��uJ�P���lR�7�%�Av�lt�^�?��aw���g�Sv�6��v�;ҵ�s��{m�q4/o�dAw~�h�j䭞�p(�]0 ����㊫g�*�x�n���kXj��3�\Q0wLq%Nn��.�6�iFKp1�]K^���8�s�_l(��� �X��t���fUĲ~�;�]��/�D!�C9ӟ5�B� �2v��,�O-�!E5>�>ZM�{����/����*�(&3̚И��)F�o>I�:�B�b�Ͱ���n���:��$$�>�tb�I����}?���mf��w
�7(o��p�μl���Шa�4xX�f.��P��1�v>Gg���Ф5t"�xGq��A/���8_Bp�3I��#lK���q��M�� � ~��heвV�cx1��{+;m�����Q��%�<=�r�˗�{�	s	�M0T0Xm�=_9CM$�$���y�$�������D��iպK
m���Z�g��_��5�IF�$1�pxH���R�ͨ�^�c���on��� \Ҝ�s�FsR�59�3�M�m�|�OQ�6��:��*3^{FQWP��!�A"��(�r^9��1��Pt`\�N:��_;u�:�7�$������#����@5X.۝����&u�w}��5�;�l�6��ͭE��P����%���������;g�����p��F��Tm��H�Ұ���R���-p	�t[E�)p}0�C��b@�: 2@���6ٺ2�ţ�SA�)�c��?/�c���!<Y{jO�t�'�.r9�xj�{���4��7�B�ɤyuw��덖W,�"�Ǆ`��3�M��BAJw �ZQ�x+�q��b��3~8�dǑ��{���}�d�O��A�#�������������xӁdw&�/8�b��������QL��Xx�ͣ������I���;��/��pJ�>��_����3q��2��>��\�~�K?Q��6\�n���
O3eB�6��Y�nO.�Se�eD����]!�3�����۬╀���';X~�� ���
�U�,\���v���{���hQi�)�Js�"V$�i��!��G�j���!*�����6^�Qs̀�K�0;���}�����c�M�N�H��U���n��B����9AO/�� E�X�+$�}U�NvR9<����n������$��W[3S-ϩ#��Pb�>Ǒ����3�Hz�W#�K!�s����
��&����-���Y�-`8�R"2�6������b|{1o/�R���vk�:���x�k	���p��(���?̏^��e
P�e�Ed��2Xl��R�o�ڈ�ebx����5��R>�r���T	A]��g�n5#�&<v�P/��n�Je�!�5�*s������-�!΢��Գ�&��Qk�.�w@s�8�,�ς� �X�z�dO���M<�7?FI�q�F$)�.޿R}��|Pg�����
�I�m�.��E�M���	��a%F��.A����a��Ab���4O�m�!E�@�ҽg��a�F"�c����>:�o������B�n0"�T�6g�83U�1P��s�k��$�.$3�!҇�F����1�����?Y�1S�p؆���8sgY��1���6���K�U���s�2V���|�n��ٱI6|*�D�����n͘2���� �N��'�/�"�/R�]&���p��g`�k
�l�OE0���@j�2�e͠o5�(IBC�n�B͂n�����1Ry���]�l�L��E6�,$0��";ږ�k<
���??�d����z�,�*t�_}�_^y*�r���0�b�N�)�;�6�ݡ3#E3��Ia��ߌ�٧p�E�K����[X�B���.Ӏ��_P8���)���k,�O�__W���Gsy�=����(89ua�@D�s&�V��a��Fvp��N�v?w�*�4�����?������zkHJ�N�=*M���� V��hQ��s�#�ɲaG"�v�dn6�'��Rt�K�ƚ��O�LF}]G7QU|/�����4>���+��2���X��t��`�ĀOn�S.A�L�����<����P`7�Scx#�Zb�[���=Dow��#)��j"xԻ�І��&-��V2�8�K���Y�"~��Ґ!s�b����u���>f�C��{C�����JC��;AM����GD�!샎d��#0�5w�/��`�Z*z���[��8��
�
�Q�vX����fm���S��f�Ωm{5�x(f=�ʤ;���-ެ��غG�Z���z���v�|����-�M� ������_���d�nPr�U�]�ﺺ Y�PB����)�������VhJ���
��� ���;i��K��P��4b��iT�������p^��0��"�^5A˸���vN�bQI�X�m��x�����䎱C��#E�iW\N/���K|�Ov���]P����������?�y�o����pK	�
]�
�Q˜���v[L�����9�K���*����g�+�$mS��k��,�]d�lVM����b��I�m�ʡ�x:e�����A6!Bd�e޾c/cB���)�B`G�����f���t2�}.h���DQ�D�;�����$��_]��'i� We��]V7�2~���A6X<�i�>,"����VY��̾�L�f�`	F�>#K��72���SVP��Hy�}c[r���*[%6��p=���rx7�9��.@���g��������X6��V�ׁU�	X{1���j�X���#6��C�	�����Evu�����񮩑�]�����"+A%	W[���m��>8�ֳba����s&�:����홁A��� �R��?@���4�Dz���OJ9��V���Qx�@�J�@6}��@r���F�f�1ݡs^��zȘ��i�$F���ܨ�#Ttu�&2AA��%@�+�����kŘ�X�_�|*#z�G��(�ط��6�R���Y����S!�8���6���>�@b��|&ϱ����[d*��]��%��(�u�R�Ce�mӓ�bi�=+��� �a����+�B�v`v�q@��π�G`���ח����S�����|ݱK0W�=�!�AHɂ�78 ���O��h�{�,\�s��b�������$�}9�B���J1|f�ۼ���{b@�o�N������v n۟�X4UP#���Ɲ~{�<,���9]mɨ����H��0G�1`����H�?���% _��e�[�'~�U�.���z�a�&;��^orE"�	9t���5l�Ml��n:s�B����yǠc$�`(�JQCy8i�h���!E-W�qC�Hy'�	�$4z��o����������+��p7�1�}�`�l�B�xšU�qW<�fϮjlɉ�v�Y�r�qt: i����݈�+��^�����yڂ�zܚ� d���v�"�Z�u�BD�|΅-���R�ɑm3..cV�CZ9��`�"�)����0�Եƞԃ��ܧ L��}=�ŜES�\��Lf�:;����A�ċ�
j��&�����39�%���F�W���bgW'bzYh��.���2()�������7���N��o�tmƋ���n:DKh*�E@���L ���H*>q��J=�	C��p������"�vb.�`99�l�{�^��,r���� #��Vv���|��� 1U��.�p�4�/ϥg��*�� �G{"�� ��e��$;3��	�~��,�ھ��z%��eZ�,V��{��S5�T^b��<����;a͉X�����ue�0���D�kp���ۜ�Fқ��`>��k�l�2�QA���ꜩ�s#���Ŝ���}��D"]D�˺�2 Ky�E& �{G��跇�~����RT��+2��6�b�T�lءk>����D|�b7�mt�R� '�'�1d�_d��'�z�j~&M���ᆞԑf�/Z=�GnT���E��0�fG������`��z]��ɳ���Ux�8�4�|ЮZt}^���E�EԁE�]�����Յ�KHyI>��d �k6��V�	!�8��"�X?���WSO�^a�$�o�|��1�r(���?�oV�iY�oȲ�h�ި=�������8��o�N���Rٕ�՛�������o�2�%;dE�HIx��ϩ*�����u����{,go�m5;<��}}�,��N �Xѫ��y�H�t���	���ܽ�,��A�,��N<V?�YrN��,�!�$xָ��E�`Y�seU� 8p%Zmw��z�lV�0�4)�D
�	.����P�o7D*7ܦQ6]�vB����k|/���.=�ܖ0��cy����~Xi����5��>��t=x$�ŏ�Q�"y�7V���s\p&F9e^n�3�J�IYQ�n�A�la1y� ����Jp`�+�F�:�qcE��Q�(��2��O�pD�������ݒ�N�ķw��]M^9U:�
�.�!Lg��A��b��_��A�~H�ŝL�ư#�i��ơ�x@��_�P)���"�6)�˫L�J��'wQ+� r� ��,��	�����v�J�6�����^d��!���(a�l?_�fW^�[�E�=�CV������)ءS�x��S�>G�e3Q+���"mV��/���+�]kì6/�ӽxѵ�h3�$SH����9�-X�%�{�S���ЃےB�����g�W����o͘�����=�,���v>�|����,�J[�#/��N*�
�0j �� �#�zq/�U��­�DC)�I���gĉ�Awx
cf��_�H?�k6�k�{��^�����z��}!�@7�j�G�B��[
<�p���T�I�xѣUZy�hƛȑO2�q��b:��j���ǘ�,[�Q|�o��.Om�9��s�l��-C,�?����X�)�1XV
��H�����ơ靴ds7J?�4�v40p�[��]�&�'�3��u�� L4v�ɺ# iB�����,�a8q)4�,4���guȽ��&������#]�¾�T�����ɭ|�jT�?�$O��BN��*�3���H�B�w�ZA��Y�7Vϳ^��D�K\�����J��O!Mp����ϧJ�^��d2?�ܤh�0D��)Om���G
��6B\������ƏL�����������I�9D<+�q5���v�/��\W�Ր�^Y�a#z�D���,�I���S0�����>�\Xq�t�
�Î8��{��y^�(}�Z��m�S�����Ŵ���� ���Q���.�D6{ �����NbdY�l'R#�������h�F/s�T��\��q��t?��$���F5�lR��y˓�og�jt׬�>��`i�X_�Z#��$y,i�u�5�̈3�$9&ڄ�惊/��a���.1vJ@�r��&�]�����]�v�J�%[)-�R��`�b� �S|�e�{�OuǱ�A�e>�_H��l�������`�&�%���wQš��X�p��bx�ؾ߶m참n�_�7U@;a�8sՌI����j�Nm�.()q�M�s�TU�)���wE�Ɏc�Ԯ�EPn��CF��πw)�ůZ�I>�l�H�̒�Ӑ%������` ��ko|����hc��=�skRy�D�~��l�8�dF���d\�@|C׍���1��6�uԈ�ڭ�Oa�V|0y&�]����8�x�8�Q"8��#��dF)q�b0��� �o�k�S�tS���L`���������7u�?��\��(Ͳ��� j6k�s��������V:���@��|V3[��'�"�v�1GnLk�8w.�O�@���naPD5���%#�@W6�Uk�W�l��zZ�uܨ6,����Y��E�u��i��Yv� ��	M5>�	$�ã�b3V������U"D��c�mi��9��$����vP	�Mgl��"�zS��	���eRQ
ԓ2�s/)�9>�5��,ݑh=���zU�
�֑�<�*VI��*�T���=�i�mm��y��,�&�@_���B=���YR�7����;TjNʳdƓi}�_M�*�A�
������Ho�o��n������
�D�C���:�}�a�%�
M9��Ʉ�۲϶x�(U r�h�;@�Pm�(Wѓ�[ɹ;>�9��	�-z����$p�D���i��O\��錟ԯ^!�D���ym4ը����J�*��;,:}�K�x��Ǿ�1�T9�vx��րT���1�̕_�lb������\a�r�N��iϳ!�l���]���� )�П�Z^��yu�DS�aN�K�W��嚷$��'`����CM`���Lj�Y�}mZz����$�E#��埿�\��|Z@6B�"6�gF)�Y�~~���t���t.9�~�ţ�����ެX)�0r��E�Y��b|}�`��b+�if�T���{R\��eR����(���㶎)�KW�@G4%�@�۳0�e�� ���hEE�a�ya�j�������So��A�T�������Rm����<�x�|*&i�DD��H�O�a��,R�-a��'��ķ��5��]Q;,�OZ�*�<��?q�Z߇�1�4h��HW�x�������C� ���f�$�eA�sm����B��⏯�hN���K|��Ir���\f�w�����ق��Ph?��J�g`n�f-$��AEtT�UҘ�H�z �2�s�r_=�b�'��������[�o":$"��C	�WL����5��[��q(�q
�O��^��6�އb���V�&�n�H�n�mm��7�dO�v%�|�6լ���8��B�Ĺ�M��;]#0���ѧ�ĕ״alt�:ޔ�P��5Uԙ/��%k^>�x�ņF�� @�j��Ԝ��R3�鼣��Bd����ZWcF��K=�� τ�$�'��_Y�WNRW�"��q��(�%|�-T��#"���(�Q�f�\6�ɏ�3f#S��j�E؂Ŷ�٨��C�l�&�^6r��O�V;Es6�l	��ð��E���0�P0$�dMֵ��s2�N��y��_�R��-��֐W�$w�+�e[��"?d�������n�3��܀�)�{�"}"�xI6H�MRی�@�H;0�:���^e�Ȃ�}�
t.�|Σ���|�=7䋹i�I9B���ʥ�L�@R��b��;�!����!zw�Z3u��|)A��2�mB7�x*'9�2$��?{r�E
�}��Ai�ȋO�㩇�S�����}R�"ښ����&��|ڵ'�*��gn	�k�un���{����Z�a���і��Ñ�$�q�{��J_�@�R��l���WoӼgޏ�,3t7̀/�K��H5aj�@�������U���y!椇������h�#}<��c��,l�g�O����zHb%��N~�Ω�DB5Z˗�0E�_��V�>�ӔiO<�F���v��hZ�n��R+Q�P'����� �^ ��GQ/��Tm�Ƈ�p��Q�r}1\j�7P��>d�N;h����Tb��-ؔ�VC�(�>+Y����.�`I�G�n�묅2xjcc��&�k�ܩD���P@ܕ|J{\ӣq����u+���pzq���$׿1�])�s4�qVf;Ά:�阥4ږ+���k��P�ă��XaDk�`lhNł�ӳS���!quN˕C�	��Iםn����[0�kXǂ
E[tz�ȴV"m�j����Ƽ#��`����b����k�y�g��6����t��}��*�D��%\���%[:�.c�fO������*ϑ��I��eL<_�sWA{��'�c���"C�)s�ι�/��C椯	O�Su�<��Zn�Ce$�͖Ha9ɷK�5����=�ݖu� �s��wg%�\B���&Fa�c��U��*M��.@\Z�ޔr�22�U�a�B`�	���)ZZ��ӏhA`�%�m^֞}���p�Go��h�N���K��C����������N��k�La蠖����.Fz*�6hkj&�g���~��S.V�e�@�#V��*Iy%�����PR}��#����JV�.a�35�P��(���0��̳B���Y����
�iI3�4���$��Ŋ��� �T^#�B���2�/��J?4�oE	H�Y����K�៧�0Z��T
O��!���uF�D.l���Go쨯�x-��d���zw3#q�gZ%�\L�O�vI�C_/�~������2�]�޷�TT�y]r�4������n[�z��)�����<�������L(�.�j+��A~>��|V>�h�W�T��krNr�<si	M���K��xQ.5�c��E^[+�vfX��dX,��f5�v��B�2E�3]NS]���`��ߣ����qx󏵃�{��0�Q�ƣ��<C$�@1�:�����D���Z�@��峁��Jg)���п�l��\��V(��c��#��o$��)P��W���-=�@t��T|q����_h���@ȊY�g(*�F�,�$�D<�R�[����(]Ý��>R�
j�5������1�aX�'H�L2��M3��	�G5�y�H��'�	Rf��/n�Ȕ�I� �� �|)c ������Ή�!��@����&�4����Rx�˴���ې��{L-UiR%.��Y�f��;k�_RV	`�$7��پ���Fv;�*̂� �j,�f���l�������E!�M�܀��'�f�_�!��@�^�,s�]�)�����l`��X2���/ݫn��`��LC����Q��ܫ'��#����K����������Z�����̏yp��^������B_���B�a���遙)��c�Sw��z�-3�7ge�b�-j���6^� 7��/#5/B��YB��ލ��b��ɴ�I)�����Or���ꁳ3hgz�M$��(7���6�����N��QZdsk���[q��l�ZYa+��na��o[Z�l؛���\X�p܀LБ��#|�!
�cل�_���{��nh`����2m�o�����6j��/C�I�+���ř��ء�fT ���ߦ��VA+8�h���
/B�kD��T��,E�/P��vx���m�A�4�%���#P�̊��K���~g��70����z;��!��D>L�a��hRd��я�n=�J�%��ksKF��%�@�R2�t��bs�_�g���%��sc?�Vաe�ǟ|�+6.]y�������f�8�y�G6��E�F�Q�T�0J��@�A���ܸD�Լ^C�\���A���__��+�y�3̅�vtG.}���Ƽ�*�����kQ����2ҕG㩽h`�ɀ�LL�5�����xD�֥��1T��W�1�����Zo�:�x%~פ��KM��wnY.�h���ԉ���W�%N����ۧ��6�#sH#��f�+��M�.�pprIB�X�s��u)j.�}���ٓv�!6��4�Z�R/6�����z͜���8������� ���q��)S4�ی���\6!EMj�	�G*��Z�P$�v4�#`���]]<��VF�3�^)^*�(n�W}�?D�v���=Y�$E��gA�Tȅ���/E�ȵ_\���91�G��X��wR�\,��[�J�(Sg�-AY��EэW�ᒍ�ۘ����y`�5�����'-H �1��502���n���;4�ܴ%C�z���6�GCY��\�\�g)]C\�hJ�:<����&����[6��{`�G�\y8�e���C�إ��dD�#4�Tș>7���S�71r:��&p����mn��k�rRO��'%Ӊ�[U��Y�����&Ӥm�l��������GP&(y�W�l��rOCX,xI�`س@��כ�<�������p���4�i*�?N�j��TcF7�l���M��OR5��¨׳we�H{����Ug��9.Av��_p�Px<�	�n�������H茜��"��j��|v����ct�pDA'Z����<i��1O����i�^CGx�>I�m�ݏ!rrI 8Ɔ����y���[_<ȡ��'*և,��8����I+����+��昘
H����R#��@_�ֶ'["�iկ0�]:�y#��.�RY��$�G���C�[�I��7%�#�[y4����x�T��a��	e��9da#`?�Ʌ���v�2�Z�<�,k�s����F���sB���t>�Q�h��C�A������<����ic��y:�;w�`(�R`����vb=�QK@���A�n7%^�[�w�i~�䧚��%r�hv��w<h��qO}*V�(���l,�%	���Ӵ���ު�7.�ɮQk�R:���=x�lq��'}	8�����Ѕ�[���ŀ�;��%	��>�1�O���u�#�kI�wBQ�̚��diö�� ���F�c�)��������tvk5!3F�WȐ�O'\W^2"@0�܃�r��w��׏����Gb\+L�*�s$�&��`3�(�jRI�~��8�|�W��j��<�{��.9Ũ(�U]WX����m��l�v����)�#�x�..j�� {z?3�wB��X���T������T�%���J�j�~�R�o�./�_�y��HBτT�p��iJ�/j ��2�(2W!D v�{�b6�b��
��z��)8e�K'!�B�ܣ�8��Q~U`[��Ym�"'�����@F��g�=$=�Pd@�ӯ0��ւ^`=oG��7(���`H��]$h
 ��5nu���)ˈ�,��˩>5�{��h�C�K6Kj �o�x��ŰS@Ej���%�M�z�V�ZՃ�[�=\�p�I���
͗o�V0%���R���i��,��L<��3S���'Ì�ո�>�b��Cy�mF�A�m�h�k�B����7)���ˡ?Z�m�BK����ʯ��6�5��~3D����\X�u1{�;Ip����	#�P�\,RG��s�L<+x#�Hs[��w�l��d��[SYb��g�׻dPě��s 7�YxqϬR�L�*�
�F�?��G~=������eհ�(<<�� �\0�_{�T\0Mi܄�M.�M��m�
28s��'={����<�"�A�S5�2�
:q�Q ��ɜ�x�☻"z�Lջ�hk�bm=h�)Bx� �-���K��#.�
�D@�He�/���{���>�"3l�nݣ�������V�����2�I�˧#$�e��Q�F`z?����){�U�r�u�f'q���s��ؐ�2[���#�z��{UχWT5���R;��Ē��"Vc�,Ȁ�y�\>��|���1^�!I�f/&%(#�*�������*�l�� �`l<a�s��,�:>^K=7>�;[հ}B?���V}�`�jH�ŋ��F�C��b�z ��'��z�W�R܁��,xJP��ᨅo�D����@�Z��]���5Ғޕ�FN�7ܜ��ʨ�U�_�kۤ��N�&��_;��$iu��?K#�qhB��Ϥ����dWi���g� _�V�h��y�(w�Ly숢��ND�O
�%pސ�(��.��LҦ�CD;��;�x|���,���|&�i'�����}���E� �d�*/3�e�C���{o�59�<9�����@K5���S"�In&��ݽ,�H��Kv�f͗�qqPUS�0}pf�G�j��;��z� ��D��b\(-������r4�;ȕJ;��?��תS`@&w�� 귥�+P:�lj�1��۬.�w��h�QكG��}�v�pd?�iڇ�� =Ks�h�o'UN�å������%U֎�B�=4&c��Р�WR�Sb��h�?"��ڌKŵ`H�Y������⯫�kc�P�����ֈ1��h�����@B���uS�h�n^�O.�Y���ǰ�ܮ#��]�V�[�@˛�X��鯰5�B�QF ��<�s-��jZ��jQ8�q	��kӑ*2N���V,��t���(�]^8�]p�x��2�[����iό�@�sl�����AK�T��tO����y��xW5�?����n?hl@�{�]rBI�q����M>~'�3f���Q�.���)�P
Taõus)b�{�cQ�XS���n;4����t��-L�@���}�1\}���Q��[����n�;��,��~/$�Cֿ�ݯ�7���4`��m��c�M7�b������,�	�3ฒ�U#i�e��9�<P��#��ꁴ�o*�YL��vB5(�#�����>�P����at�=�.�/�k�#�Bφ1.��bge�B�m+���J��ǧ�
�q����j��$f�L:ʐ-pW��}׸1�\)�P��҉�y��Fm��!�+J^����&����|-=�C�[Ŭ7����7k�r�\1Fx���D7�t ���®~�U�2B���}vUW�5T�8X�����$���%�=nB��JGf�<JO���?�i���������|@ϕ
������.�9>��mC�<�D&����Gs�`�޻�JP� 9��^�';]o q"ҶLf1Yu��i��kah�	�\X�)bg�Ծ/�������)Q�{�Q���+�=��֕p�*>vOp��� 3@�hz�<UWC���Z�^�:���=_z�_:�z�9��번LA�sm8�$�)u;�V�'ӌ��d�oʴ[j�רX ����`e����_5���`>�/!��A�ps��sXtp�ds�}:aR�A{���B�,��ӭ��˸�'�V�p�[&�S��GI�DLؒ�z֝���V=�k=�7JJl����HN�q�������	�nuP��;��e{~w�]p��� �
�}����-�%
�C�D�JM��xg�Ze�4�J�m�@j��ӎ��؛GHկ�B" �A���V��3Rȉ8I�tBXOp;>���_�X���~�4�~�H*/~%绘~ g�>��7���t\�6Zv2���k��
��}!=u B$�Ms�A��vDi|�5J���6� 50[k�kp�]b����;Xv�F�FK�K���Z5�_4��}ȇ��5��L?��F�aN����?���°3G����e�`�W�O�=͒��H����<�nu���0TX��1�~��LIX����*����� d����$�f���̵4��p����&g�=J��S+ϋ�h�sS�s�PXW�O0��FHV�#�N��Ǡ=��I��q���;���؃�7�~��y�[j] 	P��k�PY��$y������?Mܓ&~�>d�0ޑ%�Y���8L[޹��)���r�H�����ѿHe���ڀ,fm|v?�.�uƅ��<�/U�ڐ�>���9�������X�.wD��#y/���T���'�����5�_'b!�{E�-h/@�>u$�(L�pnH�X��=��A�t���n{LD�/����l�H���;���#�u,��N��V|�\�R8݇!P,E�S�>�FZ�-�N?��/%$��+���A�=���\�c�I�nJ�)��Xǚa�T��M�U���A��Ioh�u�_�hF3�� �4x�(O�ǈ�kf�Pv�h8�#�����*�Y�~�'R@�I�]�<
I'�02Cb��2Y,ʨ,�הp����ƺg�?��܍�'�'���'-xN��q�476�{(t���}�:�Fa��Z�$h��"��xt����xR�r�]�Nx럟�n��C?I�?e�_v���[(TuD��4,V�b[��'�e� ,�������ߕ)��TF��"����p\��x���us[���o����Rƶ���,�ZFP��e��啺��5�'�W�i���/-�ϒ��%�ie2��ڕ�.������n���ml[�v��%����~m�M�X"[閪��Ç��[���'-��IK<O��~��MP��JD���݌VC�V�]�������Mi��v���ݿ7��_���C�F����^��a}5H�~�b�gK]9e��c������v��.e\�Лe�ke��x�bm}������V2b}�4��b�]S��#}i��\O��[ =�9�~��?��}p�g�^̬;�In�a�L@$fVv�֕��1p�-x��D�O��]A��T6n"3=��moH��nh#��(;�$"����i]a=w/?o�w0�M?�@��)%߆�ը�j_Q~Jp�����լg���ȁ�G;Q��^���\�B{��!<a��A�?�r�K*ҝON����7߅���G�/n[&hZ�P����9lq�kP�TH2nģk����ʱ�L6�x�X�s�z� ��/ܠY���&�9�6����nlU���%� ��N�1<m��ʻH��q��x\?�#O���v��౰wA�2(ΐ^l�� �(�z�/��?�?Z�"oW`��&�ȡ� IV߅��n���	H����K���FD�&����3��g��1�Z��	b�<�Hdd"��[ҷ9���G6�ߔ������Q*h\����-�%���(s��/]�H�AEQAg5���-�>��-�e�+f���3��\�{퉌�F=����п�=�Q�ڴ�Հť������YCx��ɐ}6���_�O�WB%���ࣖ��� ��?AzO"�����sn����9����*����aoE|�.:�b�m��M(y&G���=)��snG ��I�,��+��
��9�-��0���Î�vBS�����{����gڃ;�kZY�!�qBp����}H����Ʈ����:t����2;���"�`ɣ��T� �w+�b����}� �� ��rE��8=�a�2��0qB5M��7��"�ql����3I�H��� qq�����ڧ
��6�k3��ά�u�������'�G����o�.�N���4�D�D��p(O�������V%�i(΢=�����Ж��ڮq;J�[1T�J��@%��s3,l;/ڎ{T��훱>��߭~�1j��K�ԭvV�;�-��ZJ�]��|d��;,bF�[����������4�ە]�_J��Ǽ�8�&�����>����N	�� 4�݉&��L�Y����U��{j*��Qn�M¾,��dgĮ�$�b�ŀfGo^��=���E��r�R�$!?j�V�_�0�n]t�O��Deq��3Y�X̰��X�W�§T,�x�$���$�ī�y`��VF 1`�F�"�|hܟh���J��I&�6������+�%�#��(����l��1��%������%��"�E)�6K�}(��2!G�N��w��Oz �ӋZIX}��I�uO��0_��X�� 6�~=W[%�sg�.$�=΁܊v}O�\5|ԋ?qm���T�
��Ӯvs��<���g��χ'�n42���t��儋<"�K���tj0,L�e6;A��p��\޽f"$���ͦ�v�u�M���|��%�_��=�(�p:`�N��23b�S�G��iv�}8�<Y�B�|�z-��:q��4�[.>�;���t�=��٤�����c�Ia�L[���Gn�g�7KY�oQr��."�.�l1�uW-�{�w~@�-<{-�+�tm��$ӱ��v�>[���x����e���ήuΰk����Pي��ӮwԷ�YN*��Zu4^�!.C����;����k�qV#mޏ<��}~�ƀ���)9ŭ�GLa)v���������H��)A�u/����h �I�۶Q۵��	�H�E�'��(�D�+��C�y���}+
�'��璕efYb̊�kE\Ώ�+����8�����`�U�q�z�S��H�����N������/��:�)u�5Y1��e}�Z���i� 1��w+�Sv�B�C���S@^;��SfSG�[���|��������W��[K����'[c�-����|�M���YUG�s�����y�ұ)��� �~�7%����m:(9.�U�������N�`¹��ܜ䝬�!4N?<wF/`E �46)��bR}������6.O�2�&��Y�p��E4xM���)V�rv!���>F�F��T�����˅ٺ�	$�w�A�.}�on���lы#�_��ERO�gC��2�ݚ�u1��j�q�`^iy>�k�Ş�����J2d��r�6o2%/2��������S�*ǹ5U��0�u\��8�����KE0��$��W4If��C��B[��~um D�ƕ��߉��g�8~]t�<;:���iM3:>'#В��_{ޙ���WNk� ���J�sm���KqԮ0ݙ��CD�&	���iʖ��������$6z�m��_���ո�����(}��+�K]�V�������:��������"������z�(\�cc��Z�9Ғ�q�\��C?G`	(M0��x��Q����A��?�B9�~r�_��+��fc��ǿ$tX�I��҃�E�&5w[&����`�=�$=?@�*��v��"8�.ذ�b������Y��������R{�����UN����wr�Z�0�){�y"T��羞'*��������˕�Y$�B�^2�Ku$/��)�w%�\{���_���߁��B���`����#u�n0I�ts�Q�_&�Z�4�H���\ǆ�e��,5>��~�m���ڦn6'�	��?�P����I6���Ѽ-����N�P��kG��Z쌃�*��n�~H#��:�9�!���7�8����V��U��ii*%+#O�t*4b
��ʳ��d���&]�?]w$�8�Ў��ԫ����ak"m���/o�`�p�2I���}�#�&@^K�1g��Q���ae�q������%/�J�(�t�`%���p�I1z�:4g���=3��c� +�)~*���o=(��~�dDB��k���vNz-!���@_�=�����	@\6w�3�+�7}���pH䢥�Ǎ�8�ɝHy��-ֳ�����\�%��I=�\� a�aR�D��(j�Y��Qt��/�%ĉ����r��]��K�4������� �ߺ,�[\(gi�����H$�3G�, q�{#s�W9��������~���Z{{�`��\w�\��*Lъd��t)�	>���E���$J�NvP�jQ�/�b����l��,|�!b�k��j�(q��.� (t�4�qMw�yR�`QЇH����p�x9�x�.;�1�^���K��Vv�\��(���fjJ��^ĹD�bUӱ�͇YQ�rMeL�P��S^f�	:���7<*Ǘ9���;�׵Xy���wS���=Nx��2m2�[4o�>�>��g;
�Vh���Ԑ�ɱ����ҋ*����|gQ�q���G~�T�\�J����d ��W��̋�SC"%���+Q|Do 2�Ik��)��?�� w����BLp�[���F�ĎE@gf�7�^!��c�0�8��,N��sC�1���Z�	�ߡ�$�(ҍM_L�Ռ�j*�6+j���lr��UC�'�>�G$	��e�+�����
��z����㵴�`7��V8:,wQ�sg9�o�N`���$.�3�� �HB:�{.�[ ei��+�űyR,*Aw��`S�&�J��#�97���#��,I>�j�$G}5O�
w���������q�Y���2	�5�м�1��2��b�J�/�$��~q�R;�F�:�B�%H[���]�dR=�1����r��E%7F�s������H��]N{V;�����J02���а�,STrx�=S%�5�xt�nmq�$ڰ,8�;E�}��U�a=|_�������N�ɪ,'l�q��[����Iq�a�^���_��>�o"A�A��I'��kԾm،Z�%���%��N��"��%�̻��v7=_��D�1��>�-U3�yIO����y_y���\t�����ûb߲[��z�m��{���=�����pXYʀ�p�H�i���ߑ�	](*�l�j�BA1�^"�;8�(sj	���NVG�Ly��Mk��N�7� 
��$V�3��/�S�4�.]ټ���0��9.�Z��R,K݄̯���QV�oo�K#�ڡx����;f���فZ�<,�q��#k�Z>�=ݕ����o|��?�j+��RzɄM����Jl�M�䐦��s<Y,���3�`ӛj�fE�����ٌ�\��F)l� ��(4�G�4;%�	#*�c<F�oD���|�����_�>_�i�5�lZ)�f:�j0��`��D�릎Z@�VBȪ���E��7��A��Ql���������fL#�}�{��Z��`�N��޴L�G��`��>>��w��a�_~��$�{Oe~x������I#��l��v�4Z�ښ�F����L�e��g�_6<?��>mj�E������� ���d��	I�2�D��P��e�Ҕ��&��.8���0p'h+��}���ud ��o��Ri�ԾL=���������-60��ҙJ�yW�e]�ևVN\V���&�i�UMҖ![w#7R2����ң�$�Q���jv�FNI�f�d�� ~N�y�oO�N��2�p/x�����n��R������na�N�|�s%��p�읠6߹73�|��n��D4c��Y-�>�۰����c��"�K0�}���W���+���<��(��,���uX �=cQ�OJ��4�j�}�i�&��V8{o��~$P���2_�,�9��]�@�'�@SRrh�������^��C��34k:�BT���vI��E���.��R3M�j(3�7o��$/|�jfœ� ���:�*#G�43n�y�Ğb
?7��x�Y�����Er�O���'/�5�?TU�A4�(4qT�V2/��t��˳��j4��'�h9�ꈄܒvYG���߅��5�g�XD9�y`(���܂��*_
>�× ���Vyߟ?�� P���v�<)O�TM4b�^���x� �KwQt�	D�7�l�j;�R�*љI{�M�
|[��������O�Y�Bzݕ� 
��O,�aX��F"��ި�X?��.���>�W�Ә�b&"M	u(t�Y?.�ȋ�3��h�A��ʆ�
A�-#֎� A� O�f3����A,0ϋd|��t�1�L5��7C�-#gp��j���.�-o���-���'6m�����h�� c��hD;%����0�dr��O��C
��+�{��x��t ;R�$X��H�Aɛ���d��\ AZ�::k��Wf�^]Yq۞��ҫp� }{������-���BTt�_@x�"a�~
�����Hˎ $��r��I�^�a�?[�k���[+Ĵ�zt�{����!��HW�^I�v>�#t��kj�e'w<����)�@�����7W�j��YB�
K̬�,sY�;ܾ�Z��c�X�:5b�4v��z��1��M�]�q�\Xµ�G��a#b���<���E^2B�N'X~T�7�86ݾ��n�UV��5�	/���zHj�2�y���E�I1L�h��~�A�M�d��:p�L�����H�õP~8
2�s�֨��?p�?w8��-tT#H��v&2�Q�O�?����Gw��$�_e�<:kc7�f�d,Kq��P 	��pϧ:6u�؉i[���Gd�ʄ�d��ޠ�[�)T*Dq
�-FҖ���|5{L�g[�%ӱ>�!���iE�TN_�9q�&h�c�4��r]�C�9�����*�g���1�$����q�מnQ�םN�Ԇ  s!�ʃA�ĘO-�n���v��uy���I��QtܲW0���� �A_��Hչ�򨢓�Ƹl�:黳3��b�5�c;`���N�x<,��w�9��^mD�>�FR~��z��[,�8�`�u%ԼN����}m����PYU�6ᕶ2�4�Q�ۤ�yݼ���nQ�FO]�wA��ވ+�]j��*�(����k��TtѶ�o�J_҄�CcL�(��>���W���2A'��@QT��'��~�8�̚��]x��B����y�#,��`	;b��"�h@ͨ�����ƻ���Ϳ�G��<<����Vռ[X[�/�7��#�73�l:�LB�m�Os�-婓�@��}�z�l��8�)�I��v�hH�ڷ�/f'�X�����Ke��T�������1�t��_@�l��4���A�n�`�9�_%lJ#�����}B��KOe~���h��d���ۍ�B�0�Q�uB���SՌ_O[����^����l^�+u/�x,@�s�M���Dq�Ǻ�����	y�e��D�X�ޠ<�R�%�D��r��k9�����L���q�h�x~�+��T�����hn�6`E{� ��� �xk�[��J}���I=x�}$@�.Q;�q�~(u�7յv2��R��g�L�	�.ळ�l�C�jv]�j��)���8G�6�x�c��8���~��޸�%Ԡ�8�b�� ��)Ɏ�`[D�C��L��8��	�z��޺ՕW���(
�Iv������M����YW{db�B+���Huh���]}.?.H�lN����������*寱|���om?�eP�o��`*�kۣr[WkO��5����̣&���I_*X/f�m-����=-�xL�G��ܐ%��F<��?���M�E���m��S�BH������=��B(������b:�cɉl�|���GA�l��&uj�sf�8�+�.��Nѡ��F����^^�ڤ�(��|T�����lo�6�:���,-N��R��~�R~�/��>>/�xv��
j��ْ�VD|M]_�>��^�*��2�	�Q|���jH��*�bd{i��Q�q�D��y�b�Ԩn�9ޱ�2�Ń��7l M���Dܪ�h�7��`F��}��&BhO��NJM�K���N�RC��-�J��Ω�.�Q�!���\��y	�28j�����a�H^��7ҁVM`���_o9�W|bS�'{�[�Q�,��	k���Qf�����e��ڪ s$���p/C�5f7�=4F�X���y�4��R+�q<;� y�(M�.Va.�%�}|}����u*�,���zƁ �9HU[* �4��*m�*�}Z�I�U���M�O;h�4�%lJjp��=��D��ͭ@�4"����Bn^�p���(��AZ�9G�=������i�!�*�P�66����x�~��*r2�Ho�g�2�X��OEfoh�H��?�ʩ\:�Q%����eXj*h���'7�Ui=.�>����o��N�S!j�p<�7^��F�ub�E��Y[fW)Z�9ڀ%9$⑽�5T�uP<"g�s���7���/[`f�q�����[-����v�2:ӣƓ۔��G�im�ȎG�/R�![��Sb��fyFy���_��#�$bĿ�J_�>B)��"�p�y��Vr��/B�(��.(��N;݋�O�o��>�+�H�փ��q������@0}�8�"������4v�4]A�<ME�n����l�K�j����,��n!���Ü$<0����s�k�K�Hq�~�/�b��֟\�@>��2
���glbQ5����tfd6����'�X�0:�OQ-$�1@�E:V���VM!�T��ʨZw��f��&Dތ����{R"D�5��+��iꔒ�1�����շȞ�`Bi��y��>c�	t������L�R��V��{_"�g����w���p��L��D�����͝����Q��o5U����[�Π��R��'!�������Xy������)/%B[���0@,s��*b6��M���{��4?�7�5l�G	/��'����X̪�Q��,CE�d;��x�`�n4��H"L���:�+Or��o�V��SŽ�>c�:��F�i��n��]�*��:�>mZ����i�h���	7o7�Wm����f&#`.�Y���"�y�Y���M��4�Zpc�������$ͣ>N-�<��rE�;UA�Ң>��ذ�we��?@�?*n��,�'�0�E,�ʉ��6��{1��j5 ���h���&�����w��4{na][7%����a� ��f2P�zLT�/��|�r��m�ެ�e=#��!Yp�#�t�:P�*3xi�X�M#9^˅x	�?u�VC۬�Uu'���w)�`.�a%�U3�s�|�0l��:Z���d�r��Rק��G�kw/c���5�wЫ�S�B��a+��O��=%��j�p�ְZ��/NɃ���^B�7�D�0������x�^u��%,�G��uǱ���L��M�>�<Z�����/
�~	޺�*㌁ك!+�[$��08�J�!	�J��1�.1���W�qVb�v�7[LS+����Y��Wc��I ����}9�Aaܻ��W9���$J�ߚ�����)<Wt��2kYpᗪ�9��:(�(ٙ��]4;h��WV�
��$6_���͛��6�ފ�F9���l6�'��oѤ6eۀ����?ڣ]o�~�����+j0�uOގ������
'��c(sX�1��b �p�$D`-b�����j� ?������և�}%���z�r�,��xC��<,�hP�}r�]���49'�7�������GS��Ж*���K��IiIs@".�
-;<+��AڙcM�t�v^��+�n΄�E��Ȭ+?�����m@����(r�S���c�˽�w8���8��ɯ��C��2�7�	�����f,��5H�M��Ť���	�b�z���gw���ڙa3��Tm��t�U
Xkz���o�G��9����G�0L��:F�kR�5������|��Q�u��^�;`�ʣp�'@�t��1Jߣb�\55vj��x�Pp�+s�Ђ�t비��������I.g��H�A�c��$
ѱ�!�jP� l�&2(t'/��&Bh�n��+c��ߟu�(�ȳ�di��vu�#���X��OԻ��S���̗�$���T�bGq)Ya�<u�:,�����u=9z��N�Znq���k K���;���|h��.,:�y#��`=�o6�s��cַP�q�Á�5��[��`>���X�Ņפ�J�1?[;��K��c�a0K,-V�=��|8,�+���������[�#ɇ�h���n��b��4�U�S!�.�Ķ��Η�hWmK���n�K���2 �pZ���|�4�Y��E,	�N��?}*]n[���@�-�> 8iv�J+�+R\f��G�m9-��?�·^�}:%��n�Hx>E �z98gb5���*o�wK��|�>g��N���̓�8p�0�����.OFr$?�� �����;�a�,���%��ۑ�1��Q�H��p��x ��ZE��Y�e��h~Z{Cg��2Z���ه��ԓ����C({�&�X�p�4e��47����D�E�]�)s��GБӸ��2!:�aJ�(W>�T9eH�u5=� �Kq^������a�^�eN\�&�Dc���X}aY"Ϗu0���ܿ�p���(]K�|�=��6"0N����@*�bh����F$���z��6��y�b�sO	*�����N��S[F���sbbT]̦>>�jj D��u�F9�%��3f�yP�6�//��{0���^?5�3,�/T�A��ы:��-R.f�3V4휣&M��so���2J1=�Lu7�q���� �v(�ƺ���)�kbm3-$l�ګ��t��k����*O˝�֬�/s�ﰆL��iqVX��OP�ꬭvW�L���㓎�(��h��K3ٛ���� fk������1v r)��Ub�e���FS��%5���j�&�GLo����Q���d3�&>�ª&�&��z%Q�N�/<d�qg��v���M��Sf}�k��
�G ��m���)����<;	�;q�B�M)�皰w��?��Qn�fف�^9���e�E7�뒆�5/C3��+�3���\f߆�_�"�:�f����=�v�5�ti�n�6���{<=�?�C����h�ν'fNZ��Sb��pĦ�����r&��b�6�b�*�ʳ�7��u�9��9���>Ӗ�t��G�|C�V�#��	�f>�2��K6.?I�Sq��=Yu}�:3*�c��� N�Q�����`q7
"��)L��E���b�n3�T��be ���>ޓ3I=^��J�K�Bdy�7]4��\q����
v訒��L��,���l���];��PqTW��kd���B�km�M�P��:�#,(��s��c÷��#q�Y������Hi��N��)C�i�%T^"����5Ǹ[�ˤ)G�0Z?2X���U�w��a���LN�t���W�� ������k;C���g� {g$��-� ���j-qRʩߌ�>�)(�;�@9�]9>2��/v�Va)��C�M �S��9�I��ѫ��2�si5�'����q�0�x$o�U�E �+��B��YWH|�����hm�R��:���pÁ	w�񼾒"�K7e.G�Z��ە���Q����|6:�B�Xjh�43yi%i�JGlo3��\�. W3u9�����}4�*�}Nm��o���k6��u }���B��M֑k�%�	����@D��>�d3MI�3;���[�=�w�X�����ܩ@���TY��e�w�n1�1(H�0�kU�O"��4!i؍e���}��lwZ�J�|?<��i���iH�6v��@宍'ɣ�	�Ī�L��.�]��#�o�ێ^�+m�_A4�|n	1���kfu��>Q0}灋v߹4��jFh�e�z^� �r�KO�X��O����`�j�$�^u�ϴ�<6z���~���|¶�7��u_玡�ռ��J��}]��K�xㆶ�?׬����i4^߰�Ǌ7�R���V�&O���z�َo�Y�t�DJ�g���'����n"��?�ٟ�����x[/y�z+4�>��h�L����wN]���_c��^���dC���viyd����"ρ�}��B	w����w�-��4��x,���U�.n����=�iu�w �sN�MkؽG������'G� �I<��%�)���EW@�����dӧA�p�F]� ��E$����c�/�����8~ϫT�,H	Hq"o`_�ۅg�G����-&���L���w�U�DMn�X��g�3��D�r�"�)pF� �hc(�ݥ��v�n�Hdz	bk��Ǵ�$ң*�5X蹼����=�L��U�\n|���b�Ϛ��ӣ�����u��m�M*jr���YV݋Gb9eE���ʠN��.[�l='����l��_�z�Hz|������-As��������6�g&�.\=r�Ж��n)W��V5^ꎶ�Zy����ϫ���n�>�6��z���ߔ����=�.��Et�Z<v��ϊQ�_��w��x�:���L�9�e�y��}.s�����r(_�4�)�@������
�Zc���߾�ڛ��#x���D���w��xb��ʿ���,g�p��A���O��?E��?"qVu�i��8T��c�ʉD�]J�b.�\O��c�s?��+I$t�7�So�i�P�5>_��u�L�tyU��,����)�@�W8f|)Hb�� V�G�i�t��a�kz�.Bv��3U?�ZA��܎�>9~���o�p�%p���M?�J1X�����a��	3N�^ G[ 9�H�k�{��t=�+ԃ�T05�̷ZG>�G�	��O>�`M`�D ��ʮ9^�\������$�۹��ZK��q�]�_`Hg��i�dL80��+NSM\���R��h^u�X,�6�/�_��X�HA�|��p�;���c���S �}�Z�P�	ؤ�*�<���α~`t&}\Q��d�t��}67#k��ud2	��o��m�FT��0LH���-n���
gٰ��@[��Ax޿��`bpH$�q��C~.$霘B��b��_�0&֙�Ǘ-Uo%0�� ۅ-�N���f�!'f�5� 6�qF�"!]��[�Т�}[cO[�=v�H�������[%b�׌@�2S�X@���N�˝V ��CPRQ0����%y��k
]x�>�\uV%��;�[Y��)_�?f���$�j������v��9��j��AW�y0J����b���(�D��6�N�d�V9��eى<�3����L{��;f���A�#pܛ�Cn��Y�\���SPI%0�_�Sk'7+I�`JCjw�Π�hT��ϮAס�
I���vjWv�P�7��.C�l #ȗ��Cp Վ��v�� ��UY�%|�eT�]�R4N2��Vd�sY�����Vd"�mOKg�nL�E�������5�>����&�D�)OBf���t*\�ɩ;Md8�X;�v�eW!f�)� �����Ԧ�8��l���Y$Q\f�}{2�)�ˍ�q�Sg�i'�8�T���!�
g)��FR�W)+h�"g��AY��Xy�aN8(�'���5�b��bZcil��I��)p�qx�ce��]�Fbǩ�c�ȁ�$J#&cr|�, ���R���pvO�]z-��@�*��y�m ��z�'ݟ_`Ns���E�2�CM��I�E�G0���{���$�0����R�9��O}�1��T]����P�1T�j�	}��=��� K��0�WL�r�Ͼs�����LV<��`�`�l�!ccC��"g�À�V��F��6����5Z�J=��^:	Y��_q�/Wn�|�fc' ��"d�s!��I���7�I��y��=�`rY3��o�k�6�4L�g����&��������!�q�R����^�-���$J�i�<���V�P!);���˥�4�q����̓�*!�����N��Ӈ0��_�\&�r�\^��:{������M�z�G/�HzT|i�u#{lg|n��c�'���z�S�Q�d�49��=�(\�B���o�T�~dRLG[��gg4�G6l�Ee�>�K�C!��`O  
U���c�Mx4�9�����^�p�;�\ȇ(��r`�ϱ�5�Xg�+�c�iJ1�'�̵2o������zP�J�/Q��i�U~(�n��(^��-/:*"�7uc�[��tq��V9WA�q��l�~����t�5�(*�a�����{�g9��^nL�.%$�u��FZQ����6x��d78����L��g#r�8̲N�}P�D�6@�Q�L�v��� t����G��I���$F'w�!8;�Q"a/0�����6��N���z��*4�y�[����#�V��+�_1���N�*w ��E�T?���3Ĝ��b��� ����������f��2�� {܁[��u%9�,����FqR46���~NVg9�'o�};o�X�>f�� o�	�&�>y31�U^Xˋ^�@}1�
}Qb��بZ�����o�&h�t�Y;,s�@n*�;Ih&�u��&�?��Ǩh���>=0��;[Z��#����}�z����4��O�a=V�i7_�����n����Tp�%҃��w.������a�ui��"nh��e�~�����d8�BP�a����;���-�'z<��ŏ�:��mUwi^�hr��P�媆�CV�-�7��}�?q���߭�W���Ix�6��H����嚝��3�U��"Ǝ��0-��r4]<CA7k����3�3����C �c���H*\撿yj���� dR��E���a����1pØ�<���Ӿ�"_��^����*�n�0N�7�gc��"(M�f���f}�ĉR��}Y� ={�!a1��m> ӷ_z&�v.���C?�M�y��υ��a8��'Se�(ji�ƘU���H��?v4Eh�BM��n}��6Bp�@�>S��Z.����S����pk$��F9���\ �}B����إ�i`��C����_B]���
�䍸�kV4@��ɥ�`-�;6��Vy\�l#��%�]���
l2���8��zjl�ޗ�-�ɆO��OytWﳂ�uO�l´�srv�EO��<���`@v�W0�Dp���Hg��U�A�<���vk�pH�S�����ѵ� x�Eg��x���ꂍ🛴���i��\3,&5�#��{���0 ��l���L��}Q���a�[<�T�\��a�	��M��YE�51�֮C%���.z{�����ӰrU����SC�i�L���XdB�P���-nQ�%Y"�y�5]�S�K�?&-������g�*���j�Qv\����Pu<��mv&�KS�����:~:�m�P�9C�|��YLP#G��{TuN����&�B���"��������ej�+A�ݹ&��n����N��,Џ��Q�2mîs�T{J�"ߦ��'<����n=�hL����{W���:�ڍ�vHK�����)D8�G�2��
���[���jY?c�&��h_V��P{�F��<]}� �������!"h%��������C�D��G?ʞ-�S9�Wa˦�D�<,ZRr��lG�./�G˴g�;` "�M�Q����?
9����.���I��)���Y��^���:����Nl����Ǚ��!P]���'=�ëwe�2�`��b�^3*\Rgnە�!A{�Y�{�3��s�����6"nh���j�|��2���U��JP*l1>�a�<�_��c�*����I3s%FO���	�@���7¯�8	F3�m� � �o��G�丙�ap�4�:���t�7���<kx��g ���t�8q)�Ŋ�0^V%��ϧ*�M���Y�ej����tHxY/����R�H��S�ll�S���uļ�C���s4 3w(R�*g�K���'�P!=&����Gq�Б�J<�b�GzH>�����V��,��t 4k��i�s��k���ؖ�Q�������%	|�#�m��
F6!�(���N�c�˫naK�L�.��P��$�(q�قP��hχ�B�?�jT=�����V�A���Pwd����b� Dl��F�p���#��,�r�˾���{H���dؽ�i�oCd�E�EO>���K�7i���q���0����bJzjp�?ϙ�������e�������l�,��[��_C������S��KՍ\�El��f���&�[K{��8��`M�l�Kt�P���|�ppP�iƤ���t쐜�Fq]�6���%�'�t�7lE�}@���4h��g�ymn�\>�7����^��[���CA�r�E{��?�f��=��;(9�ݛ���G�2���SWV٬[���A�;]%bJ�����D���7���|��u �-�,����}P��.\�Shd�M���}O��c���) k�g�^��G<U�5Y W�ff�\��v�YF���{����8�yK��b�+�0���g@p�r�b��٥���4QX�^�W�;�"��}F�6���'7����lG��
BM��U�D�c)?���6^-�Q�g:���VdqE.��s3�R(����>���L��e�j�M&�������qq1�I0 \(�Ȋ��+��C��"?��^����|K�+ٸ������0@3[p���/@ʠ�QEB����[��h}�
�h3�F�v�W�����_��N�eզ�(��t ��Z����J=KoL��:�?Mo��_�;|�H�������PW뎧�dF�co��(�ʜ?i?.Ϯ����-���L�����K���*a�E�Q0W��I�Hr�5*��4�q��+�|�;E����v%�PA	P�o��;�QUÍ+y߻XI�-t�͕�c���T�����_��o�M	���H�*	���2��&�'�Q�ҩ�H�l����9��pg�?��S��jv2��)2���I���ŇI��j��¸���dc��7f?��lk���Ѿ6;eT��*ʹ;I(�t�H��&G�I�/�HHx��@G�TF�m��_݉�i�"�M ��8l)s��g����X��[-.��Pz�.�P- ���7�x~��#�$qA2G��z�5�-���oH�3غ��������\|�r�}��֍5�e����Ϊ��o��}�A��N*�~T�����2V��؞pGPx�kGo���U1���HG�@��ą��$9�s��l~�W�$�8�e�
��K��`]g�4ɹj��C�"��u�*um;x�_��Z2��t�+��a�]��=�A�� �D$�0@sGX�r�5�9Q]�b�f
��tXOg����5��
*]����ҥ^M �������WOn�2kd�D�H�4ﲾ�T�34�3����n�7����L@��O{��F�[���T5kC��g�QpP�=�K�$��r̔�! �LJ���ŕGUL�~C�m,�#�:'���ؚ�=~U�Q.�]���Ѭc��M�b��Q.�i����ǍW�蝭fR�h�����T+xb�J�:�B�p�go^v�*�!��|���,� �ޔ*�!������6�a�u��o�V|��Dm ���	(��t�4�����]�I�-��Ri�pb�����h8�7��?�թ�����<w�%Xy��9]�f�YnpG��l�H/B,�h���^�,�@��)�텉t$2.aǣ
E���=�_���I��f;�?��2--X>M���q����E(�a�[O���Ѿ��p��Wĳ�^/�Q̹����WI��?O9������	�P��<Ф;�堠>�W7�U���a�Kza�)0�5t��ǻ4|A=5�S�Z�}c1߭�2M�QF��Dw/�}j�$�^��~�՞��4T���W�~���]n��u�Vm̀�rf�"��>9@�p�v9v�J��=`�U-d!ީ�Z��@��g/hM��h�ym}`��W!�@0��>A&��1+�i|�}FC�ń=����)�)M��[$��I��혃�հ�t*9D-�]���j��݀����O�wlU���+��x*CH`j�uU�W���CJ�f�<�O�C��*0*3LŦ+''pRZ\���2�;�y�������Qj}I�rs[�.aZ�u�6�ҚD@�4Jt�0$~TvP�M�>e��~;�¡��'�Fr�a�W��Z� ��(�TP�zY�{��q��[���" 6B���<�'�h~��6#���j	#>..�:'����<����;6�WE�ܯ�PP��|$ė�p[��@ou}����)�ֱ�V��8\IOk�6�/����K7�s�������{|�����aO"��@�:�O=M��q�� %K2��04D� �� Z
�h�1aB�aHÕ��U�y�ˤ.y����b�Ө�����;F2�@
G�.���M�}a
5{\��%��DNԼ,���&��M�
��+P�~���b�>�|b?9١��w�r�a[i���Jg:���}�hDF�v��2�v�Ttk��2/p���5����N'�RBv"�16,�r�e�2�W���U{uxnՒ�/���:I�ƉX��,$'��������Y�h��4�'�� ��?`��;U�?XI2n�@R�h}���I�;!J�_��r��B�P���ڡ���+�iQ��2nn�.6
��"�D�+�#z�x�I-SAP�<�2/��n�.�Uᅨ���q��Ij�$,���H�r�4���$z	�k��Nq	�"�T'��
�9p�z�����4�`)�w���B���^�7=@:g4�W8*���^�չ6��=pF�e�1ai��R�	M���B�溺����n�K��rs��=g�j�����j:��|]!Z�i�+�{U��זQz���ꀽ�0�Qz�sF��SAz�]Q���Wؐ7lnf���E�FA�$��yRӌ�J�#l^����6����Yc����cct��WIj
�,�WQ��K$D5��,�љ�B����,��9Ż�pm�>IF~R��ڏ�U�W�X�'���~7Ë4��`����X�2����qDzW�D*�G̳�&e�O� yR����=+m�����t��������5 |R�/#��
������ڿz���ț���q����;���Z|7�9&�J+���Fֹ�6!p��J��3���^|X]���Fv4yI����e �z�`h����JU��tX��G�By�oj�%,�{{Q�t9��AB�o	��\�ݥ�`�M*ά���t���%1hIjd���;$��q�0�q��3>-SUN�`�~��CP�L�=�8�)�Ū�)0-��İ��QZ)3�+O�r���~M%C,���/�p�"_|�&���OB����k�>��^жJ)�-��6dc�t�`Xcp�����$G����d�X�i
r̙���Sӝ�f[ O�g|h(���/f���zL�K3��c�X�zl6�~�/U2fN4k=D醿k��A߆�2/�ԃ�Tsh��x�ʹ 0"Q��R�	�x��*݂�Bl��у�V���Ӻ�	�sN����A;qz+	�ڠ����N�\D��	T�ld_&6%�U���[�)WE���bU�T��__�\ 4�U�!�h�3U�f�j8F(���G��������u��eX�~a�,I���ʹ-.L��B:,�̡�fU>EWp�15�ǭ��� �4��f`�p���Oy9�E�Y�JV1��m�)�;s���>߲k�'�mΒ7��u��? �^�6jGZ4�j�E��g�@�C�q��LW]#�0� �#ݱ�X.�S��[�����Hu��
Elv����>�pŒ�����uz���E	�i���0�q��(2f�4�ŷ�!�V��֠Fc<�O[
J�ʹ��{�yֺr"��D���Ի	�	��斩1ټ�]$R����
V,�@Y�����f#bz�^�QcXb7G?(Y������������F_4�XO�������r�:(�X\l�X�b<����|F��*��=W�8J����ڔ�]��Do�@�Ü9Y	E���J39ۆ���a���m���6SHv��>�,U_������[�ڼTq����p�B��b�e�e���ж($���111����U�D��
Y*���f�q�+���.��net0&���][$� �ɋ��E�8�y79���	3�+�~���5.c�]�"{)Z���td��k����1�n�@��j���%��I�R�fO||�!>f�vx;���<��ӔzWo��ҡ Y�nh���Q��vY��W���u1]adA����#R�|�Xޒ?r�L뛙&X����n��A[,����}Ej ��J��kㅲΥ��`�����ҴX��Q^��6�KLd�����D��m�:���%ŗ%�T��~��k�vf��]ZͥW�U���O�e:<s��j�\Ĕ)�#~��/E*YV���D[|��%C�B���$��2���=yW�;�E������~:��p<z,�C;�������=X��>�*ye��M 9������<җ��VN�U+5hr����q �a%�sWLTM*#�	�D����[�����c���w�olf�CPR�tMx��(�(Y+��{�>�r�>��>��<�P�f���"�X0T�Bm���F���x�8R�k���W�R�@�s<��/��Vs�G �mB��=�f��v���JA\][.UɎR|�At�\��,�}��2�	�cI�?�W��r�>����V��nfZ�aJ��T�}�=s���2��r کj̥�B�j-46�
������e*�:A����d�E��	s�� i��|���6LׂG�Ś�ⴛ�X;� �}L�Ρ� W7�������D-��	d����J�S�km��]܅D����UA�.�$EA���>���B�Y�v�/�JF�Ɛ�{�.=�I��O�i��6ڱ��nμ��;Wu-f�me�^e����G��n��;�f�m`��PA��l��F�m�9�i�z��`w�W񏧸dSY{�@���U�d>�,H��O�I��_���b���f�� �Yj����`�&ƪN�."�ju���j�T-�F.ɕ�*RDP3��,Oq��������`ⰱ�6y挗�=U�A23#��T��no���8�Hyܽ��p1وXK�l������ù:�fc K=p�2��p	d�P Uř7��S�jĚ��|��@u����-^���*~��Z���?5x)�(����@��� S@�v��u�!����f�іQ��m�\���*�7WJI~b �H�T}���J�G0%
�;[���z�?�l������"����9E'��M��B���~�����fԒ�
�I���ڽ�4�چ�s%���9*P�u�F��Z��ufR�~�f�lyէ;a_���Ⱥ�l&ё��/�<��Y��Q.����񙪦&����8�4D:M�ݗܺ�&+c3����@��ky���(�1f+�u?�m*u8�^Ⱥ �E���@/h�L�����I��*.oJ�����};�_����`�$�ퟡ`���X��C/��N�}XB2��d^Bx�����j4����KF~/_����@�)�<U6ťی/���TC�g�����E�4]2��쳏ĭ�Dl�le�?/���ښ2�L�JI�����˩L<�k�#�y�,�t�Bb%پ�x�q\E� ���J6�5�K���|���ȑ�2/�_4]����Vc	��@�;
���;�ˁ��H솁�ko)���A�v�@p�y�GI]m��e������%kx+2	��1�tlzJ�pŁ[Aܚ���Ȓo���Ĥs�W�w܈����#��I��X�����W�����o�na@$�K=9�@�WX�V�� ��� �a?��? �25<���b���H?36 m'�A4T�Y#��
]�ؕܗ|�O��V���t1-��}��s:r1��Q�W�F�Y	գ"���j�c/���ʪ$�����<�'��0�P�H�S���q�{�!nx��<}\J�{��NqAR]sd
1�\�l�䄧�ZW���^���x��3�9O�x������d�}9�̤��� �u�	sz��[B�7��!��

�=ۙ��p�=-��_y�U �V��	�ƒL'
Ni�i�)X<��F%�k�3g��g�[1�a�9�i{t��M�#i��(�&����;��k'�t��p��v�  �@�Es��g��_���{��������y��L2�ϸw
���5�C��07�Ꭴޮ��}�2CJ�h�0~����������|4N��ղNr�G�s?/	;�t!�=yA]A��Ӈb���\�B�
��w�ɥ����5�%���H�J4����4���C]3�g֨K&�WUht%Y��?Wg� �<�?h����s��z�� ��I�GgHFHm�aζ[8��"��������p'��-9�<*��^�D�*j��k|D�KR�+5k�<�iv��bZ�zϠ�϶���[ە�-@u�/d�f�� x"t��'���،��<8JG8w����kv�f���8�-�I%��g݃���������Ԯ���ʷgĈd��y@���22R��[^vd��r��D(oʴ����!u�%��&;?�G�,��F��F`in��)p%���O&�2 �@�?p!ˀx4��+O�5���tQ�q`�&=:��OK���|*��j���*�N��\/�c��c�;�0��{�����`��uvqrVQ�4�I{j���<��M�qm�����[����cCt�R�O��Ꮣ��g4mO�����������.����
�c��a�����ҧxhњ���81�����_�2�2�e��Oӊm��h���G�J15!
�h��m2Eg3�s�[�T�IU�m��]�RE����O�;��V�?���+}V� /�:������1O,�4�C7���x�lJ�Ҏ����Ԭ�J��FF�����-L�'�ҿ*ӐKQB�{�� �<����к����7�B�^
�T�}��喷����6�L.BM��ۆ����SA �a���E�wj�{L�,�pX�M�g���6L�������ZK�U��ug� 6?��)���/��G�Y�-�9���0=Jb��8ޅ�O\&^S��w�>�50�qب�'j-R�W�)��| �|�
U)��l����^���E�˒i&
|��Ҥ�ߺ�*4�uy��Se���+ya�㡋�ס�f�?5���d��|g�G[��~�����0n]qZys��D�}ז��g��vw����LE�Sm���=l�#/ˠ�S�YO��nu���n��N�I���o:���< /�+d�#L/��e�Zz
SŬ$ޫ�Q�ÿm�2�Ro./� O������ʭ�<�33�q��c��ƪ�����<�%������s,�T��l�I$W"�(��mP�.�~�U��*g���Dɺ.��Z��9o�h��^�	��x���X�ˢ)S�~�G+�<߲>��DN���kp7�4x~����[Q�ƣ�A�c��A%��_�5��O�x��O�3%��$;�*��T�v�&���ki�go�u�f˚�ʕ��0���U!n��@Y(���^�aB���3i�U�_M4�$��������<*�֣��E�<��]���>����>6a>��6o��w�������;����}-�7ZR.�`
䡮�s�(��C�D4�33f��b���yG��.�9��i5�Kr��4���oL��|�9#�5_#{�qg�߇"5�m���rU'����N���IB�Ը��_��tk9靏��rQ��䊨w׍A�p���%q�C:�Q�a~�P�5�~	��ԕ?ݢ���2�T���� ���M���q��ko���Wqĝ0gl]�D���(�D�@�н����9��[8>�-3HcM'w�녿�B��X S���>�k����n$�xne������Ҳ�Z^�K��}8��U���Պ�@�z�1�Fj�R�(�{���Y��p���<D�>e�:Y���r a^�Ű�8':�3l���y��L(�.�6J��4��	v9V����㎧���j9`٠�ܟH��j��f�Z�(>dNy�4���)f����oq��l����m��mɜ�Ah^�t�����F���A�����'��2�G �G�n�XK��I�9��!d;�"�w&�68��H�W��M�hFkb����ܿY�\/��"��}9����>��;Mh[Z� ���F�,
�e��9��ȋ���&�m\I<��յO{Mõ/�eo
ԈHer"PK��wGڦ��W�ջ�,9�2i!��	��5ҕ}�%E�B�\�Kቯ.p�:,��s��:U����ձ���6�sR����V���.�&Z�m���8���H��Rӽ�%n$��/�x� �Ή�3q� ���Z��t|���"N�K(ڱ\@��)������Zl���x~�9��ϣ���i;^Ag�gV�9�y�#p�6��<�j	��h��ǯB$�.mI@bU�S�����j�ex��ׄCX�5�#�Q�*!��d�hm9:/�8~�]{�KUқ����D"]���Q�Y�dN�M����� L�ϗ0;�hu�]�C�^��HH8g�F^!�|/�:.]���YKzN��`{tk�<��J3^�O=�Z��A�|�9�:�tKȝZ�/4�E�U��tUcfXk�C�+QR�y�F^��)�I(���;!���k����[3*��&���'eO�*oo��o��+ �>i��Tk��W˜)� ��A����V����Yduݏ�'P��\�ab��t/� �-3Xmȯ��>t��G�L>��(\�y9�iG���b�|4 �yW��_}	���{vd�My�K�ƃ���� &�s]�"�<�av	2q�jƽ�6�!$����X�2c�*�+՚>�CUuX�vJ�Ʉ��k�)Ǹ;���@��mzT?��T>�5�ŵ�OG�7�s�����)�\���� ��-͊"t;΢��p���ⵍB�F�Щ�Ϸ��:ʮj"l�Ń�ȃ���2�H���R7/���kh{EL�X�;���/}�+��=���1]8�JFEW�MQ�&����o����N��Y>��wWh���O>�O�y��-�{��27g������K��z'cB�F�&��f�:1}OF#5����u�k��#�m^���V.K�}Z_����vL�,Z%���: ��B�p�J'+֦怷X���jCol~b���R�}�����:2��0�~Z��{K(��ם���2P�\�+�]|�zQ�.����,kRu�!���U� ��׸��&b8jMڨ�젳4����j:%�\"�Y$�<;b׮�7�O�ku��ق��#���{�4�帻����O� E����g��<�+OyL G� ��Z��<N��ɞLP$䤠�3=�T��m�}�B�/~S�h9O��nj�4S<���1�y��_�(v�~�/'Ղ�H��J�4�0r�'�d��xgQ��#}�s�������c���Q//���������Br�T#¥t�N�hb?������S�K�}Ul}/�1U�)�nrr ��#f���÷���}�u���4�o��������U;)HFW�5W��<�3g6Fhq�w�\�at]��l��/�K���|���r�Z5jy��0�k$6�a��ft�K�9&<�sec8��L,�S=td�T!-ÉpS�S�/ߙ_��>S�Ҳ�ŭgh`�w�by�s�aR)���J��U2깇b곮0���c*#q�f�Y4���Y��~?������#�����Ցeb�Fv�$,pI�쁱��L��_��$PD��H���a��$�K�gH"���P'�.!�;.�cqS���cㄟf����9Q�\;��f�[9�A{�"�/�� ���K�[0�֚	�J��nm���ŷ��Æ�ͯ��d�W��ťq�J;�<9�p%3٢͖�@ܤ?�V�ב5�Թ�bL7���|�ӽӢ�`���?�1�v2��Q�y*��,�k��xOP��%�gN�b$JD�H"�Z�[ʹ�����R}����x�]� ,�IFcA��i�y�d�d��5r�z����ؤ��0�(�V9���[�8'V��#�T �U+�F�3%�5/��5������"%�ة���ty����4b�Ѱ�GY�|V��djR˘���D�l$�-�����O���s�'����PV�
yA�FG ���ӯōK��VPT	
�S��c-s6䷓H�x�+Z&�h��0%H}$�X�;ށ-3��0��@Fu�#
����6�F� ګ�n
{)н�(�5A���!������{:3��񜐕�� G&z@�p��LU���v�����&D,�΋\����y�o{ڨο�ڔW�YT��J]�]�`.,Y���=��[�zɏ�=��5.�ٝ������'N��Q�H�'�r�%�DZ�Φ��0�apdx+o-g�O�l�f>NGjtu�>ǘLf��	D]��o�nf� ���YЪ��κ���P��-0Ƞ���3������%����4$x1�$sVy��/=�F~��M������N�0}����)Юa?M��M�2!�}�]��m�c	�3h
�|��u�p"�-�췺{�IƦ��E���_�>�q�efT�S�,�Aӥ ���8��ͳ��1������U�c��z�&��"�$�"y8��X��D�^��$
=��{ʱ�,���O�Ya��������t�];T�~IW7�ԛ��+ �H<!�����2�_N=~c���T�an+*ee!�f�~�iǂ-龫��N��+M-���YJAm������s�.�ciO�(t+���MY1��˅�S�&e��$Mݐ��ƶ�[�S�I&N<�g��C^۳�J& �C��D���}&�p"����Ô�_�)��O�1m{���Xp��e��Դ�<��M��&'_�@�r���z���7�U�,F"�P�Bt_��ѻp��"�}ls�b	�+|���-Rћ�o{��1`��V�Yu$}��Dȹ�Z@���<t����Ĉ@����`kD{�!2��Ċy�D��9�8/ 8'�#�V��EU<�9݃:�L<��oe�P�٥S�w��7��js��5�!NpDVK캆>_�Ș�/�'���,��Ip�Ӊr���B@���K.�|���Pb�������q$�����TF*���PV��ʑ���=hb�5m�0V�)���QKM*]�K�`��>���>����{����]ڦhF�Dլ����y��0�{��1d~XU� C�{����GA�
�EFIh����	�U[\��M�	م�p�T{�+-Q��y�Ҝ�'!(}=���9�gx�=��blw�Rm�Ri�*hc4$�7���t���@��X��f��6�&@d��F�������:a0��nVŠ�����RbE^2 ��c���I�5u#1$�ޟ.|����Ϲ=�_bf�����
��qq���i���0�y����8��<A������w�w0&��@�����%�40�qw�&�ӓ�Vüy��v;��Tb�{K-Hg�_
O�����5����j0�'m.�Tc��S;g�QL���^gAÿ�\�ܧ��q�& �pWa���-by���Pb9	9R�z����y�5��`���g�9ڀ�Q�eS�{�M���d)���Wv�KZ����jC��7����W:�w�Bs���G�܉	�iAa"wW�z^R;��ؙQ��gۍ�������i5��ؓ����6�Ѕ�B!f�(y�1#���1�9���ܜ%�4橳��}0A�fGlU0m7^�o���;�UP{a@h��[�w�wQ�u.������F|�X�)����}?c�A�#�8���(���+x�l�����>�޵^#�J")�@3��*V^|��,��N郞�D4���]̂@gw���7(}=�#�>����Ge��[��DHl�o�f��\���<X��6x+ �z�%��/WM�1�,/ +�o%��-s��GRy�X���,�Z���O��[M�?�+�G�t��$��Ԍq����hXF��t�c���iƆ�u�}�l�Jw8 ;�T�LLBZM�Ҍ�dJ�=��kzV�nAXy�b9B��|tpĴ��$O-vԸ�/L����Iͳ��%�eK3}�w����A�N�{��Cf��	�V+:���!�r[/AZɁu"(��5���l�sY#������5#��,��������)�oC�`��~�m�7E}gH蔏n�J[cϚ�'䉪R�4【�Q�!�ӽ����ڨ>.�u�E+b�9�<�i��g�
O1rGF�BS�|w-�Eq�->D�aK+Y�vR)n���^����D�xx��w�<\��v��J�b��\y&�PS�'�pLo�h�(�q�x����)ɑ�Ef�3������O�v��H�����}]sJ�Eq��5����D�]�A�4���bK5t�1�v�fM��9��"��K%_��A�;a;6P�Io����6���3�آ�H�
֘=��3�݅�@b3�ѵ��#b������LB�C�^��#WOL��r���cLNe�Z��x��:ϟ�&,��;�!�u����Xh�䃾v`K���Y�
�"�n�|/?j��8Zq�4��ƍ�벆~�SIj�@	DL��0`}�elFcv
 �RILm8�`A��IU?P��w�
�Sߧӌ�1�b���{��|�F�l-���3�`wu�Pc�B��P��`��ǂ�(ߏ�&'��"65	,��p����~˟f�[Y�#V��+ev�?v��F(�u�sM���L�,=$�A�~��j$��&�+w/+s@և(6ٻ���<F:6�L���B91��A�O�a���q��o蹮�f��L�|���]U�����9�����I]B��a|�-A�Ʈ]��T�<5ߵ������l��{-����cj���F�	on+��<���E��@�/��Q��Q�N��N�of���z��d�lB?Z:4#��(.�Y���-ud��_���ZJ������Z�?���rH�Qhe|�d�k��t�U�Gla�gk�X���gd����~d�M�[ n�^�� �n1h
T�L��DJ/ ����8+� ��۹i��%�\��{篂&X:�4�nӸ��,�4�j��H��#q��=z'� ~�371��7+��������
�(F��B����W�ߴxȓ����!��$��ש�{��[�� Ƭ�o�va�8*_��n���!;��	���F?���Ȁ�:��R��ɽ��zock�����hOt��y���Z�<V=k��!?I��t\�������B��W����F�+�%��EC�� ah!�)N���M"�E�^p��qi� I�zޟq�C�c�w�U�\E�^��J�ͱ��� ��=!�g��Ϧ
��sn�.��B.K���|t&�{k�g< �ޗ<�b���-�-��s���4R�ȩEܤ���ʮ�>����9f�V�i<�}�ؕk5jWn(�
�X��Əm����C�BǪ��A�$r8T\�� ���`ݵl��9,�h@v�cq��ժ"�o� ӎQ�d�X2�	5?J�_���ؾ�X.0W"�2��ͷ��0��J�W>e=�B^���0����WE�^�;f1v�r(�j}(��$���`g)E��5 q^��[�-�]�O�?�9D�>�h0�E%V����ސ;�ĥ&��IM�Q�H }�w:�E��d[�B�8��D�Cf��.,u�Z@KG�<��|�!� ?��d]]�+������5i�U��f���z�&:~�f�@�6ˢ �1/P�������0�=���Ղ���@���MQ~����6��
�N T ���=�InL�|t��17��e@�JtaO�z�����WwLq�1FAf�Ƶ)�۷���X�h��TS���5JI�/�}g����m�MB��j�]U�m �8��U��d�_�p����z!? X^.:?�X4�}��B����\�/��!���ܐ�X3���}�"~o�khm�%��ɥ��NCN4�Swe�%���=�on��V��u�� �jǻx�g���l�*	ь���<xf��e�]��:j�U����g�y�_`Ƴ����F��7��d�&&�4�����*;N���0�M��&�Zv����x�i/�r���!Y�iI��v��0�[35S�Y?c�(�n;=�k�]9n��y���n�Ҥ"�7��HKdȧ+aQ�G��C��E�iN���Yݴ�"oA(��7ǫ������T��&��n��#�j
8�R�b���ʮ�a��Z~�ǉ�~���ÒьO:��	{N��}	��vX�:N���4�嗔���X�p.
)�m��(����ꚗb�5�#�X��+z��}�>D2��q�pEr̬F擜
&L���mS�z�d�*d��.�c{�^&��e�z�^	15������b��r��R�w_Y�*Xi4ǝ�}4 �4:ph�sea9�w'`���n��@/ި{�=ɼG),Z6G��������^깕� �`�ܸSAt_C$
�y��{j�u����x���+��A���f��8D�MV�l�:XGE)���*8px�k���(��ݘ&�]F7l(��5��%n��i[���I����9l��B~����d�Fu�l�&|q@���"��W�����?�Z�C��\���Oy-����Ev��GaԞvH��l942�fnEp�|
�x��� *p��8���:�tY�1Iumfh�`a4�Q&^����];|��o�S�~c�j�2�&jwٞ�#e����^4Q��7wG�g� �����_Tآ��3�9*��x
Ԛ��O����sᔌ���Uհ+m�ي���U�Q�%O����4�q�4k!�:N�;�l�������Y���`.'S�sȃ�В��eL�:�+22�C�tx׸ �K���.��p���[���>��9$�H�Ci#:�␀On�Ta�'�	��:掍xw,e�e]�X�#B4
@G�'�Z�&=$֑���{S}���=�o��,�";?�k{�Y~� -~��f�+>Av&Ј��9�a����ܑ1� �>�#���}�9O#T譌�!V�����w�$���/�|x��g��*�������L%xp){ڷ؊k�H����&7�e�(y\k�(�TC�Q�?��0�Ex_�)��&��:��.�&��:�ly]����	~иa �l돃���N	������M\��Q>������w,B��u:����-'4]e�lt�83�ܱ3v3��ʫ�{N�n�93'��k7��P��'�.y�6��ؗ�{|��A�<F�����@��r3�r��1y�X,���9}���n
�$����[�?�WJbğ�סf�)�0��l#�Jia{����!��˖Р-W���vsw]s�����~d]I��-����9�}�R��?�-��.�m�g���@�Ү�P3�f,�|
�j�oq�2�b�ׁ�*�JG�����H�ZU�K�q�,4���:��,���h��W��cn����ݮ@b�g�~�h�������AǍ�M}C.�E˃Iu��ůW�C����V�۟u��x��Htw��{S��ߠ���`(��.�`���{���)4	������2`~�Ơۑ���M_��4�$�<Ϲw�+�qK�%+�I��MP�wOK�Z�!0սh�`��NψaU�)�� �*̹"d>]yN�J ���U�ι��j�����	ȃ^�&4&:Hz1��K `d�$M�?JUx��Ԣ���|����@��~}V@՘ԥR����C�k�΀L:"���4�,�U���gfH�x�d'E�`Kc������]`;����2��qк���=�)��.��g�� q��o��o}z�XXL���v��F�K��+��� ��V��jڔZ3F:�1�5�����E��H�t[r�z�Ռ�A'�д9��TZ�j��x��L��˻*p�y�.�]��l�<Ļ0_]vn�.��9��ɀ�
�-F�����OƏs�{�aٔ0}VbO�7�di]��t~�ع���eO���IєK�@��z�N�m�y�W�!I�`f�����͝�#l�;���������] ��;�9��� B�;���kSe�cj>L�;�D��o��6g��b���&�|peE�pT��8�M`]z��F�I�t��;��ˏ�}*��d:���G�pz0��Wg��4��!��ܤ�x�N�~��q7]�.�_���p��j�'���73M�$ ���W�ۺ�	���*�񳜽 ���n�Ӝ}0a9�\��mw���K%�Ae���n.�#�Ü�9���Z�8�L4�]�4G�W���ª�K-�'��h䶃�<ẵ8��9�i	r;0"�H�냏���h��C��`�ƽ���s�)a/!	�_"ZIt�1�O%KI�������9��d5�֟5��L|�9���Uk@׿��)������31'G��Y?=ӿeX[L�+���^r�c�t���ndҥ�E,	�k[Ȭ���M_����GzAe@�d_�0�Xp��Rn��;�~;2����9��c�
X�d�}J[����;QU�[�:��$�e8ƇGY��jW�M]���
�5�ֱoU�c�6Hÿ����B	�5O44���-&>��n�8������,s*�YG>h8Wvd�!��[�}�!�&mQ%!��'e���Op�Ac�`�͐�#Q�[�v�v�=�D����J|��
T���bۤ��o?!����N7z1wvH��!W�Vɤk�{cb�Q��5��}?����]0�L�Z0�%he�z<�#����0���#+�`�v��'�8<E��n���k[���2����K�8��FFR�/{$X������w %:���U��r���]�y��&#��؝J=Y�\$���Д|N_�b��F�.��%'{)�B̘��ig�-�f��x�����l$�]�A8��D�Q�04�O�C���P���Z�C�-�|;PU�.�(��hu괤7��� �cI�1���0Ik��mW��?2��&	���=U���k�f�e���mL����TRڈ�ћѢ��M� �n���؇VڶwGP�|���`ǈ�B���Y{�=��rx\+�p-���m���Ӏ��(mདྷe�F&I0U��a �~�Ü0��g6��~*��j�61���En���P9��n�k�T�������G9]F��U� �Z�*OC��n���D�!b�:��~9�:���e��p���4(\}^q��6L�$�,T����,p�C���U�4��U�� �㤎k5�l��w�� ں��)���OU)�,Υ��+����|1WR6���0�)d��B'��p�	M�,��$��#{�f��[��Oe�i�{5�vJ��`��q�a���`^/i���D*�cs�U��5[bs�]0����E�
X�on'OG2-�2U�y�F_7|��B�;I���V��I����
MG{����eGqٰ��n��&^m��֣&�k����*�/ZD�QH�:,���!�@eh@C��c��ƲBƧ%�����7ӑ�X�|~۴� h�Gn}�Y��`����f
O��Ot�\�]ώ��}�����,�ψY�_�J�|��Ss&q���}�Z��>O����9N�L� ��Y:2WU��lkg����q$�)��n�0�{|J�,�>r�ܷ��p����cF�Fh��b����.g}~�0�=anF��(�X<�����E �8Y�<��E��$����!Y�.u$��$���o����D�x�����b���)����7��8��ӟaFd�F�P:��3��|�%&�Ɠ����v� Mz�R��\����a�j�ϱ���"�{�#E)��3n�YȈZo����M 
���`;A�)"�V�1!�\��Q~�tH��mifz������*��!�����K4�����������:�M�e=���O��7u�fS�G�8��j<�w��rC�Wd�����v(˔��B�K��}� 璴�
8��7=)֕��଎A[���כ��H���O��R�K&ʉ�C?���7%���,O���؉
�f�(����I�(��\*7�US��v�-���12���h�0��7[��\1�t�N����;3*e�Ȣ�<�����p\�bcC,�HsnҮB��YjJ�����C�5�tvCMO�E=R!AFx��}*ҳ����Еt��R���E��i$�qa�ll�4V{���;kiV�o5r/�a�S���E�
�&%N~[��Q�xj�'I����y��s�����]����|A��w��a�i�]dq���M�i��m?5�kJſ���*V�R��.V�:i�)LS��6�t�T&͕�
�x:��r���xgO�1���I��8���h�С��
@����K�E�`f�)��ր\1�E�*_;v�w3􇠩11��;���2�������Ɛ'�7�W��#Ӄ�����Yz�͉��(�/����x��R��JD�:ɢ�]�,kB^c���:ǎ�>B��L<�Mi�*x�^������1��*X��c*��	��	����8���l�6�J��b�K���<�?A)gk��P⯼w�aD����>&&l�˵���v]o��?��l�3J���^���ky�G3Z�P���\���Mʨ���v�l�k��6U=q/7"�gkd�;L��S��B0�1�=ޯ�,��%�P�@��(n�Q �2���"�ndIcw`�-�&�R��^��� ����g$J]r�U�6޲���T(�Bݣ�2�O&��A�'H���:����ț4�)e�?}R�Ģ�����(X��T�o�x�U���kl8B1_��߃��\J�Ձ�`'�;;�G�u�:z%����N��;� ����!��Y���b�3���r�:���Sp@�\��KY���٠*��S�R)�8����YKJ�?U�>0����`j������ؙI:7"��+�(>*<������,�i�y�_��5 W*��R$�Y�]:�m�]i��F�,�`fF[r7.tG�M�"��Nc'�6{'^�찭e��%:���*�n� 	�nN8;����"B��u͜z&葦�\;��H�`y�C��|�t�3�b��LuNTV�ݢ���nFErw�5��e�<i�);&"
�M�(�lҷ��{���C�M�a�}�L6���59�V�X���D�9������1r��bq����^oY�#d����@�T�R;����Ԋ1bah� ?����N�|�Sڲҏ9�I_��R�-�H��!�|�i���������;g1)�UK���w^ޑ�_�mrz{ń��0��g�h7#�BHn��&$�.M�2'��K��2!������;��Q���Z��9�!tb�"hm}�~�����=��h��}�&]����Z`���p�ݙ�������k����OU�,>e泄a����uN�����|�����Q86$���+s����̛��y��X(��jБ�j�o�����l��PN�r���_Kh%���Y�<���;C���D�,��3��\��7��$����
��y�8 (�ꜷ�(��G]�:ײ�dL�C0�ۧ_���"�Tq�JpNh���W�l�h���Pc�֖�I�}���f F�\�km\�z�V�m�M�yz�;��W�B`���џND;ߒ�:�{eE��E�<�5�Yˁ��	��x2v�B���b�pe܋X�~��a�������j�J��_���iW$FloO:9�d.�/�N�?}�֬FL���dzI�+'�ɯ�e-�Ql���>	��"�����ޅ���_�"��6}�/���e�>�6z�׶��f�:�<'�����[��P�G�#<b� ��pT����AP'����h��N�|���W)g{�)&JM*ϡ��	&o[&�cܯ�7�Uf�VI�̧�xmub���?��d�<������S�<�-g���q�ԕ���irFڠ?s^�-��4i�æ��j��qTH]`dj&�2⃀�����h�/��^�;&�Z���Is�����~��p���t��خ�������>���A6k��rה��먮'��g�&/,P�A� �#�������f���*?t}(����XNB9	.��Q���TJƁ��H���n;�h��h�#�neJ��Kǣ,w�<?*.����KF��,8)鶜4����2��?���D~�"[����)�N�v����Յ\a���NgJ�`@R"��x(,i�E�A �Av߽�s��h��X'1.X�W�ë7.D����!1f�f������7�w���	�}����_���&H����0�>�*0�s *�񩲹w:.�i��a���,��w�\^ss9F|P�W[ϣ�L`>����m�OmD�������'�P�F����-7?XD|F�g����}��3�M��� !��	%��>�	
��L���������Z�&t$�5�^'�*d��;"��Q��۠���$M7�N�{�LM2Lt/�t���Ŀ>���L�_�)5pk�A67�P ��4C�ZL��d��
a�gm�z�N�����f��bD�/�H�?62]u������Ʃ_���ӓF5�����Z��Ԗ���p��Bc~R%&SH����&(�C�����wB�պT@�BnH��7��l�0���k`<�{ң������r��S�ħ�&��#`��f"�J��!R�:��/�"W�|��Ɩ����ъ�
�5r�Y'7k�j��n��P��n�aBKR@�C\.Px�Y�5����R���c��uS�+|c^�BUy?��dQ3�8�� Mn��v�t��.->��Q���23b�����X��lY5ղ����kb��q=e�cR��žؗ�� ;l�=��v������R�}�f0�K���1���y�����3d��_9>l‗�`S{8��شW���ΉUߛ��H�̤[���ә��I?�D��V~۾qH���oi�ɝ�vTfO�i��(a^;QyL.�����M��0UG��gtk��|��qj����V�)���|�?�n��uR�8���? ��^!��Aqn�H�-�<���zUMs��F��|xW�%�!�ck���4'�N�=V ���y�D��o�v��9�KZ�g�o�8м������e@���=�>w'�	��U#^�ү�J�&�y v 9�9[�P�J���S߄�!���|=q	U��*�ճ��H�e�<�9�ۖ:�9�^R�"Ϩv(_%A�K���BD��B#��x#'�o���㘼:m�$�Bި��v�C�.<Ȥ.��!�RY�2l[J�	�Q���D��;��y�����&�w~8[����#��8[ɯO~w�8՝����,�{JΞ��± �L�4a���TQ�cW��_�to	�_����M�L,u�����nW�� �dZm��)��)%[e���ץ���já0!���l�FW]d�Ңr'�������2;�����g�ZA����y�6;�K�3��4�o>�B
_ȭ������	Ü=N��w|S^�^{L�Gc�BY�B�.�i!.>�%zEH�]��+{P>�W8NL3�.�V`�DEIS�#.l����B\�k0�������//�<����3�8E'����Y�S%�����:���y\:	�.���*g��G���~�B�'Q·���`��1�ƉڛYT��[�臉8������W�Ά녚!������ք����p�*>`��o�c3�i��՘Aaq�u�H���5��~�%d�2 2�h�vT��q)�U�v����f������� @�]ҋ����Ը�9�|�k��N'M�3�Ǻ��c}4t��G��i�㤓?��aO�����Q乬�:�J���|~m�#ӥ�@���}	SF��,(#�>�HA�3,�����OV!����-�x�c�
ۡ&8O�O�hj.�"~��M�v�}?z�*<�BA-"�s�7XM�������0�u��4,���O�6h��h��[W\S��hE��S��q^�@i��t4���َCm�E	O�;�t���*Y*v������('��X�����л'u�d2�>�����r��D��Inu�n٪ߩ�h��|��De#����5	FiF��h�kڰ���4>�Ļ���oRx�7���+Eu����F�
7��΄���xGH#.�'Vלk�2�r�$�n���E ��@�F�O��'��h�j��*CP]%��m�'���`�"�?>�/J���+���c��z\#H�?OU�2=9���A��`�����/1�`��x�Oj�P�?��A,� ��]�G�T�����g�B8NO�L�X�zg��(Q)[N�M������F�N�2۫m�0}�^6����8 TZ�>��M�JYJcd��]��ur���sK��R][V���4y`�P1�{'�j8�����pP��Z��)Ƥ�~/���+�pV碕�ΛԷ���2h��s���⩤�:rq�<��Dw0��d��N������.�����-�3Q35��7�S�;��Al�WN50S,u:[�~;�����Z|bn���ZW�P��-zZ�M�<�;0���w~��%����)��D�a5Od���=F��h(�31�7Gu,9�R�i�nm�*�{<|�3��5Xn	�Bǅ�Y�5�[��q�����C�,�_�����9sĔO�Ge�<'���8�IX�]�JH���!~�L�f��G��V�q��x�g���i��S���䦦�|(Jt>b�4��V��2H�����=��y�E���ֲ���`4�fpÖ�
`>�.��qK�h��?i����T�h�1p��BH@Zw��}b@�|Ū�
���X�d�'D��{���=]~j�䕖זţos<����D�`��Cug�TR�N��JhK���:vM��q�"kܑǟz�sҸf3rj5�v"���D7���ՠp+���:<v�O��%>]д[n��14�*��^!Qi��)낈�_�?�\0�VGo(HWZ������S�^�b������V�_}Oc�~9U|/�Kd#(���O�W5F��z��a��$BL���΢�%YZ�a_DtG�+�{uS���w
�Ϸ�q<�QHBی1eN2W�t�ncˣ���h]��2��x�6��?N�Ͱ��wt)(ֹG�&g�͈��D�>%#�
;�����<�&=C���R���2�t�;@U
��[RNvu���_����
��A�ҖK�~�ϖ.$�9?hLՋ�`F��^�Qpڨ^1j�D�_��N�k}E� �������^��<]W4���v��6��&8*����F,�#��E~֭$�(��]C=�mvUR9�Y�p[s(��%^ej`�R�$�NF[D�e�uޟ�y��hɁ���o�i�C���$0�����w�3:F����b�r��s�W��Z��Lׅ(���}��~�u��S�U�c
���h�{��=�j�Qy⎣ԛ�تEw�R������v_l>�#�6�x�>�	�!$V;�,�WF�g��8
G�W��������[?����ȉ$Dn̜�&��U!��4u��'��c�"������@��q��8�D~��l<�3p�N+#�"��O����� /��Z}�XL�Ӫ�xG
���倂|�6�L�^�87�c:�R>�&z�,��
f�@�ƾ�#��1������h�}��*M�t���\�g칼o��|�R����M��| �JPt��[�Rl�����Ȑk�!��E��s�X���,�mÐQ�ދfVjZa��2�:����څ�T%^�9��c;��_>�4!j�;���@�P�v������I*ZxP6 y��D�}<Q��P�[C u�Ѭk�e�05\ȇ��\kq����n��u��Kѣ0��a��p��}~l��� �|�A�e�,�e�Lb3�9|:k2��V��2N�T��7#���٭��y��eP��im�)�W@r$�Z��]b͓�����h�x�� �Zz6)l0"��R�J��G�wD�=B�͇���4=��9\{��]yvަ��Z���\#�d*���X��Q�Cۧ�+Ӛ���9UH
��FX�⡬���"5���#O�Q{"��TIe�Y�g�M��
3ĵ������K��!��a�5�{���P���,��RFg���џȰ��1�rZ� �!��<�F�>^�"�����������@/&��r��̺���/H�h\�l�CC?x\V�p�օ���)��|�\6��m]���"���rԄ��Џ�I1����)�~�D��\�����0�-�S������3���(�����`�Ukuم'�<�`���6�`�Ht[6��žc��m��������u��C�:4�me�B'�kOZ��LF�Џ��XG�c$P'�C�&\��%EiD�P͈P�r�����������V�p�$ޱ�y�����kr��;�K%6���WKV�Ͳ���P���Wq��j�Q���	���	����Y�u֞ǭ@b���7����:y�#�*�Iӷ���y��<�4�B�s2,��^4R�F����K)y�e3 ����Mj��0�U�TQ��`ih:�嬌'D��"�����jf֠#i_�	?�|��93�ꄘ�2B�jO���J��Wr�uA	C_s�c�VN@��mjr.&,��+�{�0ΠӸ	Dݙ�Z�*(/�c$X>����K��J"���ޘ� f���݂1SPC��ܻ�!E-v�FێB��cc
�o"<�@�kU�=$�Q�M7����Ɓ��E� �ހ]H��|0�R���e�sk� ������4�I�d���i�X���p8�J��yܣ�s�vz�z��#�ٰ�s���Gg�Dǡ���$%F���@m�0ģ��0�kNkk�jf��0� �nxh��Z�>�}����å�e�@��	��͍SZʢOl�{�Q��)L#i��[ĺ�E�H�aj��\M��g7z��>(�;���0ۢ�,���L��0f�;�~�{�r�?�*���Y��қ�Q�S}@&CA��Z���S�O�N'}�$�0���=�f�Z} �7b���)���������g��2B'qTkdn�k�n�	U��g*��n����;gz�:s!�c*L���I���7+�*�a精#�gt##���� r���f�d��^� ����K��!&]�?	b��PF����z�\D~߮i�8X�����vE`F�\���E���g��rih���G�E^ ��,y_��n
і��Ic�Q�&�k�R�v��9s~k�ߎ�S����>��SN4�ki��JO�C}�Z�j�y��"\Fܼ;�P�x�ܑ�� �WAS�I�m������`�������c �)���w����rX#���L8���ѽ�Bj�%X��2��=����ELFҮ T^��3��t?��ٰc�Ta��1�S�B@��e6珘q	Op2�2̨���ָGTD�a-1�`���(*�(�������;�vL�<Z;�M"���X���Ht��՞�ɸ������Vj0�ub��ě�ƴ��7h��~ԂE|��Z��	>^?>���u`�lgq����^�J������m��K���b\E*W��K�Q��֑��D-'=�2����S�}!?����0'g.�h�^eyz�H5�r7��	�b���z��G?zМ����m�.~�:Ȭ
D�E��`%�\f��޽V�{�������xt�~B	�wm��rČѝ0�`.c=Z�.��]�'�<Ӂ���'�o+�.m�w �ܜ�Γ�?�
Qχ�FWkbȅn~o�r9�k�	����_xU&^6t� �& ��Q�q�-5k��9ΎDN�G���}Pq���3(P�R��s�˘>��L��=˭ǿ%�:R�;R�%�h>�R�w��=�Bk3�κ{�I��ÿ��|�/>NA��3���{k�L����4[����8���V��C��^� ��N+��3l������������*
!y�t�����l.� I�2YE`-�Y��*�'�f�8�-���ꓞ<c,Z �C�1�u)`F��G��X�?h�I��ܖ�^����.�3ùrv��x�Ӆ�W)�GU�u����@�h��Ae9��Q}�!�0O�x�l|L'��K�8�M9�����e������}S�ɂI�f��]�<iD}W���8!e��I�v,���)Qb�:]=Z3�'��8�Fe�l�Y���>��DS{|_^���c�����`mb#���u{��`ռ�cĴ(�$0���y�v�NksN2�gV"����dB�	�Fh�.u��7��Il������5ē���;+��牦���\�-���y\�`X$�ާN����l�f3As�L�O�V	�ro� o�ob_mNk�v��Q�����_5aۻ��^6��mM�*o�q��3J�|����o_�H)����sa��*���8/4�@��+��{h�9����as���Ӟ��*o@ԃ�9�<�@=}�7���u�?h���d'��$�*v��3��ϡ��hL���۬W��Ȏ�x�X�i����D���]^�����*�y��̷ͯi�<�^m+�C��1�OFb���n��m��ܘO}��_����l�I���~�
�J����hA���||�HV���a���ARǕV�fr[�_%��|(��
�+"�e��0�t�i�oP9#d��jDO&-�[� �v�z>z�6��w-��(�jK��H�?��٬l�V��a��g�z��2���>aUOI֊Fԉ��9'�~���!W\�"�%F8&wF��+�Vu��u�z4�{g.w��!��g}��x�	���>���?��g#����>�����c"n~�i�/md����x���y+Ԩy�ŋ�\%�`���K�����3�c�q���;܃��]|��~L�T%�ޛ�
��</5V������'B��Ec;	��F_a�\dLx���h�d�����IH�
�1aYj!k�$^q ��h��}����8�r�@+�14�"��C6U����ޤ6x�R�~�����c�>(���*��+Wֵǆ�l�4u�m�H����	=La��� �ΦQ��>��q�cy{���2�^�Y:߸hٕ���B�Z���K�|�П���HFa�a�*^��#�����
�*+۰��)�b]�h
�K]/�}H�C�O��'E�:�B(O�L��*+?H(�Ǥ��,���I����ܻ�fo�:"N��vR:�o�ⵕ�$l�@��Ƽ�8�&yıq�S+s�*e��:� T��<��.�Ԭ�G��D7�<*��+'��@k�B1'�bT�Rt��ם� �'�B��9.����s�ͬ�	#D�I��&E�%�
.�l�wdnD�d�k������V��v��Wq:�/(M�J��Y�������4��#�}՘���_J+����LE=��[��e��XW�o���VNݡBK@�J�$��N�C� G��Nt�xP`���l����M� }`�#k�IR���M��6AKG��A`�[�r>{�g��K���t휽��rSN�_c𶇶���F)�#60�ԟ��(��g>J��O�1������SRx<�+>3���1�0�Q��D-'�Eֲ�@@��~�r�1�e�jJ�����b<��M���Z���H ��a�%~�`iœ�7���꛷�n��@6�ik/��;����������	!�&ʽ���|+X��ls-.^i���N�U��;�R��#݈2�H�M��c-�N?��.��jjȻ��Y���V�j!_��wk�j!/C�v��r���4T.�d�@Ӻ��`�L۵uW�����m���ɜ-�K��̜l��K�i��Nn;YI멧q�i�k8���3K�6�pw���E�@��޹�kD�+�(;OI���Q:�ꐥY����iD���6��SKj.��ki�_G��T��T6�#*����'�e�������A�������$�����p����I�&^�f=������n�*�`"xqi�J��g�CWۛ_���a�X�&�9@K��EQLౙӈ�ُ��`��PQG)3⹼�:(ۋ5�黏�A.m��I�y�~g��$�]���B��3C<I����B���*�kW��ْΘ��A�����M����d� \x����!R��0@�S��L�����b{�v�|�	p\�>yvLs���_[��Z%Lw��!�~ۼ�,l|�t3��!} �2��I�:�ݲ.m��9��7"����σ�d���u���H�njGg�p�+��8O%�R4yS����ҼR;�+���gGE��� 
+�^c���V`�Y�~����*}qDy�K"\j���b�nxJO������5%({�y�x����ҍ�����/��K�{W�&+�+ғ��w�1�!��c����2&�����@�}��7�{u�:��A��c�8w֏���$}z������=X���H~9��K�m�2�37�[U��V��Ew�Sg����J��wq�v��/6�y�ߠ�fc�M:/��]/�k�vS��%����}z��؁�)L����&�1:*};ߜ��n���I�����R�2�
qG��b�Ϣ�c��	[[����]%}D4���˭�������K�)c�8�����:�!��v����͆}� �������
J�Ϋ��r�4x�]�2�G��J;4�,��w�9`��Oڔ�@ݏ��W�KD�r��jT���O`�Q��RR�AM��,ӌǢO)�@��Ug!7Q�aW�~&uq	�B��s�h	ߢN�?՞`�0����N&b��~�GQ�#���n�� ����!\R_1%k:y n�b�,t�z??�!Ҥt+��V���b[��
&�������Ս���=M�xhw&i�5)�� H$/,;�@%k�>����!Z��	�R��J�8qf�b��q�=դ���i�)S�R>�ݞ��ܛ��Y�a��+s�����۩���o&n���X��ٔ��>3���^�M̮!w�sEC�a�,��%��%��N�k~��%/�g[u��[9F�ꈵ���"U&�BP�|R�vd	_=��Nt��/^����F��D��M�����"��wC�I�誯�c�S�Qe���h�i�wu*2�^�j��y?����;m�j̜�:�1.��8z�Z������Mug�z��-��x1�eg���~��49�,o[�&���p�!�O��1�T���H�K�*������8��`� 89����{����N�B{�+O/)@�������<m[��-*X����i-���o"��L���E#o_sH(.{_a�1��|�|Z��U���t	�xS[�h��R�R�f�6lW�I' V�۾c|����Ѷ��:`P76M5u�]]��"�� g<�~}a��K+w�	ݗj��.�*CJ�U�aLs�e��ڢ�@pP��#��.[�&(�z@�>i�b�7H�Nk�bX�^+m�3*�����}�*Ex�pZ��l�%1�@i�X����6�v�qUv(K]|��yb�����9��r�:���R�Cx�e,��h���?��K��f����e&�Z|ȧ�H� ��U���I���P���@ҰH�����7�h���a���t�4�Y��W߽	��Mp�9@��#���{&��dO��<��7Nx_����1PE����bqHF��� �ѡU|�Q���5g��e����*�Z��
��0��_v��q���������ɉ�b�������z�֧ݛ���D;��j�E��4+����L\S�6A����F�~q$4����ɉ���!	6M����*�rY�b,�P�2�K�X��QwD��#y�!ϑ���������jۉ>N��Ċ��N�_R�B�l���qS��9Ǚ����b��W��I�Qj�L�� 숂 G�T
� B��f�2*����0�o��;��Q�?@�I%��_���tJ$]��U'�A!��9rZ�_F���,fU��8����^�GDBN��[�7i�[m�U�Mi,#�'�bL(��W7d�Jj����¥�q���������T|6B13Әq�hg_�/����4�ğH�8�ćK�3����a�(�#]�'%Cu-�\ň�����2��A~�@ՇDAu|,oP
k�,��=u7��e�S-��.�n	ϴ�:��Fe�n�T��+�sY��	��8a�t|qͷw3���Ed�)�:ôTt�!�}�c��EcU�IUk�?�T}`K}�A��3�
�I��F�wE���ͣ3��^V�,���z�u��C�&v�k%��6�j�΄�L�8��ֽ,Qp��_J�u��OXp)��6���]6Mןc��Эè� 8sj0�y\��E&z�+�����Q,���Ǧ�]ooT`֥�!�4Ю�ex��#���rZR�&-�/� �	[''8�~3�qn����In�:�)ɼ����^����(�=����hܗ"n1�F<R�B���2+
���]�8��A ����z�E�y������Y�����hO�Ѝ�G&�r�x����u;�Q�|ìt�PO!�8��P�!Qe�3<fR}j�`�*�B��4���4���1�y���e/�?�(��i�飐��$�"	RS|�9%g#֖��7���n�4���e��]\ÇG�8T��KF��j��ֺo��lP�%�j����7n�~zӋ��:/���׫蟤�ߢ�^�29Ɗ{�ߔ�����g� ����/O�����b�[E�/��i�b}3=�]�E�/����ެ8�'�P�i���0Kj�d��lS�]�� (Ih0[�r�>� �%Gډ�Ш0{��]+��㫒3���-Eί �\�W��ԋ�,@C�v����:�Y!�#>4�2��^��ʠG�82wT�v0/ߝ�;ky�?��T!��iy�d�F�у�2��7�D��0��}ln|(�ߦX <ߖ�C(ށCrA��1$$�Fۤ���Gwu����d6�}�$��ܻ�n��	���)�>����O�5!C �-�� X�~6�Y�8�BG7��	��s<	=��3����]����}��Dt ���Sԟl��'f1`P$�����O+@��?Ʃ�>�j���ү����XW����ŷ�Xf��b����u���W�@�յE71�~��I\6RtR�B�����$"�=��om�=�C �����b�x[	i�W�f�&b�����LI�9��Fvx��j��K�����B�L�� h��N*�g�������d���U6�F���¤�G�N*��\\���MR�hϬ{c7VI����VW$T��v��~j\v �� �G\az����[�X�o����ˊy��[3o�O(z����Qla�E��*G8�I��F��pD��AQ�f������C!4к�U�Gtm��rڥ@����!�u0�X���"���0�g4���������X{���Gk�v�h�e���&@��M��,9V#�
���'jKq��nR{vAI����t�p7�J:dp],cF������%�����x�S�G}R�մ�2��8�� I���Zq���(!��
F%���w�hP���&ٝ���&[v�c]Y��K�ַaD{ �@��� ʨ��Go�%���0u��3{'���*�V���`S����`>�>f�*lq9~�T� ���򿟳�XS�-�_~�%$N�O��j!`����5mʮ�A2��KS|g�֡㽲n�]y?��n�N#V��=��4ឱ�ga��A<\`r-���20wscu����L��#�*��u����-դ� >f�@�"!%����&��c�`8����l� /�՛)ۃ�w7Ur{NBr�S�q�]-?S'OS�h��@0��/fQ��!��g6�n�T��t�xP)cŞ�w�tQƪa���.)���l�4.?�
e=2��V���a�!z�j=So���<��Id�~`ٶd�@ ��8����8w��+��E�L�+"��K���mZ���x/����F�4�[�pm�YN�l٥���d��4�V��W^�����_�Vw.�cW�G��ՈĖ�Ul�5By����gT�J?�A\0<]�&ٻC��bf�/�o_��C����,��G.%]NX<1��v�17� /�EыP$N9����10����<N��d��}?�J����pɕ+�L��Iz���9ȉG:��V�)��P�\��k��/�z�e~}�_���0ָ����q���j���g��L��2ox	E�:¼
B!��n�vlQf�*�%Jr�dt��{?$)N����]5�'덱��?Ӥ'���2��vb�UH;5;?�l�D;S�%��v�ɩ�z��QX�#\�0 ��,�6��1@5%}��i�i�d'����a9F��C;�u����w+_�)q/�_҇�,�`����!�¿w�G$Y�ژ��<c�[��@`f_�.�U��Tw�;L�3*ъ�f�'Т@$^�+��j�;���
�,�M�S��PN��rݽ�P�J��������r��0b�B��^�H�$�镡H2w�?l�a�e4`�^#q��-�
W�USD[ӓ�2��_��-{ԘZ$�:�e�!p@�ZzzJ���.�?�a΃+�$&�jG���t���-���m~���ٖd��-�'l���r�<���䬂]��	c��
�����:o��t���{��e��@�G��>�a]&R/l�jS���\����yarg9��[��SI��]_f|��k6H�'&��"�+�u���Z�CVOxM勾�E:�s�C�_�
Ȩ�������"m2�d��gD#�k�|�0%|+�9\�2��+Q�H��e�.���֯U(a���.�o�U�`R�����3sl@�?Km: X�-�vX��]��#Q���a�g?��pm|��ǋ.�Cɧ��#��7�G)q������C�"<���,ѫEK����f���"�V@ӆ�m�j� �(���dM2���<8�8C�0�XG����v<�3��i=l�q��V�q�ʌ�;3Al��#=�UF�C�J�"����[$�b�;��������<y����9�n����0%e�,��[�畱�O+Zk�0�|~ e����XAt�6ͬB�p���0J�蟪��O�x��sq��W� fz���E��%w��F�4���S�n�ؘE���O��8�JZ@fĠ�'���R��6���"|�i�g��K,�䈜�/��:��u�}RP�;�>��,Ѿ����(̕A�~�(A��i8H�!�%S�xy�K�lV0D�Sc!(�qL�_Xj&���Du��i�ϒ�� Īk`DbU�K��l]f�>��2���f�goKݬ�Z�,J��a�����Ӗ�R�C���X&8k���UO�k܄軥4�j��@��wn�>��� �κ�|��-SL�[ţ�Qӵ�9���\鵂S���¯;�����X�70���z��d`[u���D�����[�̢���qu��n���6�2C�Y�d�:��>}4��`Y�+'���܉���y�#z�V�s̎p�2����]����C���)S����;��$�CJ1�)��KC���'G	��d)���O"6"������1u��W���e���l"�/��������ŉ�c�\�5/G��E�;�:У�����G���>���P�B"_j�Q��$��6�G�%���p�/a�zrެ�T=]�����V�4�	ќ�W\d����Sa������Kݖ�^�m�T��k���A����-��!8�b��Z�D���%܄\�|b��[�������Y��lYk]q�/�n�k>��l���5�|�B���=�]����F��*#�\�\" ���f�����q�_�٩���I�f?�O8�C��斔ʀp�׉��RE�A��
$;����ă��2���Մ���?�r/�C�@Xbuusd��Y[��}@=҆��,k�?�<�(PGv��rfy�f0���j�&�P�0���%Y�R���tG�/��t�"�h_x��^�n=�U�a'�?b6���S��ޟ�$YՅ��of�*��^t�l��Q�>Ó�ƽjf�n�k���~�o�������uGIfD؃��ϲ?�����&�>{�
�$4T�޳�k`�@X���49LV���#���\�_PO_�a�8?q�����e��J�n��i>>�d:謯˼�3�\y�g~�/��3v�A.�!���@Ӷ�����ˤ
xŴ�-o��f�QF�L�����<`�
>�������c�^ȳ��"��f:����Q�{�HE�H��a9���I)~T�(�9��[���ī��U�$cώWy��Ϩ�'�����(Y��?�F���S{�F��|l__Z|p�+��6[��.�.8{u�=�Yŵh�J� � m/��[�����ȓ����7?H�Uu��xqW+�Mp�dL:�Q�|g�9֓�z|�Ѱ%j}���%E@9�U>z�w�/d3�ʖ=;Qzzs54Q���qnT�0��wC���y`�d�����~_�$T���E4V7�w��H�쀒^IN��Ftԝ�����Ms\$��&Ө��{d,�\�N�ck�Z���ń�h��n,4
~(��[����j����+�M���5力���$be9W�䙣<֘RKU�o�����{�i�D�.��O��4j#�r0i˟���ȅTA�������5�R����~��c�7��>=4~!t(|�=uʤ
RC_�� x���(��9wt���>x[b�
�/�J`�s7m�b�slɦ��5��R���]��I<1�+%��=��"5�w����J¢�c�7���n�ycyv	�!=b���9��2[3J|]0�Z��]n�M#��)Q�W�����VO�?i���'~D<�3*�����..n�tA
J\�т=L��kt����X��M���CZ�Wk���Z`2�҈S�����l�;�V �p/�e�
�x����f�:3�Ǚ-��.#஭��!n#���!*��	�*����A�5@21�t��1�C8�����y�o�x��!�T���f��-u��(���\��:�؇-]�ɽ�Ҷ3Gq��vӄ/2Ȧ֒-����xf>�>*�P�J_��㹴��x$�(�⡡��_���9�폭,#��i���J�{� �����eQ��D�ܥ7���_���z/��4���,�� F��ruk���4�P&�ŐUF����tjqWgn◦n�0Gr�i;����Y,U�+,�.+6	���~�k$4�q�����U7ђFa�[�jev�`%���$bO�~b}�U��e {�Y�"-��7�,!J���
��`�w�ZDߊ�����SܼE8���;�����ۆ�u��kOׇ�SM�p�S�"ZH��[|i�_�+�{ōhL�4�u��Z'eW�>J�Cn����c�^^��矟�;�J�cYd�z��p�p�8XLюH�"�Zg��!�l�W�5FZ�q,*���Z]�>��3��dY�<�#���{�Cl�N���px�V�3�����]�To�T�R$f�f���/GK6�����p�6WvX'703���s� ~�1�8��f@�����n��K�T��Y4(P2�!=����h�ST�E� 1c�$}b�|�!��``#��sO9��D����`'FX���>�R8��dms��c����ZVw��6��(�n睪����/�_����"�"�)�8��~����)�e(��W?����垭��YM>u����g�s���}KÓ�Κ��T`��BLB�˦Q��w�<b�Y_'�#���0}�T4˵}�x_�Ʌ�	�������9(PWb�z�j�Pq������ݴ��{�@պ��8��s��0i^ը&�1�WZkr���7��	�u�ܡ�'�����A�y��{z�x(��l���&�ϋ��}������ju�L[�o��g���
�ɖX۰�*MJ�Ä2�H��I)�Ae�*д��菇�hm�@>�o��GrC>YU��]!A�����s��L�/�~|�:6���t��WgWU� ��91��A��<bW�������u}�bm?u��L��򭹨#��Y��RL@�q�R�d�Y� |@�vh+�仹C5�-P��^S,<i��2�TLHc)����jߒ����2���PHš?C	�Uت/�qu��?�Y����T��꺂��F����d�߹v������~ �F��"
�n��v��<�Rt���.W��[���	u V\k�|W�+�˰�ݕ[���}(,!�h!K�l$t��]�����i w&�f|W���#?i�H���n�fd]w�U��i�D�fe��U��;��$�Z̙�v��N��L��K.o,�XOcJ�p�q��	���h�pʔ�s�]�M�p��T�����c�\����cl��*�]�8��j��ǙA���1��̿"��X��x�  ��D�~�.�P��+ ���7R����IP\�h�}hmy����Ӌ'�^zM�4�n�Q�?k��a��^U��!C�j��;� ��^�Q�I}VQ1��SrpT�5ƯR��?�z�$i�ߊ�<�����*�c�bp"BĮLQ܁�:�F��W/����=�'���g�-{S���b3=��H�ct���غ���
M1��Q_kS%�>C��&�w��)����Ƃ�����,��<����~0I~���~�>���i��+�ݽ�� &�����67�G[%�Z����a�P9<Y��`=�{����o��݆��kG�ZΰƔ�}bWo4����3O��1W���v�z�� ��J��ȴd�@߹�{`��u�+wnl�Q�F�q����?kÃF�߂��10i��kG[�0$��,AZ����݈Q���){!*�37M�*���t��֡�n(LZ�9X�	�(��md�@�M��d{��S�Nz��p�������<0i,f��jL�m�VZ�j�P�>�8��O}��I�*�8]1�v�O���𝸥H���c̩�Ŗ�0��W��k����'9E �E��@�[CB������� ��~8���7��qx�#�DC)<+�����&\C��-�V%Y��R�rS�V�LU�
����s��Q7����R�Ȟ�V�]��=�ixdn���2�ߪ/���:S[J1���D���?%{+M�p�`��]C=pIo
}��X\p�O���!5����1�7�«"���+�{K��VW���z�s��黦�&H-���bΌ��2��z�8�Q�g��Jަ*�JE���i����c7H��o��~�%G�C2vE�
ߥ),�q$���,Q�I�n�ƿ?F��G�ߺ�{TL�+����pjܯ�}Ћ�f�������@,5x�RU9.],�goo���?����9%����%g�D���|MZ���L��֕�Z�����9oA�]�����=��8�����u���3���>e�xE�S�A=K)n����Sg���顒]O���	�{F��O��b������4�������=�4�׫ރJ ���a$���ʸ2Aq'�me�(��@�Xx�x��ᒲ^�������c�O�Uf��zVB,U��"3Rэ>"�6I��8�Yq��f�@�����ǤT!�R�3 ~�H���W<�W���,Z�n��]�V�O=�`�b=ܗ��j�77�����(���Ȇ�Ʈz'��q}g�<�g�����9H��U��N��3Z�7�r.�������v_�36�V��,�a�"���yhC��3��Y�}e=��jT�����i$���&$-�0El��$��ckW�v��⒜ Jaݨ�
��Нǚ��	O+v7��+�"�CTZ&��<��ѡ)Cc��=+t�����͜]�E�E�[LR���TU�^�ݵ���N.�$�'���'���O#� S$ogr��s˼)�N>�G�m�-eG%��yJ�l�m�Q�\)�a�H�jz�,{c��:�ob�C�pJ�HXy�U9�":���6��>�!4o�������EgTd����x8nKe6r�-܇
�=�"ݿ�����`�$q] ��1�Wh7�YY�7�q���T��0W�B��F�$;kF��u�F����(�9? �UC6��z1�+Qlcl�!�箺���}�
��6����[�#]ìb;w�PHt���"��ũd�=�r���Ҁ �����^��z�� ���(�8������k\�ga!�ݥ��L1�JU��{�JT9��F�6 �+�2����?�F*{(�W&P��VOى�|/�``rz���!��7@�SV��D��N���F�y?�&�&� ���t�ȑQ�F�r�y���`�Z�6~h�_'�03��=.7N�brv����؉8�Ŵ���c���ﲋ(���y��	���0F-.ቋ��t�@B�:� ���w��~�\�e�\�C,ʜ�3
�^֠,���jnf��E���B_l�����?t�]Γq���I��a���X�e���i�0��C�T���?�
h�X�x�Ԟ4A�-�*O� 2D�$�j:�c�{t�Z���S[�1K6p4˖&���U8v[��<���q�L��k��Ĉ�!����I�=9G~P��>-Q݊EA�rp@��y)MǾ]-�L�,çFo�If��Mk��e�?�*�ɩJ��|s��~t��m^�E%*��o?eoy���Pډc���x�jV�\<�q��#��Uk�eg�ĉ"�1� �]�Qc�n��4DJ������������wh�s�F���ǖ���_7*PQ PĮZ�'�g�<7�,�ؗ�4H�(��(���hT�+��B�3�*��A$:�S_!�@���s�2����5*2#�c�4Rq �ڗ2��S��0�"�1�l���@R�q�X|��赛���&�1�n����bFt���N#�8��������G��#� +��Q��pY��/Ğ�E�j��%��i�����+XUҽ��jH��Bs¨� �x�Y�.7*�n�� ���|�՝җ ���H\��C.�@��&� ���u<��qd��p�-�`}y�]���[?�vȧ��)+RY4�L��֨j�e�@f��;�w�4MM��Čޘ=�$*��=A��l�\���rd��R�g�x����Q��5��4TI��,��(�ExT�-�i)���,�e�ơ3�Ǿ[ɴ��_`^�`���^�����f?`x�<Kd��`���B�q���ܳ,Ήc�!�R���W,A?���P�0���t��Lg.���}��QH�6��0^�e�Μ�o��,G��:��|/�G^�d:�6��1��o� ML;��ۋ�1��O�=��ȶ�bQ��]G	�3c�;%>�\8�.q����������5�.�IXi�l�2+Q1��6f#�&��,IϦ�b1�a&5j��{j��f��u�jHv �3'̪tV�|�ޜR�q����N� �?���;�RpL �ʋ��Kx�'M^�q�����_a��|0��9�ഘ����h[`�����o��gԊ�fL2���^�Ę+�^˚��עSF8c�1+�y���u�E�NL��cbZ�1T��G-:o�0������^�1��U�tKP��ŭ���������6?d ��:�J�>�*i8�kd�<��b�!є�^�E�I������}�+�8�k:��\��ɣJ��0y�%Wz�I��G�w�+<�9L���o8�..�e�g����<�⾾�?Y��e ���� �c tt1�:6�^Z�In'j����p����"�3���b�;{$ۗ�,��(�-���N�mi�?�6�D3��K�����~%L��EY�8��r���]B�l9�U�*c�0����7���0����'���(=��1�CD�"��	��)����aTe[S�WFh+�W�v�8�Rx�����2�)8� eĥ�����R�ו�&3}��D�2=j�G&x�_�-�t��y-�>� �2��a�{���I���#�%^s
0��'yC/l�8�Ȟ�3�43w8q��`}N]���a��ݵO�Fp�-�%�G"x���٬.�>,PD}v��Yl����.O{�8n$%�O�Z��N����HZ�)~i��:V7�F�U��⠖�ڇ�k4i��4�)���� �,"_���*K[�/��=���ӏ�)�)[rM	���	�:��R��w�<��]���
f����/SJ��^�i|;���>�ao�c�Hi�4�&e�2�݂"��N��`�>7��w>��UR��A
�B�[�$�� Eg=Sq�d O�M2���RhF�qR)�]'�}"�ކ��	��������Z|�U��N)r���]i��`�� �	V�)�<L�d���K&�������K�{�B 5�q����`�w���
�7�Gh����Ҟ�K	�,2hy���	��`����ĕdJ������B�w'f$�j9x_����M�y�*
����?T*tzv�PCm͒���:}����b,B��I�. �~�E˽/�O�ݓ�i���抜��y(j��9�i���/<���/�k,���fpj�������V�v83B�ֺ��D��6la�Q�D�������<����ZZ��Q�3H���MǄ�#&T��(}����@Y�g}�T��J
����vҒ>%ﰬ
����ǜ�����oޞZ��a�
s.�A�v�U=���'�ً��6�s�K�N�z��0�NN�V��9M��)? �s"��M�e}�>����)R�d$#�bUu�]���p�)���T������!�g.$0�:y%�	��#ϞY�q�SZ���	��9gC�S�ܖ0�=V�t�{��P�Ҝ2m�B�n�z~ٌ ������rO$���G��Q"�voY<�?�M���͇ͪ����o�%��X�T�pcӇ���Q���2�ʐ��L���'���
�{-v��}U�7USG�������@s�S��i�
�:�͍G��OMH�kOrg��Yn���}���ɌѺ"BLB�-WbiC����,:S-բF=�}����#]u]��Oԣ�zCW�0��5���������	k�@�+��夂�y|*mP��t����#�\��#X�-;ɭ/��xƄ�l$�dQ;��(��d�KfϞoB�����j�A��O�`�`6$�6K�������	�k�i^��ۚ�=��2n,�^wJVA��uX�`)>ڲ��H�z��X�b�eB��K�����4]�;�iyP�L��&yd���X��t��
��'���!s�/��I���]�_�܅����i�ig�9�w�U?��J��W���l�$�T����"�	���y|~1>7-�8Z����!��}k���qZD[�b|��d(��7�
�P�H�"y�+V<�:�"΍:]1�DzR�]7'�fc7A�X�U.cp'��'�?���o�
&�>�C|�Ҭ����Eq�Yʼ+~�'�&G����w�N�Z�Q��+����i��L�R��"��o�r1�[(0��e��\��5����6C���fp�ʯ3<7��f��YEq����� oM�/a�^�C��x��/jt*O��wu��=H��?.2;���"R��aLy!.��̙�z�d$��as(���~+�^U	���ȯD/�t�ͫ��or�ďj:�\G������!ܧ!�m��	&ڗT��PS����� $wf�F�V[N����ʹ�ԸL`���𛹥x=�(�R��5}����)sVJ��@W��<Ƿ��W'��1�J0�v�
��T�E	�_�	�+�j##BbZsF�	����-�s\f�tg�����׹~�^�)�L���2a�?�պ�[o��B�[Ċ>�C�FM�):�>�Z�	D���`��l엿t3[��@��Yߗ�{Ҵ�b��|�L����0�����R;��,�*]��C}:�ب
��L�H'<��A����S\?Z#�c-��>�-��L�C=��c���!�{�2�ƣM'�n.�H�@��4���'	�4�s�4����)�˭���'��Evc��s��D�[��h�+nx��~��r	[�2V̺���l�a���G��U�[��!k��?�Q�z]��J���j@�x�a����Y�W�g�'2�O����\}�&�O����{�PwrsZϛ�����Jv���g��x�"U�s����;�@�"|y�b^�nS�'�
{���]�>9�V8�߁h�(�����߭X$�?^,!1���� ��;�@�78��څ��6}��g���D�x�ΰ�OE���R��:�=�Tҙ�n����2��H�,d�k7BD���P���ak|� ���h<��Jnl���m#{����T�e�Y  dC�u�y?&Gd�q��4�n�I�a�I#ll5%��(Z��� l֣�/�~���םO�nt���*�~rOH������?��_*y�>���0e�Į4iF{�j6��^�h�,��[�۸7�M����6��YgL�H)rqD���ƹ5�c�`�����.WҤ��hO����z��H���(�aGE�%jYz�W�0���(�.�5N���jC����2۹#���bS�� ��q��@0�4O�;v/��;�Nh���JH{M)����B��?��N �f=g�Y�����r�겛HW�۾��Z6�'�`��,�3Â��S��T��v�0��>јKPה3�Qn�͸���(���=O!8��~�zD��M@��zC4%v����ap����?��Ws��)��H�lR�S�`��G�ԛ�n	���M=o�o�_m�/)���9X��r�g�� m����r��$\Q�˲*nr���C��c�����~�'b�_A��+a����8D�h=�v��4뺔�ɟvP��p����E�y����2� <"-�:���GZ�H3��vV�!��Ey������E��Xe�Qr�ш�݌%���Z�� QH7F@*#fzK�6��\�M���U#< 0w�ҌE�`�)7�3R�W��A-����|pE(e���e��8ʛ4�ɴ�!�YP�^^f�o���e�Cv�c,��}���՜��H�7�-jY#�%qtNf�Uj`��o����Kv%���؋���y���'�&���d`e���Ί����Jh��8Dh�<���oD�A�,�ĳQ��C�n��n~o>�m#m�Ď$4�%�5`�J�S��ms� ��)�P����ӊ+MD�S+�6{w�����V`jL���YG��a��im�v��$�ƢLv���`�F_qSۢ�>g�x5�K�&F!s�P� �h�����<F1}�3?±i���*��w�C2�sL�d���i;�q���`��H�c�J�v��}G���-�O� ���y33���{�`+�z��Ԋ�z�� CK+����'Q	�N�JO-�X���x��l|����"uE��
�;�x����=7JJRr�G��;~�c� j)m9'���!�Ӡ4�w���)݋&O��tI%8�����-PPHu˂�Xj�O��d�@4�}�1 �fT��;���wF�?���jt�
h���̣
�
�X���`���!����L�F�M��Y0�Q}�E��%�*$�R"���OG�;y)�+ ,$��R$SND!�"
���t-j������U���lA�V=�G���lH���5�mnc�4hg*��I׆B��� �x�c�@���EB,�g�L�,��!�Ь0%?q�������j��4O�}�Իd�ྋ*�M���7�CĨcB�֒���f'@�x�u
eb��S�Ñ�����
�~��8F�#p���h���O~נ����CG�u� dx���&�V_����VUi1/�90 �0�
�(���(ki����\��׬���!�;�?�&�J���L�J��0�c��3%�.����J³l�w��=1}��~�~CJDLWT�6��Ƙ���#���%O�H/��Re�N{�����n�ܰH+�]���0DH����u��ڥİ㥁t�N+�
�J��n=q}vސ5-N7���^N#���K��_§��!��No��8����r�O2����n��h�\:���F�B`�rKã)y�̘�:�e�L��R��W�^���c	�bq�r�o�����	?�����Y��jĹH6����i"�%��Fl�B�d6<�8bz���1~̅q6��S�	�ĉ���c�������}�<�oNw��8�՘���ǡ��O�۠�d����H�49���!��}q.S�J�4�)�qz����a�`�n�;*��F�v]�;-[�L�|�'�b6�)�B	[
((`*EZb�~Ԟ��1>��L��r��'%V)�\�m���II�+��\R�<���E�P�}*f�^��W����x_4��)n�_�lW�ψ�qZ鄒�a�@9��Т�j|%���5�ˈ���ujL9�r:�Z ��V��{7��Pu=%�ݰYG(���j��U�Q���@�s�W��+!<����������uB0��[ �X�������7۬�-܁W�Q66=.=ǡ��jn���R	�h�ɒ�/��Z0�A��]>����>u�P��\xk,
c"S�ݲ�t�F�>o:��G���t��ێ��@��WO��l)nFQ��H	���W���FP���]���wM����ˎ�����\����K�D��q~ �����~�R�[:d����ya��0%~wWF30
��m�X�E��F*:-SX�W3�u(��2uLc5�5��e�5x��������fgr��E6��=3�ώty���<%#*q���l�Գ��b��쌦�<=��	�-G{0��6��a�R��fo�����"�cΩ���϶��*^�"p�.x���m?�,����Wc-ģ!K�/�8Ⴖ{�����t��%�4� ���) �V�7�^^H��LR���퓷�>�9ͮ_�37+H0DZܺ�<�4�ZŖ�W�5�z^�Ơ�^)��y�}���\bç0�
��jT����S��ZS�:.U�	��t�s�^�eMh?קr���d�,S5[z�V��j��ğ-ދ�n3��(�7nKN�L�5z��(*�O������~9P<��Vf���۩0D({�Hr��| ����xz��G��Q4�2��,�<Vj�;1�ٜ�����q�0iF��Ɋ�C�u8Ρ��.�P�؃H�-���B��V���X�J��:�AF��QA ��w��9�ή��3Q���(�NYdk�zFM"����鈦�[��d!_Sg�@R3gY���b���Y��:��t�/[�w �-�6��2V���	h���HG[֚��ש�b �{�8XqCM=C��A��489�<_���+�	4>��k�S��<!�]�,��P�zg��:����n��;��cK��`M�'}J�쥡��&�˵Z�H[���[�.�w�'A&�Ŝu�1ݗ��kz�����p$r5L'��3�9C_l6�����{��C+T�k+;���b�4�M�l�K�W�55x7�m���8�S]�p/r����w���g��5fS�q�?�pzw��BI��qf�K/>j�2>��g�����`>���`��	m����j��7�W(�+5��[�d.��eJ�1�5�ۀ��Q����$p3�6�p�s�\�����z�Z�Ӧ��MI����xs�t6H*��UOw�n�NjM��.^9��-R�y���u¹��v%��׌?����h4*��m�r���������AJ��s�#rӫD��>��}WNeV�u�r�\�!<b���(�D/�⣩V�\х���&��a�4���%\9���+������H��S��YN/C���1��4�o�����/���C�l���|���B9����G�{y��+�!�x��N~�3B�#CmJg*S�/�+C��dHxɋ�Y�	�F���&$���RF�*d�|.ʹ����CR8�*���V��`=��;V�a��FsEY鋓�]p�� d������#)LK ]3ʘY^���pe/{K����^J3S-A1g@�����700?����L�5��)�-+(o�z��E�%����`V�n~���t5I&A���}�F^��O�'��	D 3ڟ7�pֱ� 0b�zTR+�� ���x
��	l���K
1�'`�'>���ns�a�a3O;m޾�*�Ev��^���Jd4(�\���S����.bK�^��e�F٣��o�#�m���ƴ;J�I�z��~(�Ҭ��>�|\����wi���H�U�6�mY�)��V#FX��h8��t��������G���n~�c>\��Q���k�bC��J��p���gF:ϭ���i>�d�p��� ����i�����-*]��̰bs05�U��	��usmX��yH�/��\:��9'sK*�4�oSg��7Z�k<n(�� #��O��9~%߁�S�!Q��>�怞���rT0�|aƫ�}����u�b�l����U ��a�J�9����|&,���pϱ��"�^��[C'��R>�ٕ2��5сz��)���fS�P7��������Z��-w��c�A�� E�l�����Q���l���j�o/�����s@�7#�}�AZ����~�"���}�-�Z�dr�� QZ��{���N�SV���t��Y�+*�W~A����¶���jz�j�S47��b.\1	_ �.'s��ا�J����v�0e}�o�y��A6�����Ym8B/3�4��$��Y�ζy�LY7��|���}�-�
��"�����)-�G���X�lu#0����w�QeZ�t�V�.�VҎ}\��d�/���w�"^&�ř��,����JsA����� E�s�|'=)T^�3��ɦPח��`Wx��CFCw��^հ�)m1}'��&�A\�&��1k+p��ѧ:����Y>9mZKB�=v�Ab��K>�^WB�# ����wL��c{H��^0�-�r�N|Y;����
�����(퓾w�xgR����{�k��R��/4��Vj�����H�EeM�tX<q�j�g���Krs7�Wm�/���u��׽��f}�-n���=��o������	@�=�D�z<�����j2�F	��ԍp�KV&�� �0���X��l ��G�Ga�<����t^�?=�'_�{&�dm6�&� ��/:��	�l�W�Cc�C�I*�>��1�h�=��ƛ�j�֋6��%Po|�Q�,���n��^Ǌ^1m�Qe�.�न6-��%۳��$��EЧmn�[R+�b�zlޱ��*����`���#���A���4�BmA)�~�ND���P���̱�W�~�/���o�6|VĩF��V�*��EL�d�2��3����?��F�^�q�fG	���	�B�T̃�
��0xb� }��%���vI=}��&�#K�Ϸ�tJ>��7�Q����O�/�M�O���cB}2�z�|�uC�&�Y�_��I !с�\�7�p����Vy�$+�ړ1C��9p���joȮF�*;�4��,N�w�&yT86�j�&7��+�ܾ
�/���ԋ������ �
�����y�-�Hk��V�*5h-��Q�5���ⴺ�	'��G���.���A5�yV'e��*��4���2ʱ' ��v��V��B�OW�H\]A\�9���_�	Z�Ih��F��>I>_8��C�j���J�|�3�F7J� L/ۜ�ҿ��c�8�Y��<�@��x�=�Ƣ1�u؇X�@��U�	�+k����/��æ��TV�0&�·D���cz�}wx���\2:��'A�+�y����O`g��_�œ�(�N�p���o�i@24�h}>%�������8�����m�)`���f������_`��bv��yE�H3(^^�r�����"�aAֻc����%"�HI�I4�S;����]�X�}�\tKSF+h�:�12�S��T�_��uw�aӄ��rf�n9���\���4�?��)���a/�1۝ �%�� �:��~�>����4��Mcm� ��:�	|ςܪ��Gg(M�s4�N�1�k8f�˼��B�mLFh�Y37ꥤ�cZ�1$u�۴1vB���G�ME&3IG{V�5I�&���$u�7�n��w4�������w��'a�j�/u��)0�/�F!�����y���(������;��T S̑���!_�7�$n��.�`���2���/P�pk� d��LҠ���4�.0�0�p���h"z��Y0�- <�;�B���0�'�4�M�s��>�G��Z��Ko]�		����	�_�@��C���®��8���	Zc��r�s��[�W�m#����ŪG��vWS7ly|���*���W�T��"Ut,.<���f3��Ԏi�mK,��/��}d�ZV_��m`�E�/N+_3�"��0s���;DP=�'ZOJ�H`���D��֭���;��|E��A�@�B��G)��v������]e2f�')�Oâ%OxY�?Ԑb��U_��،|C[r*�Lr:L�<���a_���I��Γ�OO["}�;q�?d��\0��8t?)
�|8r���e��)\������)��,w`�l��i�!��MH��R�x�=��|�Q���cz���/ � �j�=Ԕ�]p�y��s�ۣU��ƫ��y�[{���$0Cu��[�/%���wME�$_�Op�c	�e������%�u�%<rA�WRa�).�S`�	�l�f��O�`7;�ʙ+�s�ce�w2x{���)6�C��&�M/��fN3d�h�AGi��7d���[3�	(�Eb�Z��AS���@-�����,[�6�c���Q%��Xg���1��'�d�?׋�9=׌�ld�o �*Hc07��<(��2ób�Tt�aF���gK�~}_�������'��!�/h���D��X�s�.U�^��`&����:Nz��y��),]�Q!UU�<��7{��F��ӈ��D�_:#��U�S���}
�3�^R��XX��]�-	q��Bs�}0��}�M~�B)���! ��P	���g�z�V�����[V��S��� �;�^q��*dڢky���UP�:^��^X�5�!�I�P'��}��Y�d���aH/5��c��YW�����t�r�q����ڿF��q��p����� ��X�ᴔV�aw�Y��&�l˜2>�((vf ѡ� D��l�V}w�r<'���-����Njɶ[lIUv��YV�ftu.j�]"���(�9�%|����:@�0V󷕅_۴l�%�S�y�~##���e�O��lO <�'�T�v�V8�a�����L��;���;��tX�Y�p�l�B���T��U��:�Mk%�`�fW�uv�V�U,��\h���L��Y�s󇖸^*�f+�6+�����Bި���1;Y�K��4��M��8>sV"�b���>���Jܜ$�!~����6�re�v똿���~*�E�N���V7�	��4�K���NSƒ��^�+*�α��xS���|�%2�~B��a�)�,eу��1!�>�c��u�0"%�!�vU�gI�_/&�6_ ۧ���:�t��/�pB��_�* �J��3�$rv�_�飩O���;.\�,+�Q"@P z�z㸘�+C��!�H�/I��7��_�K�{^ }F)Д�Y����9��m.��Nx��]uZ�H�rh�h�΁iw�^;��l9�J�F��d��F:C��C��
��Vֵ]��|7�"ΰ+����ǭl\@<Ū�{����9ﻲ���ڂ�t?��]WV����v���"Z�[�#>-	lV��l}��I��~��?>}����|�����T/�9cٗ����8sBh~wG�gٙR����cc�
X�;�ܔYS���q�V��m�0��q��If�7�/�܎�|�C'ч�#E��~Bi()_����0�2�,�s� ���"i�4�����Z�ف�`G�������G�d9����\&ܰ��̑�d0�X�5�+����v}����rn����\���%t��pO[�B95��3R�EhB���yr{<�|}K,�;nV@�9��0.��f~���ER	8bt���*FJ�?��n#�����Sj���?��J=d1j����섦i�|�W@S�b�s$�����ׇI�@7N3���x�)���cb)��)��>`;�i''N֕!�����G�s혒j� `��پ0&�8H���K��l\�~�O�?vj�]�F|��45�v7�EP�2v�4�ɹՏmFl��1U����/K��/�Mх�^�q�z�2��cO�������o��������Eo;$�
�3�-��% Bzb�3��,��+��yX��s�9�d5N
�w��/��2������ͧ���}^���O�,��Av;�Qv���K�9���gi�0� }�]�`�����Z�r �	�������cY1��K��0(�Lc8��w�C�)�@
���BĆ��}�p���a�sy�ك8T�-�o�	��5�^c �>�>��t5��7E�d����$'�FTm;���c#vU�):C�Ɣ�nj��PФ�(t{�d��d0az���Kqd��w�>^YU@����C��t"k"�WC�\/L��Ӧ��ML�؅��k`mw�煛T�o{����^�v�XS���hb"%☣?�3r~��V2ym�]�"�y�K��RF���n7Ds�L�M�X	H�m��.sf�jT4��:5����$�9X���Es{�o1[8�5�B�V
ԝr�F3uI}$	[n+yı��E�΄:B�4w�+�h�
"(4M�+�v�Ym0`oP�PI޸u��G:*��ИhB;:�ɾ���b	Μ&c��"g�0ʰ�{��������iy�]�=�s^�
0BTk�ѹМ��lV)����Z�v��J_rjF5A�7�>�?�)���%75��4U����G�gN%�ʎ�@�t^Ԑ�E/�� iw���Wu�-�D��qC���Y���x���|�Z�cU����Yŵ.�uڐe?�R_����9}�{�ՖnZa���NF]��̒������D7z���6>D����*�/���� �a��z�ɹ�׵ $)(�o��;naq�����I���	�a�A�%��tǎ��"�{�����_�f\;��RG�c���[0�[���A9S��������T����t�����:�ƐL����\�!��UA2o��=K-!՝&� ڟ����� K��Z�L��H�~R�h�$���
�luX���{^��	n�p� �J\zG�r�57w���~f��E��P<��p�H5d�#��r�v�6r?I��{%f,����Fi�[���WJ*�q
�q�!M���gV�{T @�bND-u�	�79t���$.��xE��3��{�Ї8�p[�-�:^��c{$��Y�~{d������{��aM0ka���@פ���=���xm���ހ	���p�y�/_���A������;1ҹ�d+�eA���9��D�W��Q��M��?�0N� 50��9kV���Ralc�B�!/fE�����A�"�����T�>"���V0�J��L�go.@�f�E%`�{����B��(ɾ�{`����whB?�Hw��&T���S�"�D��j�f*6}Nb��W͑J/��y����+T�)�OXeъa����P��
��E��M� �./�}n_B��'���0!��2�rP���=?tK9'����Bl�P�ݽR�ӓ��S<�PH�ʋ��`w�Ul�]G�C�M�61�z�lt���$��� m�f����b�] !T��`;�xu �+'>S���i��"��v�?{+!�=��1��8(�`��(�M�U���]��/L���S����~FA;CD&�z�a��-�������ȧI�}D��j1������n~s~��e6�"
���!����uF���^31d�шy� ��� *�]��N,�}f4\|o3FJTfzI��)f��K�ͨhv�}� +-���1�w�ry�	ygA����>&�QH[�YbD�`��������<�!
lڑ�gKj���E̯?Rǋ����9Z���ǿ���{Aij�I���R���<�ؐ�+Ķ�*,E�S�k4,z�R2�����֒���}(�s�y$Vܢҭ��~k�>�}��_�4��g4����%��}����N��� �ޱ*5û����~W� ����x3��� $K��Yj�Hj�(".�4.��*�{b�]36�7G����rH_�G�*/c�����I�g�Y>#v�m�&��nۯ[��ƍRn⦥F	l��:�kߜ=.�k���5C/i3�Qt���Eq�)2`�@w4-I��{l誡9Q�Í���j�9�E�=,�ô"Q]�TA�&uX��.��}Anǧ�B?�����$�����8s�Y����(�j����&�o��2���!|&�V�+v�E:uB�����\�J���R�iK��;�<��*�� H��{!��z�^Hɱ��G^��[��Ki�D8�k��BB�gԳ�q8˷�.�cG�ᾝ!��#��;{``��a�رJ:(6K�w�~`t�����`���>Q�o�9e�e!|ݪ�5�T7Fd/8���tk�(=���7�N���@Vv%���S��.�%8B�t��2�U<�i4�3���7��<��5%��Ў^@�
)둎��+����yP0���l;y����?!�t8������/
��V����{ >��	;��N���I�&T���˯+ˊ��A�������p�5"h�F�e@����z�iU�J�[7J �~��mR?Z%���M���{�P�o�9��g�0r��{�j�'�ؠ�7�jl��bl���B�F�{� ��|�p7fv �ѯv6�rdԪ3�7�@8B�*d&!;[��'��F/d]:�m���S��]j�1xt�O�X��S1���ʲ*J���wc�)�{�.��@|�/��TigO����N�^�K���$�q� �{�̭�ڌ��
4,��Tqf;)���m�<�sYk�f'�<�.�=+:��2 [;	��k�it�ݰ�Sj�oe����A�c�̞�Q�F]���"�~dwa�r;��F*�����sk���p �t+���@'U��o@0�!瓦~S�7�u�o�_LB8�C�
b����k�ː?ِ:̛4R!���% ����E�Åd~�����C+Gێ&Gc|��ʍ`1d�?�U�m��s\�7�;�*-��-E�����j��5=n�3D���g�������v�)�?��ѓG=�z���y�QShn�/�F
�s7�d�D�wH�/��T���_��RË�M�����p�8�X)��+������h+� �	B��e�����Ps��F�D~�#R_� �	�z��h;`Z� �c��L�MI00��q�p<�4�ə�tPm+�@�ÙKnvՇ��UyXw�D0ERp{&�(�]�̃��@��� �|���N9E����u�\�,���G�T/���^%t�\�`U3e��V������nsX����>ƭy���{4���}�������.��Ť,'c>�'�
�9��nQ*ߡ�ϡW�ye��%T�:�;Fݺ.��6{5��Bcpaڻ�j��B$,KZ�.�jP�&�j�:���Z>�z6�����nn��u-�=7(���S_k�p�zOl̰*$'O�KQO:Q�t���ٺA��~l��p��f]�.(!FZ��q����_��*[}\�p� _�vZpLʹ�/��,�u5	xC�Z��?�N(��m�����)T�̑����[�9u�i�웳��A�!��6����y�a����V�x�tq�^���u6sNp8I��9�Y����A��Dѻ�������E`�+R���6+�@z�6�F��St k��]���v���`=e�ءK����I��l/+WB��W&�4i����M"��s��0�� ���G�h�\�x��o�$^
H�_�n�ʮ�Y��*��d�"�X���{�=!c-��A ��dS�^ۇ;��n�]U��P�Q#��QJ��{`%0^i�^;���s��6ؒ�D2�
���3JtM�Luѕ�¥�0��c`Z�]N���S���/xPA��Sq(ݜ���:�!6��"Yʲ��H��~M2r�[נ,�Yl�~�FHϮqV&��<F|��qh����U�c�{#a��X<%����ɦ7��h�j'|�S
���6o�6���� �5\��gb��;fDwv��2���+̛���N}���_����V2�.JH��8w����®[F0Gx6-_Ȍ�m�*?8}��ٰ�&�o��Q����������n��.�C��V�-YG��[K��(�xK�ǈ��U� '�xn���fW��ݕ0�K�1��"�(���-BV��}���p���KSiV�3���}�}ן�G���n
���+!����/m��S��M\�(*��x�`Bޗ{,'��V$�`�ch�4����H�+�-�%�����"�8�dn@LxXdS@j|ug��Z'R�R ����n����_7�I��N+��K�~MU���d�X�4ړ����=?/��\�P�hH�X������	|H~�8�,��IX>��M�#�>�ᆤ3ݺ��H���r]���<);�-�H��zNן��r�A��GOn��F�W������$�J<��mXVħݤ�nWf���ַ�0�d�>*Ħ�;G�ݸ�%���mw!�I�H��:�y�IAl�����G�]�%����d��}���%,��}Q=�0m���4=�H%f��2b+�<pրPۅY����fe�^�:��~�H�T�1����3��)�e���ԣ�*y��O.����`0`K��%v�O^-�NyK�_�ck����7R��z~�^-�w����y!a�+�W��$Y��m��Z�H�"�~�L�_��u�ŷ��D�vb�%xHD��p/?e���r 	dkDc�h�5^�S򆉲�dqQ~~��{���v��o�k�mcRcmr�[�0N��:U�u��Y)'+ye�-�P?��y1�/e=��A���������S��.E����Y���`��Çm.3E>}M=��ߴڶm��o�N07u�v��Ӟ:xD��������� �T��Y����6y0�1��y7����,]�,��ߎ�9�4�7�o%4�#x����;��q��wm=Dq�8 ��gA'6���x��B>�J��F�3h�{��_�/l�˷)����*�Dt�<3KŰ���	�6ww�?�J�P�0���3~�Op�Ӊ#5	������p�y��U�3k�~<H��n��Q��6؝�g���R����oC���e%o)���i�?���A��o�%��{��ZS&����X�Ǵ��G�04� �><ߗ~m�s��GM��_.{wG	�2D�}��g�P�t"C�q�fX��ة��?��;|	�;!G��M�/��?��B�6s8�-�Q��Z�A=&��m"��H���v|��=����$�v>}��������Ya^ɣV��Tƾ�g(�6rHr� ��N�@a�Uq�#��"-y��Z�kl�ʇp�,:f��b��Mہ�t����L�+�'h����ק�Uǳ��vas�˒g��޽��@���`��`���a�g#P[NL�������L֕�u����Be�gu�������C{rh�n$ y�Z+�a�7��{X6��؍�я��Nہe��X�LT�����9�5�Cy7���6��HiQ�̿�B�b`N����Y]XMT�&�`qtDA[,�{�q��-8Έ�-��|V�� �}^4��k6r���6�ʿ���6�7���+�·��	Ë��&��e�Q%,����4#��fA
���tB�s2xY`	x�m���@&����"M�f�KL�_,ex�Q��J�Y��y��J����53�jW��z��S���Q�7�K)#ii5�=�;	} |LZ�0��25�R���%n}'z*��8��7o�����UQ�W ������Q�i����L$X�4�����n��;UIhM+���`�M�@� yEo�S"1װ6�]������M*����׀��2}7�gC�����(P��u{ã-�٬�N	Xj���c�����A�d�F�:�17?$rT�״#�M���	P�K6NyM�H)�Gf�8�~��T��vr�a�jD�d<L���A���1H�h�DU�"�%X����
[ͥ1Bh����{D	2JH��<�PŸgCn0�r^����� t@��=A *��P�-/�K�6���ti	����yH��7}Z��]x��[ ��"Q�����:�Hron�����$��Եo�i"^B��_��zsv�{N�|���0��w���	�SP!��79KF��S�α6� 6�:fr9ɘ�}*�)o�� ���}s����="�#�i=V׊�y���d�-�4�3ά�Q���ȕ�̓����ū�N@�Š���il����W��ƽU�P͝`�p�48�h���u��"g�^�|�Ʀ��èGɒ�ܩ���ȓ\�@hrRw Gw��9��r�#
8A	xE4h&�퀙X���Ԛ�u5~�	��Nbe��q�ώxh庍!�{�g�fn}�Z(>b�qY��)����p�e@��������SćaK���zc ��V�	����p�v��y��ɴ�agn�#��JG!��:��.M��T�v�姆���`�A�|&jf���:�8��+j=�¡D��P����d�}<� ���g���˓��|��7�=�N��w���m�r�ج6DD��jR��nT�PP�x��������DubCC���'��$�G�+"/���g���
<�7Kƀ�J/�w/ѽ��cq�>4��;�9\�r���R���J/&�a�Q���'�FW�̝K�|E�4�ׯFZ�;R�?/_ؕ&K����ԁ�ʫ��ö���j\�f��H���<�BK؛A?:wK]���ݽ$6o��AqPY�c�y��#~%ϩ�Ng����Bjz��dÀ�a" ��"�m��`U�ˉZ���H���Z$�5C�������0��Ua-����oY���J���a.Ap��9Xm���G�����F4�'���r�5�63�0L�G6Z&���A�|`=Z�1����FQ�/D��N �w�a��j��1��<C�,�B��Л�'�T�rg��J��®��*9U�X#oox���Ө�l��Ԭ>�����47_j��XM�.7�@��:��ڀ��R6�H�W�A���k��W�4��J(�����_���S�i*nKO�	q���v����n��j�L���LA�f5+��N�>���������2\8�pYxӴ�w[�O��I��s3_���** ����	�R���@�U���]�ɼ?aVq��1��ٙ'�AM,�3.h$�f(�jZ�e�+�'E�ΎAuє�^ ���6�k}GI��yk̞���1��y��q���q��4����
\s�\�@\$;E�B켵�Ǚ��5����Z��@���К���T+���l��l��k=x2��葵��$�=+��럜Y�)��^V+!c�H��Y���F�iߺS��S�k%_ځኞ9�g�ˌ���P+zDܾ8We/gS�v�irJ��+� ���Q����2�C��v'� �#&qb�L_���zhm�QVcr����C+���w@�&W䱂�b��vqz��$��-4}R���+ߚ<M�Y��^ �	zb�(�MwŪ���+�T� ˊod4�y��y�u�\�l��ė�0�0�a=`��n���R޳&A�#���Hr9".'����cpܘ��������D��s
D�3FlIV.A��U$X�����W4j�{_���e��N'�1l'�܂�������u�7�P�����\�T�$j��&ؼ*�����,\2D���@Is:w	xs��2Y`&��$Cm3�O�;����L��=��.(��}����\R��0d!2��:b%8o�PN�/���G�Ɉvi"�H�����~Ф�H �"9�k��ƿ[SS�,�e�J�ZUC�Y���xA|�����Q7��8��%.�yR�����-Ȓ�k"�]���g��Q�Ԟ8�&�l�U�(0op2DL�`?�Z�ɥL� M�@�Jp���1�U��Z��X�ǐ����C?'I�n�t$sb--���f�^��S÷5�kB_J���������6�+�k
e������ur�@���Lt~�«@�WO��8�m�:&��1v�ê�����]e;��Z-@;o�m��z���e&Mb�7����m�*�� ]N�Hm=�����WѼ�eu�25 ��U��[��-�YT���n�_�У�T_y�9*�D�p�J��vMFF��%a�|(��_,��P/x����	!E��ڰv>eWC 0"�9|Y=}6F�����|y�p�S]ZEC�E}E�;@v�w��ۨQ-����s�'��oAw}���RX���SEH�b#e`x��3�ԛL|����Z����b���?jLO�GS��U�B�7
��E�z�<�<����0g�|�K�
�Ƌ��%������o�y���˂Sw6J�����_�:�'���8�-�"�1�� ����	�n$);a�I\L�Y��?��X%{=
����"r5���4�1߰$�<��y"Kv���e_��d�����s
�<ט��������^&ێ�~���fK=���s�V|?n]_1�Q�e�<6��?^��N�e���g���:�6 Pt�R��R<�3�q�eZ?/�����&z�����6�(�g{~��V59ZPO�����`#?4��Y��Uz5�@���7˅r����w�mj��+ɨ��+�C5�')~M��/��'\��*��2B���������-Z/h���xj)A�������C��YW*G�B�ߦaP�A�����%`7l�����RS�<z0:�E�x�.�&���/�]ɳ�A�����$>v�Du��c� �Juh�W���'� 3.]r)��7�G�'�/�I�!x�8Nk}��"~��A�^j��y��Y��g`�E��m۩!:#҂tn䒁�e�����V�6�d��!e���o����phfK`������n*��*�<�ͦ�C��ڏW�]�x�b��FkY�T���L���!�\p}���W���E(9��d��i��5�m�n�xM�������[ay%���8�c`,�w����G}����YP�&lG�l)�A!8_���w��oR��p���bM�@g,4�7�-��W���������x��!���x$:��j��{��6lN&񁟀�ǀ��2�������l7��� ��׬�;��{���]����d��7c 3;G��JVaL@�)���5A` 2.p�e�Ӡaq�@8I̪��%l��3E�����[�݀H6O��c�p@m�z�VÎ����
��4���T)����L�s�mܺf�kyYoa�r1R��������[���|v+%� tn�{�A��t�=�]��-���+1�W�����E�o"�_h��!����HmŢ6������i)��<��]�:�2��E���%�/�:���KA.^��x{���[���uķ;m]�x ��fg]�.@$7#)��(��	 	�����i���u��³���]9iIS��1�rj�);��{U)�n�hĎ��8�;�>�>�p��3c���/ɦ��Qx8�
�^�#g3�-SUL��:Rz�����ݜ��(�g%X-I�y�J��0�v��2E>U���qx �Y�B�x#�C�� c�HQ�5/�y�q�"D���EXZR�`�*�(ymY�&!JY}���`{�.�T����^��m�G��P���J�G�ޏ�Y�o�A�~��|�Y�AaT�H���+Z�1"�(f"!���2K�0
� A�z�[bF�j���(
5pr慗��w\��Y�J|� ���E-�[R���a�[̈́��G�VP�4�V���(�h�oPV���SJmꔅ�k��` ���[�T�ӫħ��+\A��l �0�[��Z9ژ�'�Cw��yeUE�P�����%�ʪ��t�e�kKD@�A\���&�e�҈8�6�I�9BCȕ���XI��t����a�����ې�`�±Cj*�>��m�"iW���IF~��j珪��%K�0M�:���#׻���<(�|��.�t>(�}TV�_l�}qr�`���e��Zw}�S �s��펠�q�֭�a�x�ݼ��H���k=�^��*`ޣ��'C�UkC��������	Ü�:h�Hu��OdG��#(���%��DY�`��ќ�D�[>l^ܹΫ�̀Q��I�m-�}'4+�����֔bq�W@���+|���"�\�����v���bk��7zX���q�sd�1ٍa�R����v�����|���2�0,�r~�Z$'Ms�{�ۺ�->���`�����`�k����!����Ս:��JY�Ő���S�O�>��u���ҍ�)��t!d���p�F�F/DVK��5`��N�a%��&�c�A=K	0��I��Ĕvg�O�`44VoH�)��wm��9���<ps�4�M�?��§:� K}�Hp��Nk�[LC��!�R��$�? �R�d0?�n,�*��bѤ���t7_��M}{K����|���9�nAet71c!S��������ƍ�}~��<l�$�]f̎əw�I���0J'X�P�N�|	��f�\U:P.���5R@�|c��WL�\�j�L��  �V�@/��MPva�w�dq-�U������|�+���C��<l�FJ'��^��F2�\0#DZ�3�]����Y�Hq �U�b͔q4/'�� ~��v�6{��ߚe ���Ğ�-�=��&rU�Yi�V�3L"��*�Di�ɨ��tJ�"�o�,W����*�I8/��U�;��O=��� ����FLԓ\el��v�F�fo�e����I�'!L��7g�Ʉ��������=��:��u�̐����6�W��U�<&��p���&FpA! [*�Ae)�>vŠ_d�'�:��U/�����#�؆�yF���A�у������8��U�;5�O��,�R��e馹XC�;��,�Ztd�wx�~�X�Sk�)��X��K(�O�ɞ�M�_���^#�����WK4���Ә��Ě:�ȵ����V�"�`��0fH8��FH�n���QPλ�0☟n�����Z�۟��~v����k��x� �f�gA�q$�I��?]p���,O>=R��>N�ZO���Fbn�DqCrG���Ɂ!�b;.eX9��*��j��F���+�='�HA�u2v�WA�f�ziY١���϶���;��;<5����\MS<��q�q�)�_�����;?��YK"e*S|��~��5���aO����Q<g����!k�4	�\ ��n �Sv�AMx���X�j���d�� :>��U������p�?w·��dNW.�A�b7%�n��
���~�f^R�G�k|"Tw4��6�%%qY��'w�.�7d�!�&�r3+�{Y�Q����kb�PX�R���T�_��~�}(�(;����?�c�ML��f��ot�Rݵ�������ӭ]l��
�j���x��M��w��GM9qR�ѽ�ZȜ�$��ESm�MmY�\�ے~*r���#�r>�&G�e��b¯��l�>�H�N��R�z,�8����s$u�7#�����d��U��jc�W�t̀
I��X�fw-�^��5@�4�A)��Ql
M=�$��J�*�$|u�V|�����)q�v%������k���L���_V�h�$G̶~�oe�a�U��L�j�B�M�����Rz\��1�����u]"�D��k"�3d3,TT���"���|��ߖ�G\D�mý��*ò:���ξVp���7I���]K &]�/��2�ދ+��E�A��t0��S��=�Ja�5��R?Y�����Smt0���I�_8Q��|=�_A�2C�1�.�b�@�����i�'2I^n��S�^hE6JM���"'̮�c�㦜�P��,~܇E2�䊽)�����Q����o��%��^Ce=��@��|L�r��H�
��l�[I��X��O9�Z���68v-A����,�\�9(w�^��~٪��߃�vr��1+��dz�5������TK���Q��������v�&/���U_���9�J�nư�Ϙ���@u�&�Cх!)7��`���#�J{H��b�3oM��'MGZ�,�&z`�x�[,��b�B�,Uާ$_�%��O�k_�B�������H�P��2��j.)»�5�R+�*�z��H��\�b����:���4#�"�ɦ�՗0wd�vhCw�N�G�g#G�X�m���%s%�С._��e��(&��f���""�/���G��(��W=θ,x�lKސs�l�������w��v?.]_�5��S�.�9
+���֭�PƊ�L��_Qַfy���b��)a�n�7��Ρ?f��D�(��%�M�4KR���j�v�4n��9���3zj�1o�-�єA��Ÿ�'_���S���ηH Rw�m���*�h�]5��)f��,�.}q����/�B�>��`F�.�;'�+g'��V�����͈��	��������2]kb��LÖr͟w(@�{�;��BZќ�Y͝"/��s{��"�R�����r+Q�>�K ���.?G�E���eb�Ґ��W�]?S�a�����X���i*fT�ms�Y�N�1x�M��}�M��0�'���*�����
m��创��j��l�����At#���!ܛ��m�>��:K5����S^$��%
�zO���|��J(B;lQj�bd��s�h�����"ܲ�IH��C^l�^�xTz�`�P�������1z+uػ0��d��Ĉ�r�8�{OɎ[vma�^`pр,H�IMt�x���h�#Ǜ�ĕqȍ���9�LHx�Y��*��l���ԃ˫����I�üq_�*�6���M;��cYGt3?惲�(��a��/ʽڄ�,��j���Z��c���q�I�:}�I�����3�������66i����`���.8D�㧃��5�2"��MPp�r쟩�0����I�҃�'��0�m	3����;7�R�c30�#��ɼ�ȥ����F�K��W��h���ü�^�a�(�}�A*�Q뮗�m��W#ɻ�q���rB�?f�Q�I�>�b�jH�������M-�5$T�!VIp'jK��v�yրSJ"�9����q�`6f��l>逝9U.9��h�׺h.�{�6%}�#�o	Dk�S�1��¹�	}je����:7���8eh��0�O�U2���������@=�^�er��~T�����+���Tt�p�M�_�V�@&x,xN��h���υ�B�¹��ݰd��O�@3&�U7k}���9N��Njn�A¸?���� ����{��/�%���࿐Gl�	Gڈ�A[C�>�>ͨ�e hS�g)���x��Q���C�9,�(<��]{�.�����R�?)Y�
�~�ŧ���1+</�㊎�[�G�|�M&�5�{/%y6�H���k�l�.E���8p��,G�`���N�G������Tx��R�����HL�m�$n���Y���=G�t���Z��E[�_��s��U�㙭Z�"�Ϭ���9��Tc^�)Q�]0��]��љ�i/��S{��$�7�zex��0�컿Ev1辷H�	�u�P� �C�'E��x%�Z�(lϞ��[�_�꘳�����Vx��(_bw�,�[��թ�9g��剹W��reO�ar}5�9��[Zi�T�W����dHl��5����ݏ̻5/���C=��b&W��������4_���}��߾;���|ƀ����t$� �� 4ͫ��WX�2�[s/8'��E��m�6P�H%�ŋ.l�w(��X<B|�Ӿ��ì��j�<�˩�H7���b�~�cޔ3X5���$��i��9�ڨ�"�� ���}/P�3�l��DUQ [���l����U-{����GҚK�D4�#r2�+]f��� D�]$n���qg�\�ܪ!�q�]~����d�����vʹ��8���9�F�X1/�)"G�8��C�����r��Z�考cӞ>�P�fWϪ�/{�`���(�-,��4K��(���YE�_�!�#�#��ӫCr8�'��"-��c�q@���*��V�����pp���\`��\5������щ���8�z�2#�
�´�Y�ŢHVO߻BS;xN��%S"�5�jy4�I�DO�E��ީ�'c�Ux����2 Zr��8F=�I��{�P�^���R������R�j9���YuY���#�͜�G�Aꗚ�.�$���i(�k˽ܥaE����� Nd��~�^�}��r��g�3���(��3;M[�f)��RaH����q4�3H��}+~
=�p�/撓�狓�:�	!jl��E^+��r�+�.Q$��6��i癤bd2V2N��y�}��7�Β�w<��i�W#R�U��+j�T-?�=m���஦������~���tZY:�ν1Bd+��]I��e
`�q~���l�ݖC!��Tb��L�nڶпH������:�*I�w�4�G����}�m�:�
μ��R:�2�=�SY)?��,Ժt	�-'ߥF�h��Ʃ�S��9�[ ��I|���pp
�̣O���t���������v�.�[i'\2�� CٍS�Ɋ(�^��ŧCK�������X^�'v�;�,�C�{��.�)�K�%}��zX<�Ċ���螺$��Dp��OW�#W"Q̍����+g��r��S�	���0{�Ab���%5�i���*�N���/] ����K��l�-$�����8�/4�m$N)�$J�G����,�������)}բ������P�!��	�	ﯳ�'�n�DL������%����3O,�o
��ʀ&�����ʻ ���6��)���x������-����K�įhn��,������C��-ߺHD��s[T��Ɔ��VE��?5����u,��d4'��7Bt���ݿQZ,v��X�&���A3M�˛���S��nY'Fk��h.Oy
5ʗ��{�&�0�Z��Iy�A۸��|�=TH|���!3/T;)���T�0�a�~]5��g��0��8�ʬ��C�X�)(`�;�a���I�^�j�!���>�E`���jEK�Dj[^�{ǾR�	𜢪-}�i~�{3Z#��m��.�*��-҂f�R=���AxI.�%�=���8*����d�����w��z"��B�Z�a7�&��S7���>{�Ԏή\��C	�����Mx@j�vr�,�T�}�}40�]L�]d���6߼!����-�ǻh��,)kȬ���y;z:�!B�����`�/]��(_��������[n8j2O\`8�ee2n���<5�6f,�I��8��3�5QT�բ��p���au*�]�LQ��MU�*�߮AQ<}DY,�y�.s����T۴3-b�����Il�F:�mZE�ăͯ�SzD"�,�/��;k��c�n��S�@/|�΂����I �������[NU��kt��+s��9��әO��y�q�8g.�N^d���к� A55�i4�[�~��>��j�ZR�Y>J�wn�k�(�K �D��	!�u,�jiS�IX��D*��'��趞���$�4�4��EeD���R�^`ȳ��(���\{/	�]&!���v�u������T�5�'�F�v,Pl1� R�Q�^,�_BJ����d�A����W�w�-|uQ���>y-������ә�:BlW�(Stt�y�L��"�Kc�1�l�d�����	1Z� b�̓x�"��T垖��\gS��݆f��	�U�B����PD���C�;p�����l�  ��0t}��U���Ù�6�ʞ�e�z�|Z/#�e�˶N�s�;.8?���v`	��z���b�I��k)�g�����S�di/��Eنb7�$��16o��|��'��Qw�em���<D�b!C���]l{'2qג�y�i/�{jHB�����q�g��ґ��E�R'A}��K��V�f��ds!�:�]��vs��S!��CԼ��t"��M�cȠ�1�@aa���.g�[�_w_},o�M([�
@Xq�5����I>o� 2X떔����嗴�
z�!p��e�`�G�j�a�
pG m4���.Q�����ڌ�=�� �Ǌ�u!�,o�uQdU��&���C:e'[������M{���BQ{=M��nl^�Xe�K`+���	\Wi/�>l�ip]���	8�%�u2������d�t���D���䰐�������6�ϩ׼�� �7MŔ�g1\~ces��=J�����o�k�|��KG�]�^��zI�޼����gUz����v�=��N�{ۑ� Y�:�vU~-ce>��G��X��8�}7������{����cH[4��+�i�fC;v�R\��f��H��x�J��u�T�����+�3�̫���Wd7�&�[-������w��R���и����^R�n��I-�g�Px7���2�г F;���s��y^\#��KJ��?E�)T��	?�^���|-.S��v�_��M�g�1.��
�K}�(��D�{zcʳ��u��n�1Dn6�x'~2O��Xn�\�9����į���>�S�{P+%y�L�~�D��q�}4>�H���f@���64���յS*���JB= �jJ���J ��-�&U�)A`n��D����'�]�öo߼s�MX��Х;�8�~HpMh���ѕh�28�i�6�g����Æ��J����׋4ȴ����<꘵�hV��ɼ�S�X�	rC�Fh\q�F�a�H-!;9Ju�Da	G�_���oR�|2�����4>���m@��gM+��3�#�P-���)Yr�ɔ�&�֥�u��ҙM�00H�����[� #O��z��V�{ŏ���R�>��˻ᾅ���/�����,MuKIZA�.ܾb!I�G���xͺ����k����s�3�����Ӻ�,LV�q�ǽt��1�K�O��`+w%Ľ���*�؆)�b����򲄥 ���0@Hw���.:���a��5�}p��cD��)��t���:,��ՇFZ�k�� �ˈ��>��+���ˏH�b���Y��v+
�i��N�u��w�� *,��X,3�����8&��?+���;�gm��%j��oY�$�KΡ���Ȣ~�U�C0�̏8$䓹����\��Q��V��/��w�v:�+��]b]p�v]�������c��dĵ~���DGh��=IN6�=N{���¢6�9����P�W�k"�O�.�"��8Np�1��L�zV|d:C���W�H�e ���]^Y�9�~!�5�{������2��W�`_��d ��<:^ygU���h��%����/:�eg���W}���tCJ�R%�
�R��lȌ!b�;�y�z;Û*��;��<�,�g�{���M��<�r?�W=I�Y>����al������!g~!�{@ZI�ZL>�2օ ��Xfp9�c�T!Ey�X�Z|��!�N)��.��=`C�𝧫�����-͝>h$�B��+s�X�mԱ=G�kuI�n1�����ͯ��	P�wm[�v�H (���ꬢ��3]�k���,�����<p- �J�4��"lS�({�=2����w����Q,{����Ɯ�|���j�j��'�YӼ.�-�w�'p�>�΋��؇8f,�9����X*ߕ�(�hv)��I"v{>h�y9(_��ބ�cXf�r&�ܻ��� �74����mA�7�kF�$4���jNw�[}c�Q��wIU��TUb�hO��W2�k�@�S��l��$b%
4���w��?���4�6�cG�W(�K{�k��_z�nD$��dZ�{ĝ���̪	���vJ��P>��ʵ�x�k^�7��Z��A��$��3�%�:X���G��!������ަ��B����ң��u���Q�H�RsU�B�ZQ�������G�v�#�fX{ ��&��-��O�t�s0���l�H����#=�	������w_<�H:���Ζ�v����G�ye��j�=:w�n<�@#�DR}��ߘ���E�]��h��4�3*�E��e�^�z�X���G�tw�O�8+-7h ly�Tܔ{�`��BH�?��q�d�%�29S-��I#���@�nJ%�)�i�[
L��=J���@e�����x�y�����J�	��������A�"�v�o.DZ�����׋�� �����v[�ݘ���9BTǷ����m���(A��_�����S`�D����~�%l���f��5p4�+��������� ���'��ƙ��`ˇ��}K|��Ӽ�h�˃��&����w0���
�Q�������^�8V b�A�̐�#��/I�̘=6Տ�����#�<�'l�gɗ;�R�U��=���<��g1KA�+��)�]6GԿ`n�:���"T67�0b��m��������:���	eq:\�+<c�&D�xf�5 ����f�̆E�#U��|œ��]XqJo\f:�6k��	���C�1��vG�Ua!j�g�,]������)y�*�)�GW�ߜޖ�7���Գ�ɦL� GKѭ�C
��G�SA��,�$qL-|�L-%���9�?��<:J�`����H���[�c�'ꉑ<{Q�D�2p�	�T��.o�����"AGXh{'/�ޤq���vE�#~_���%�o�Q+��Ob<��CV92^c��j�tF��wN ��TD|�R)	���*y�҉��p�μ�8�oiA�)�f���a!c�Qlzx��VY����	#�ۉ�%���k��l����󀟀��u��bGk�A�Zm6|��f~���yJ+˔툩pX��Y�����\�W�7��RX��Ky|�����W=���"����]��d�D���>n;��dP�mk��9Y5|8��uWr�!C��z��3@C�^��˛��=݀Y��2e��T��H>8�Xb��`�WO��� �W;�}f㎤*PB�����6N{��ri�zrs�_�2Y`�&�~d&�]�s�K��w��bak��������Kg�	'(���;G.�$�}S+����qq���\������������+s,z���f|�TLL-��[�|��j@k���(��Tl���Z�F���}P���K��o�_[�d�#���qB*CI�I�Q5��ɚ篠1�}�ܭK]����I��,Br@�Q9�r=6�����<6 ��"A��|�����j�?`ty��ʤ�ϵ�)qGG�`'p����#\��07��ɗ[�;Z����&��bl�uQ��]�V�6�u�1*7]��4�=x�>�ΈG�\���A�B����p�>պg���q��<����Ĥ��Q�)��2���3���_��~U]�)lr��dW�^П��Qsϟ2��k�	�.���^K5)�PE�+D�6�[G��	�"�sj���"�J��H)(;��A���,
�ڣ\����R{���Q� �AY��}�'z"����Zh����?<n2_��c��b���J!��]�i��u�d�uyW�4��q�x�<W��D�N
�@�C�?E��5��R�q�E>Z}H��\j���L �(��;b�V�֐;�ئ���]�Ŋ���R 6��GW�xڢ-R�R��2#	W?�AҎ4�P���J�Ft�茫��ta�����H��>��P�f�;`���l�Ж������o\ކu#��9U��K���`X��W�8��}��ؐ�j`��Uf��ƈ)���7X��㸮>cx���"�*���[$��J��Vo���\|�6�ch�������� CW2DubWb[�$��1�<hT���ow9���+��g����"x�i8�W_t���������Ş��14@EJ9��=Q��Ua�n?z�����ܥ��/7��5���ДZ�1���Y����R�%�%��%zݷx?%g�T�ݓ�E�W�>�X�(X��K�R5����s�
F|�/�&n�7��}Ȉ�ze��T��'�GL�ߖI@�Xq���	�q�pٷ����?c�	���{C����﵁�0���Y�5_p&�OH�/��p�1��h��,���/;���m)�;�*��m?�3����:u/�"�����{�|�z�ꈋE}6<'(��ڽ!��Ie�����Q����w{#�ͬ�Z�~�^�j��Y	R���ڙ|B�s�of��#�}$�w)���;���|��\B�#�j@�w=Rc]����
�
;�
��g���H�-\Zs_�
�.��򧘽���y�������#,�Q:	a�˵� �<��_ʻR7�FVAt��N,����Uz�br��V�g&hԎ�"W��O	���&ڃ��:>�q�n!�>������`,��$�yV�.4��k�5Y��"2��ã�w;�z��Ĵ@ַMZ46`�7Nx����%�m��${4:�Z��w�)�ވ�<�<��0)2dr���ܯh��݂5P�i�3�Გ�h���7K2�[�!�����!0�P���QrX^x74�2V��(ӊLA�f��) &�G\�i�Y�W&�4*p>f�"k�)%\�8o��M�T�2��w��x$%���x�����yee�wP��H�Wy�|��l�����FR?��<?��(U�PM�.��g~��@j��-�f���j��T·"��ICc/>D���@��/���ɵ�\��r��&�PJ1[��d��%@U�}�hz�����p�[+t�~��(�G�{�����X��O�Ԕ�@�11y����������!e�_���5��&g�&�CH�E��"�:�r%���w�mA�Rh�|��8���'���	9���i_���=m�
<����:t_�<𴓴Aư8y*�|	��Zd;(�����r%�k1�`<=�n|C� �{,ol�Q׿I>��V";q�cM��Ԃb�u�0��u���\Qg�
�����"�����2)>&G�{���V���Q�BS�Zt�N߬T��G��B�)'�����SK�X��m�����6�G �G�Y�P!G=0^3	T<��w�C��'��/ߋ�i�l�46��U �K9;KU3*Ԋ�ѷ��贋^, �L�Bo���9����|-��$R�Z�%�pzzR������Z��:��"��C�@J������\:��a%P�[�����:.r��	v0�^.�Pjބ�t.լ�rt�fe�啻�iy���O�)�%��b����Wh�<�l��͹]E5 `��?�tV�_H�}���9�W���/�&���@�����g;���gQh��<|�WC"�g@}���`��k��[��(���|'�����0Df����s�4/�U��C|�����5eP�.Ā2���+�`��@��J:nE.qt��t��3�~��G7ðH�0���OMfJ���UJ2��n��&�C<U_�n���aI>7A,�i� ��$��͓�C��i��C�
�/�)��s��j��EYE-w��A�`ۿ��ZVܿ���
9�熍��=!7�6�F��Q|�G�h�0_6��<�_�i7^���>��E��.��1�Lm�����V�c�y�U�u>z�ԃ�w� �	�y�0��]�nj����]0r�����H>�C`�Bi��-�B~O��� /�ftW����#�)^HOD���9�<R�_�����EUÞ�X�|��F�0m�vGǉ*.�3�σ�V�\�������G�8������-��4*�z<\�}��a��6�قB�[�ErwZ�(�/��MS~2��ٱ�C��!>�Ķ�FS�c��/#��ym���_����଒�C�
*�a [�ܩH1e�H�V�)<ɒ/�`�>��mg������e�}u�Q]h�c��N�0ق�ֵ��wA�nX}`�<�Sa�RPC���7�H���ǂ�M�T���1�m��_.��Gca��4��MHB�P_0��N��H�"C8B?V�ׁ(Y�����Ӆ�-s���y$���A��vټ=�.@�a��d��hs�����ȬLu�ێ��,E����є�R��bT�	��6x�-��\��.|4�����������XWݰ��@�1�����M^�]�%���Jǁfn�@{ T��������%N\6������5�n�j�k�M��l?�O�\�*���/�������ȍ5���aV���me<8�Y�L�
�"�j}r��/�mټ2FQ
dar��6Ӊ(o�ĸ�������1uyUw|&���y)屰4C~2�l��qƅ�\7��8o�9LD�N5��ܰ3Zn��e�bs��-Դ��x��o(~�82��߂�	ۣ?X��r�gX�:Q���jlb�r͵<|���}��4l6R[�<V�*�Z
s��(��/bYr(�s�a�w�U�8&F-�Z���̋@�D��WL���<� ]H]a�W���^1�P��Tq ��H�0�7�����!4�B���!4�=���-gj�� �).�^B�T�����=���®q�Bs�L}U8�aB�Y1�< �����>4:����6�{��Bj����Nz����5>m�Ϝh+8��<Z��m%��Q��5�'D�wC`�&}3X[1�������L��Ȕ�o�B/p�n-��C@�L��-� Ϣ��_ߦ=��t?9b󒫋�/�	���k+9 ���f�j�Ue�0�C!2(ݢ�(�vV����mY�"6�5k��P7�淽�(H�qU�{���}42~��P���V�j���g�tÊBM�%P8�ս��y'h{�I�+jf1O؅\�t/��rue!;�W(6���ԡ5�e�W�맕�e��P�)�Q_.�6�S��#c�kS�yWؼ�+��sA�j"�f���4w�
��A�r�5�UwH8V��T	�{�Ij�d���4��:��������gFT��Ǵ��X��vC)�R�&!�Ҽ�)�5���Þ��c0�j&�o1���i�\M qaa�bq�a�����G%!��A�Dk��˷�H������C,�!@�! �l�#�@[=�����7A��S�o�gS0AW����`c�!dU'ϮL�j�ܸ����}*����.�J.)]���!H�-��Hf<c�� �g��l:`��mE����t�t�K�u9V�X��5ɕ>U�:�*��łC$��<ŵ��ԇ���0[�5���6��<�LD���	�Z���j]rT\�1:��b��U>�}Q�ʤ\
�O�\�oٻ�F���JI�E`��vj"��노,�[8�B֫*�ZC�e� ������f��u�3oR�B�U��K��K%������*�.m� %�شUXX��t�
h��.`P�2���׌JMB�yy?M��a.{���4&��}H���?�]o�ka?�^>b2���"�l��!>��lA�֌�$�Ӵ���щ��vU�V!�^��3	��঒����b+Z�]éy0��c�����<��#%����E��3*,U�V�Q?i��\�Ŕ
LGx�&U��v�1�i���s�[D����y�bv�Ƚ������x��y7 \7��Z
���֡�M	<��:� �r���IQ)q�QοM���M��\WM�j?s�/�mb_ӣ�1`,,n�|ǂ���C�+1C���-���]-���������sQ�R%�� h">6�
S����5Ǘ��Z@�3��C8e��T�u����R	+a�):��VuJ�t��@	S^X��n����&7���ե7�֚�9�lN�n-OȘ���������򒃩։�[�D�&�襟�J�
������*P����د��YR�k/Tv	�Y,�LDM�}���A����;z@�����L��y�c@Y��В�["aß �RS;�N�3��u|��C]Ʈ3d)�@m��03�>�Ȧ�O1k����$UF6dZ�d^�һ��I��hT=��;���J�%���&T�-�B��a�-9P���=X7t��/�3)GI���I��rQ5,lLL�#�����/�.���� �r9f�����˜�\h�ּ�p=�v�㟣��e<��6'r����*�F����[���tS:�Fځ��g�56t�)�sB Q<�Fa��#:�l~�ڽ-�|O���,_��~C�䧋�o-&=B/�0�hA ����{�6jr��xhε�m4wy��.���'i�0v�Uk��-�&�Z��`[��F5���?S��\�b�n,y����k���[؂b�R6x�wٗ�"����Ջ-)���{�|�f��wm]���%E$�_̥(/�x�$��p�ۧi�s�S��ʹxz,���h�Fe�q�z7���-=��e@'�b�<�a�F ʹ9h*U��l��Js�,�@��)�G�� �k�/����WieN#u��02���u=�lw��?1c���F�,I��}�}�v������JN��y^���"���-�
3ux�� �#t������L9.�� ���a�j�C�~�
?	��H��Q��X�8��cjF��I�R���q��@c@��GU�����?z!��ޑѯ��Ę��*zXs����$L�0k}VSwN� V�� �f�V�����jcq=&sI
�����>MB��q:��0VI��m��z����I�o�T>ܙ��cƪ���
g��H�L�����0Iq�;��͏�Y��mU	�����Y!����^5ȯ#�j�Iq����N����X�����h��ᆅd�RܐX�oq@ļ��-��q��Fx�N���:wF�bA��u��^�	��(p�(�5;d�����:A"��_#��jk9��؋Y˽�u�Sea+̘w�B�)������������=``�<	p�/O�$<yñ�ߐ(�m���W�A���5 �� yM���aiZ��w�Nn%�d�K�M��oܖ��P�;ڣpDHM���v�����$�"1��9$��}��M�9ׅ�bn�ߔ�6E�oi�rLo�U����/�VW���-��1�ۑ��W%����Jٝ?���"#��b D{�L�(�ݥ�O��r-��^� -.�W�/_�ic���lSn�"�83��zJW!�����1ƣq_{��uR"5R��͊�X�f����5��)G$!�x{2�K��g�1	-R�'ɋ��� ���#Jbe6�b�	�f��� ����B��{n1qn���qK_W�8����yů*Ua��~qfL>�eg�r�=J�D>��,�7Ӿ>��A��u��m$ �|��T�9?V�`(�C�R�_|D �!v����� �ZJ�Ik�&�����GF�F�ŖAx9)�G��S�@�e{���rT��S㝖�����/	|���X|6#� �;*B۵��)C�'{S B��Q!r~�la��1[�rK�Dʀ�� �I�t_���w�h�W+8��ϖzKy��'��h�%gj\�Ps��~u	\i�2/�z}B�䴍���j$���%���U���2C�v�h 8���V-�H��7�T�=�29J�o�� �䵯I�:���*�2D\P�a&j�ZT��A[��}����<'�}-��瞁<�����M�����El�Y���dś����$�@\J��z�������-ët�g	���[�[h"~��0��k��,����{�l��6���.����O"��ao��j8tw���̠ߵ�)1\
8�.m��p>�)9' e�4LpA��=���X���
>1O�I�:7(�}3$��/�6��՚o��1�gBώ�ڑ�A�%"�1�i֖j?��53t�а���-���V
Ǘe���T�Q-�����?����[��w�R)j~2zl�Y�R�y�#l�����
�p۽�y��ˈgWڽS�ʥ����W������Cs��ɩ�Ġ]i��ɴr�߳SI��H��S�zfi�{�g�c�.ڍg��s����oQ���-r�@�[↵/2�`�� ��EKJ�X�$~� ~c�"w������+�K{������H��z�Y��_��|X�D��T��jG��m�LrV��ʆ"h(w�{u4*z��� +��W���S4-eg��nUy#���#�@at#� ��;�Ԟ:�Z���0uZ�߹��*)/uʅ8��먼�3��>_њ��]%�M�V��⁬����F��Q¼��6K�=��f�U�_LG*ŵVhԷ��9������}�\�b/��s��G��%
AD��Y*�hWI�.�&���Q Q$�V{m��FŪϝݵ��Ӕn�)���/�e���<�"͚%��Y8��\�q�L�E��#�]J�w�l�EA�lA�N 6TF�+a�JL�m ��S#l�>
CPn��[�z�P���Z�9\�F_����E����	ҤCbM���ݸxp��垞#Z�|ډ=�π����FP��{@63|崐	���z$ˁB���/�75RD�g��������z�fK,�U�f��#��+�,iۂƎr�[��BX�	��b �(̀L��8��;|�����8L�G����.]��S*t�M
���a63O<�
��_��k�*�?I>�rh���L��A\C&<��V7vb��ߞ�xzη��w�R��Ë=w�qV��A$$3��h�:J:�_�ۄ�����RA�e����;>�Q]9�;M�=I���3�̖%U��Ի*@�R/�R�~^���������ɥv �(�����%(5�8���4���D��>�r�^ǚ�5r��Q�h=�j�Q�ByL���r�w�%T0	�0�v�o��җ��L����3O1b	�uɞ�9�7��#��3j$�Q��&�'���^���+xA�8Z(��ƶ��jX�}���;�3=蛧3�O]���o���[䇍E������̎��d֕^��wy['�R�!Jq���eY��!���eS���q^;䀗���iT��}�ۻ�d�O��k�u�?i4�IL�5�ܕ�5K	��������TU�@#6�x�D��� ]�Hd�u�]�s���w�z,����fH��,�ϦI�\Ih�9�z=8>�Dp���wf��T�!|"�H�5ڳf�
'K�@�<������"V�]� ��.=� ��+�Y�sN�'��6^^sV#L�8���jL��m��b�� l�%��+G"nhg^ՅC������?8��d�j���P�zk�w
��)[Jpk�D�L��NeYvD��IǴ�4S������;Ӆ�r�x�@o5
��������M���� 9'�P���랗��� ��h��J��]�tH6�F���I�Q3jJ��#О�1*��c�\�Z��1�Ų�M<���n�}sR��/�l�/�%�,�w�����orJ��w�ܪ���B�-lF5g�jP��c:-���y���=��k��MϾ3X�@a���ЉN�X��a�w�������㾎�n��	�%����D=s�kˌ���Q]��{�p(��:�n&��ka�]-��:�VJQ0� �C:e�v�at\�w���ж���@ڠ�<?*��\O%�Ʀ�tS/�2l�$}-7�ӄ�W��fy{t_����[vk�������}ϾE,�*�҉��'w8@/���R��?���1#�������>B��}�Q��5"u�CŨ���^�����!����JW[J��-j��N�,Ɍv�ą i���@/rK�-v�B���=��u:Jq0�	kǷ���h�X�X^�����V��\�F��
�^ފEL��h��;(�?�D�\�/�!�i�,���8a�0;&���O�}v0�ٔK�oa �7��$����}�f���/��
�i������A���a�O�2�"����D���Ou��
�U��˰��j�!!�T�✣0��o���텥����W��E��H6|��<`&E"|��o��% `7 ��\{�v�D'�tcg�fZ��=+�0VZ]�Yn�= �m#�?A*h��A?v%�fg,��):hZ��&��a4ޫ�V&�$���ۑ��}�\�������5�'S/��mH���+\�$�����6�B�4��A�E��&���bU52�W�[Z߹`< �e��̺]Py�����m%n��4��I�X�ܦy6T��n����@ՉP�樘�O�ubbL�p<O{�On�FJ؅\���*	�Q"���N���f�|��ɘ4�_.�pz�0�a�5`�ˎ����ۦ�!WMi��ЧEL��2����>��Dz�P^��1��[F��4�N�2�`f:�Sz�17C���m�2�#rz�G��R[�BЊ\��3Ds�'�%��l������L.i_��WS����:$X�l	Mj�5,Q���B�+�LyS�*Pt��(�Ih�þ�|�ł �))�b ��F�n׹2v�W9��.�+�g�´
U�i��s��4S�X奊F}y����	�����,�ɜ��nFī��+�nz	wr_�݁v�,�4�b���!�k,���Ü=)��їk�w����_���n�{ك�ℯ|ЪO
?�H�~uT����/���b,����|%aUHx�R#���_�R9}��J��g/h���VU�>��I>d��&F�2���;I4��1JR.7�4쭏p�J�FGֵ���4��Q	&'ň�0˹�?���;h��T�`)�{	�:d��H*L��ݲn�`�d��N2_
��'�?ÌzH�v3ㅕ��EԕA��Nȟ��؋q�S��7y��z�'Yj�\ļ��w�v!�!f���R�F��G�^����y��_c��x�I�;+	��i�(��A�S��q�:h�D���Y��{#�����Jbg�@���b�.�^ã��yB�}��e��2f�H���ҔN�{RaA�{Ǒ�����nM��!�l:�(�"o��Z:�)�2rbst=���任��l����ĦQ��0�|�#oa7ս�>r���u�%�o���H:�e=/C�eq�-��q#�ۓ�k76"+��PN����m>k�d��Hq[Ġ
{���k�_�i�#W�Xf���ĵ��� P�(ta���ebsc?+�Oyg�KE|��Z�(z�ɵ
��I)��ȯ�{*>ǟbG0�1��@�$�(���fW�<W[Sm���ɗ�������<��]��5��a��4Q^S����a<P�G˃/.����y}���2���b���Z�[�κ�d[Z�̼���~9=7�wg�9¶ܡs1J��[�	ؿ}V�4�m�'#��n9h��:Q������n�#P�L�v^pD �L��U��p�gxp�d�>�$�R��떭B s�올w����$Tw&x"7���I���E�rg��=�W?�	��h��&HN�%�Z<<� �Љ�X�0�Y��W�U~]��B���A��H"��J.��	�(��+���,��-�ciw�L�tw�Nn�W&���!fak]�ǣRI^�`�4�Y-q�c�A"����9w�6.�ȍ
Q-ƙ�ߛ�v�%D+���M���f�|�F��bi�bjmBX,�^�UAg/��r�G�?�rM��z��gq��v�xV}��+��=���*���_�@�-|ѲP����}p�#�#�o�C�t1�-�^V`8٘�	o��AJ����O�'n��<,6��	A���aS��Y��PШ=�� D���UL�Ĺ?Q�P!�wPf_Ғ��Sড়��M"��u���>.H"�5㮄
���7�lz��t��q=y,.� �@]%9�@;�٥�ĠLPh�u�"�J==�nW��k0嵬����`*�Yvn� k�?3�/�����Ͼ�i�+1��(;ꐧ�����UͰg+���9�h���&��0���s���-^���D�[�A�,k/Z]���t�Ǐ �������ՔyS��iBY�{o�^apY0�;�/fy'��H�^��i���8n�QG��K=�4����bŞ�k��ݸ=X����\F�0[��N�0Wn����r}!W�.H�:A�2wѼ�Q��9�|��$�~���N�Z��z�r���p�2G�
� ��L��8L�����xID�?4p@��vh�z��c̀CH0]��{w�4<̲s�!q�R��m�'�:z��F[�\�{�o��J~l؟��`��0�m� a�g�����`Mӄ�D�#���}y��
i��!
��:�.�G13PE��#-���V<��T�|�����~s��f�
��K#��Vx$i�n<Q�1���P���f��{m�Rr2hh��v�9�N�Bz=!��GS�kj�U4�~NmM��Tܭg>�|%!+rk�a��7����[RK��}/ν;G7�ɪ?]��2��M�ug��f�F@r�����d��9[Ve�F�D2�v��z�fy��\�bg�s��w�eY�fL5.�ne"Ŵ^7���UU�����c��Q���]P;_����bhTq���9D��^���Cxq���pN�E �gd������A�F$Ʈ�M����j��*�@1<V޵<�kj)κ�;�;e(����zpK�!�J󡃒��~��Lj	�~&*��$�jU�B�\��g�(UY�5@qa�=��jb�^�<0	���ڀ���f����E�!�����0E'�	���r�3I���<E��&����
씨ƮX��/�K>��c<�ڦO��ypB������hI�Wַ4O���/�Nz݉�,�p�=]TݵR@��	;�jɎY|Xbr�3�@BO��2�y�l�㍋B	�N���I:�ud� ���<q���"�U^��G �[R�H̪#q�%w ���Ғ�4E[�S0��?�;�nq�ˡ��v�p�Y���Q��Edw��V�;q�g\�z��<7{ x[�,sڟ�e���2�����}6�Ë�ե.y�-*�x7?���]v�*�@uY��WSźꙛ��Gs�=���z��#����EF=�*��Ha4
]��r;^ZR=���t���};���''��9U��h3��I�L����y�Rs�\':#�xg�2<������ڧ�~��ji�x��\����֜��.���R�
��<���<fA=�]rTP�Rܕm��W���+���b[����L4��T����j/���>>E,�i�-��:F�U���L<��${s{Q�W�}̓x���D� �jz6����?��R�.<�C��7�r���`@����6��_��d���ՃO=1Q�T���c�M�ك�3f��\OW"�yy�/�n�U!��,V�e	^.k#�xr�����������Ibna��|�l��-�����
�O6�����j��'�*�B��2[�=m󭼠[�a�Ge~�	j������Rh!Nn�n�h��D>���M�ة���qS%��뙩_��p�GŅ����0)��*�:��9y�d(Ӣ&#,�F����3T��i�w\��\.���sh:ƠAr�E��(���a�&6�T��]�U�4ַ"�'�q*���%�Md�U�?�(���];��*�)����b:X$��冓�r�#A�yI+���ʽ��`�����Si$qq
������Q�}�߰�'��+�l��"���&(R���,�}��m�)������|%�j�
�M�#���rXM�V�g��+QQյ�A.`�U~���Z��I$����O�­(6/�p�ҊXoWx�zp.$��#�/#��F	�sW<�Q.|aױ8�z��j�#=]��J��v����1�ӧ�`�uK��4�(�������O~|�:0LCp���{�K�Fl�s�hx�F���a.|uށ���>G�%�<%�S5aZ�J����i�~�֍�ꁞq�����<���W��БU%{�|��w��4dj	�㻟���MՅ�^�A2���9V�i����#A>����4���/������gZ��LqY���'-�A-�*l����D;u����Kd ��)YD׹��S�:5d����+��-E��f���ʈ��(�*�h� �ρF���̋� ��K~Ѥ�Y��L��m�DU�8Ӽd�+�0��,����MW"-}et�_���S(�;	�-�N��#Y23Ϊ//ǞLo����4e]��t�%G�1����v��!������k����<O/��eƣ�{�E]��g��^6(�_����*r�߆����F+\�v@u���~��~x:���]\p�.����" �*�/'���0�JN~�#�Z�]!덿����)��W�$3tH(�,uTO;L� ��r�Q���{X��!`ff���i��7����.|�c �a�H���mV"$�nJ����V�K���D%F�(P�����'b��D����3x��G���W�Mф�8.R�;�A"FI<����	�A��e��^�Q<GR���=?ܺѽe�w��fu �"8���WM����������{:F�����Q��s╨I��KP_�U�}H�N���'��`����Ʌ����d(��o2�;��[O���m��|�J��Z�R��޳e���^ 3J�M�!N{�(�V��@�a�G�#���2�8֊���0��Dz��>�f�E�Y,Ng3���`���w�G�ȓ�E��PfwE��NJ:��|Dπ(��I^��RZc�1���o�7����쥪�Gɣ�.�|I�.�~�dת-æ�*�]�-<�B�"���k]@xU%������~d�#Z��a~�y�}+���Ń���wVфz�ܞ�O�$U��b�V��c6��m{[mnw)�6|�R�����/����:���G+j�{�!*�Z3��KȺك�]�M���U{�WY��pU�?��2�=�g��s����
���VuD�Ν�^��;)�g�Eİ���4�����,jH��S�`�aP�/�c}�/�("�%����x"�l|q�֍�]S�b�.�c-m�#�M��0�t^ķl��Ǉ�0�	&��W�]-4&�$�MB�?�D� ;�E ���.?�`$(ѐQ�ABJ���9n��Tx�<))ѿxۨ�
96A̾G��
��y6�sJ-��/������p�t�p}�d���<��W@����#��}�&>t� �.�b��iw��Ű�p�M_�һ���Q��f�2>I����?{�Rb�s�ٵ�ݔ�|�bȆ3�U`�����t�ƭ 6�o,ʓ�:�?U�:�Lo:�3V_)j,B}|�l�Ӟy7���Vv��W�}[�w= ��"Uy;�ט�z벢�,��[��Y��-����oD��πf�����֭j-i�$-S������qf0-:�n���*����,�uة���nפ�$�4���,27P�$Bb�q�����Z޼Jx졅��6���ˏ���z{X�l�
��aa}����$X\������&d�D��9�M�v8�O&1IK�ź�w�����H^8Y�����2��D3�Yťo�����Z�OM1s��hܓ_z;	R�O�ޝwbĐ$J��e�S�F����QϢ��Rasy���:�正�`q�^���P+.��:�����@'i��X(FnWIӮ3���^�!���%b&$�I����yX#��ȹS˨�-�ޝ�%�&��H�p��|1�ל?�gׄ�d�a���ʱ��l�C��טx�p�6L��i��Ep�k���*7�f�l�
c��a����m��'��R�[�@��t���Џ�f��_\CI@�6C�4&��IŎ�0�Ӕ��ʋ@=0�cU�Y.���s+-A���e������S����1C�Ɠ���#%\8�R�៬�> �~b��H� �{E,մ	�Rq��c5��`.N��������B�=��@f�K���R�^=r��7^�Ͻ!�c��܆
���9��򰋗^]��I���ki��"�ˇU�sZ�o�?s�i�=\�ڧ��D�0�Y]�v�O{��S-��ɫ#6�\�`:d����&N��l:�<(���|�S�G����
w=Y��V���u�)��C����j!�IŗH��5p!��>����>����E�Z`�ڭ?%M�.��e>�"��>�� �Y�K��u�Α�)Tg�E%��zh	2t �6���A瓃���A�#�
1� H��Kg �� >,ok���$ۉ�X�JY�G&�n�Pv���1�� ����+l���o��&S~�(�����X����e�2�V�=Pi�U}2=�ʌ4��=$�k�,k�5F|���ps�%gd%48�09��$(B��d/2�y�;"�ôR�6)ٓ0P%��ȭ �\����Z���2@̵�g���#�'�I����t�s����@�[�t����lE��c���T���a��fC�;��*�E��D��b�?�u�eՍ7q2_AD���~��7��gv��Lv�Z|��(�U��>+�?�"�|��}�oͩ`���.K�����xjN�� K�_��i'=�K��`�;���OA���<�s[���،â_�&���/�s���[@�Z�>2�M8�i�Z��
��:3���P��R6o���X�8�ˁ�0H���J��4I��m��Tw�X��i�m����7�Q�P-��ƴ��&�#M7������!7����o����/-W&7NZ&���+�H�T]ii��{�b��U1����é�zi�'�������v�&�/;O���2�)@��<�cw���D&��fǈ�~a���<7PW�;����T�Wס?v�����"3`+.��g�Q�q��Bu`O�i'Z�Y�k�]<2��IF�n���݇ ��Hs��2�4B����2`�o����#D�WXD�����`�� ��qK��U�nH��PnrH�3Q���K��g.��6hiV8,cR�|_�#��Q�,/�څ�앉�C�P'�>�i��<1hQ�� ��=�6��R��yo��|vT�R>�_6����'b�a���WS������xj2��'�ak��3�r{������&m���d���B��,<���R3E���h���������No�����e�f�p�.�.39�RQ�
��g���V"l¦T<�@8�����*!�A,~���~�r��V�c
7����;\�����y���tI�$�g�jr��.RmCZ���7'NP�F.�0Q�LFC^����A�U�l��r{���
!�N��E�8����^��㯡�y����紆�w_�?�B�C��J���?�tb�pF�y\~s���|Z�T}e�Q�Np?��V�`���>���2 E��.0$�I�ihD�J	���޺FK���,8i��gH('��=���&�֒�l�I��=Sb5�`"�?ٸ���_�)m�_>�g�~
����J�V)Ѿ�4³4!L:'�fZ/��pY�jxߊ�t/`���MIVn.�P,2�sW����~>��x�1�rr��`��k�ͯPv�|��A ��*���>����l)��D(��W�7�T)��@B(FA��&c�����fi�o��ି�ɳ�*���ҏ�v��=��g����c�b��<���W��>�1�vcL�Rq4�S��5������/��Ÿ�6�.�CBv��}@���]4GtO���Q;GM�&4�EfN�������!�u����\P�,��oX��_��SL�t̟�ke���t�f-�:"���7tMs?@^{#l��u,QL$��ߒ��m�k�����Ӵ���;#D������^��R��D��kr�7�\��5I�*��\z��P� ð
���V��B앰�G}��R66'4��R�0̰
#^��\���5ֽv���?��i{N������z0�7(A'��>���1-���9I-5��~�XD�FM���o͏�;�ug'�?og��l@R���.���}:F���Mf�~̥�хHO$EL�\�$:6P��Z��ną�S�n���P�X+�~���ݏ���Z��׼YăT���6�٦���=*n*���Tm~��-���7*��*Gpx$o8�\��ꊘi�7bQ��fʦ3���	p'����I��D�i��6ml���5��0�0�g4�8`>:�yw�+Tﻃ�� T�;X�ဩJ��h�E��xW���CǪ�.�a�v$˶�=<h%���~B�_�ă�]�K{F#�`$^�����ԯ{�#��]��ƙ��td���[
�:q�i�K�t�G���5Ꝋ�h��l������|��2-?gt�V�?3��-|@~h�*V��$�"~�.A=�}x>XUHN�i�GV(�H���O�[�	`?;�L��P�Z��3~�T�Kp�Y��7xx����Y�jFNS
�݉⹛�xYH)�ߔ �����[8�}�9�/CL^@�<~���z�zb$I�y�H��>�C�|{�o���/���Sw��C���������'��K
߉��\u"�����E�����&+�^���mN�Z��L��=P4O#�@�eb�qL?e������oA��b�1�sչ�V�頕_gUx�})C��\��]�MgA�w���T���l:nBqHy)�s5�I�Mh��Y\�%��%.gh%8�hy�+���iF _M}��k�Z�`�Rp�ȑ<�e��4���gk&�t�YC�	�0;����,��2�qzg�.����v�yp4џ��t����k��e�]��/o�dI^���^Kf��#�g(:9N�Sp~�5��~�`�Z��dB�IȦ��ia�;gq"6��\{^�+�`�Ҭ��޽�cw.�ɶ���*D���a#_̹���2QU���&��vp��c�Dw O�v����X�-��sK�ohb�^��F�S�J)��[ٗ�� �Ky��0��U�B�(�47.����a�kH�tU����l���+?q�<��K�C:��B���� 9�3����ƞ,�6�kK-���)��X�I'ذf��</����B^c�d�������a�C��C��-T5�� ������s�^�<	S6��n2�0�/Ϊ�� X 
:�Ò�]M|쾹�'TrM�|������
��T"X�w$L���g?Dc��g�O���[�����2�W]����Qcb 	�I���̊`o��{�1�]'&�˩���XTٷ��(� 6+|P�F�����)��x8܇�,��S�y��j~Y�C��fj�,����U=Nܬ�� $F�zR������)���3	j�z$0$�4�h^�@E\Ze�P(���oC�`����$�u�~%�����>k�^ �Q��3_�e�^��0�,4ḤW�l�]+^v�]�#� �=So�1©Z��H��f��ls�H��&.�4���;z4����~��	�! ��;dj�@p�Ur(h�W�;%;�D³��%��4�e0--F��3)^�3rTPL��j������]���	���j�`���ǇfJ`\V�h��L��^�L�h��k��H�~]���*�D-tT����Rj,ܱ��~(��CpO����Ê����<����J$/�(�mj��FU5=�i�O3�fF>/��:�sU�7ځ�S ��)#]>�)���ī���bY�iV@۝��%G @,��y�LA�_"�vu�(%������|�g��se"������-����	5��c&x�K���'\P�=��Q��>�AN�lMQ$˕n�4���g�^�*���V������ɀ�����"���E�>���q�zs0��㒆�xt�q�?ۺ�� LyC���$�K�AN�>�s�ug�r�I�@x�%�I���CC�ױ֜�i:(�����V^�<S��*=�,�������A�P�.�V���I���@ǝ*6���G'*�Ȃs���WOP~[ �ܞ�Q�}� �C-��t��&����Ǵ]�c��1�é���&#i ��b&�dM�Y��(	��ci'����eu͖ݶE�p�P[��70g���Z��Q�̤_�lrat��O�.!�U�{����7��C0y-��B��1&`��o*��QO
��d�!��_ZA�c���s�3���|\�&�f���b�Ե{�AGǠ?׊��:1!���fK�j2k��^/�x�Pمe�B��p�+�V;ߟ�,�Q�h�����Qד9���8@чW݊>f��a(戟~gԳ⬃�B�Z���Yo��J����c�h�?"J ��܍���V�I��˱�>@�}��2�`O�����c\�b^�<y� �d���|��V[�.���I��dg�ŝ��� �l�9�L(���F\�������U��ƒ|E����H����h]�u��ۃI�7r�[-�@R�$B���1<���.cd�b�}���-ȣ������1{m(^�'��*(C�_��7P�p{��)?����}c�${&�6G-(�.f������ʖ�8�8�O�7Ǚ�Zl���:����V�JQ��}dcڌ��S���Lc	AI��A;n%�{�i8�L���������t!>��0[kH_� �< ���&����0�K�v�e��+�B\�נ{��ԝ��$ô�څ�;C�e�H|�턉�4Y�Z"x6�G�9Pq{ͤ����cD���F��dOpeN>f���贋b���,[���CJ��F�k(Y�dW8<�@Ff�i���:@�wzg�7v7h���>?��M�4ʻ*���c�,��՟b��
�J��nD�C��$(�<���oa������<�����n��t5���a�iV�$>��c֜Zk�i����Y_R<S�C����{{�e�")���ܑ��cƙ��vI5i�3d�q?�(K��Iq�ty�+��cی���	�$C&%g��KAx2<��ح��e�f�����ś���)�D_5m2�a�&[{�[��K��UV�U�U�o�Ѭ"s��M��K�c���B[3c>W�J�O��NM_�=n`�-Dm�Sꏶ����g����2����Z�ѺLʝ�5R)���A��)u��MM���53� 2p�B&�ٽ����t��m� �uk~����]��2���@��E�sfmW(����%#.��t��M����w"�[/��h��`Z�W�/9pω�dd@c`yKY'
X��Q��:V̽������{l���A��3��T���&���8�,q;�	��ǱjCxp�����~��eS�ٌ��=7��kVmW?��*\!)��h��'�\�es�q`WL5���ɚ}����bv��:=�M#��\�&I����)��I��}k A�f��J�܍ S=�����=��6�Q�8�5�N�ǖk�l0�A����f1���꾋;���������u�;��kVmG���X�Y���ת����x�KE����x-A�XB�G� �A0�w����,kΡw6'̦���ӫ�b�DT��堃��7��y`��+R�L��o�c�s�g9���ŘS9�. �-.��~!�0��f��v�\f�9裶��N�6��_z�a]bg۾9����W�d<a�m�iWOl����ra����k��>�����9�A'�j�#�mj��X����@��Yݞ ��+�O{���d	��)(�Ν�Ig�DP&&�A�t@:-�OR�tYM����x�Uj]��u:N�G���A�	�%����LL`P.���R��#��̷���G�*�g�U�ʻ{��c��^�Ux@ߘJ���A�m��U�pvB�~��dA��څS�λ˺:�5}vm'��H�S�k��3�<g!-�Zi���X�DI^���"��8y}�ښM$�Z�S8hX�OZms1���.��lM��+J<I|��L�p..�,�DT#���c�J5`-��� �u�L�g)s%v�X0���p��碽ªH�4�r �!�ۢaKe�� 
�l����K�������n�rEf�@vKD�>ˆ~�v~����Cb0�K��(��;��4B�����y-BA3�S�� 5�k�6�',ݶ�
m\�"��
�YQR�!m�?Ns�lu� J�?BB �:�36�Y��+F�]��ņ$tH�w"f�v.zLz>���]5`�t��V��D���d��Z�[ ����S�O)�vp�$��G�'?ά�9w0�J��b��/��Ө��E3swg\^f(̗�"i�l��W��pN�绕��W0�[MM5�o�y;D"�ۆH� ���.�-��Z/\�z���1ȡ>�CV�j��Zݩ$<���!�e>}_Њ|5����d~���w�G#\�;|ڗ��ab/+�K9ʎ6��\̃���B�@;��7��#�g�8ܢ���ǣQ���(�8��اQ���n�3\��G�u^��2�-�2��̺������W�+殩{��'�6r���єe^�o�3~�ؓӥ�v=�&l���zZ,F2E��-"D��-P먧(PlQY�-<��1ɐ�M�/�R��>+c�'E��"aB �JI���+��-!�� �L0Z���S s�2fR�}�W��Pz
��p6�10�q�9F6����L@b��ҔI�C@�����{|X[�*����O�@���I1� νc\!�T\{�)/�L��|Qryu]��as�����t�Vɞx$Q�ꊲ��ѐ5�y�*X8C�S0��u�i��aM�q�ׄw��`����6|:`3��`��1��vZ�6�ي��_�E�jXX�@�2�ݳ7|���hkhW�C��R_�IHMC��h�9\��@�-�*g�i��Z�l�A?&G��<�BQ�]SmHM�c�M�0Z��_�]�6��������Z��d=��}��q��Dk�ݢ$�F`^	Hr��rL/qytl�|ߓQ� uP����.��8�p8�\��$���q��E�N��s��\�)ImR���������9�r�jy�O�F� o�66ʖz�;��+��$�%�4�g�Іi����>.��<α ��]��#=�s���p�Pۭkx���d�d�1�
��=�����҉C�\5�Tl����]�� D-)�)]5���H,���@�Q���u��dOM��-_L���NY]�/�er�#��c>7��?!�����V�dWg9NJ1�f/���5�~π�Xk
�Q���
��tZimf����=-��!�,
�=x�K�3�܅�T�]h���'v8��m^\�be��=�=	�{��}��z�O�ak(�ó�ޢ��h@רҜ+�F���g��!c���P�VY\�Oᯆ��I�*��W�rmԺJg�x7%S����z�$�[��҄r�0������r��Y�5A��*h�`s �^<-�6AQ���Y����r�OZ���ⰍJ��`ǫ��A�/��g�45��93P��V���|��*�s) i��X[�}��X�w���{���Yn}����3ͫ�lBU�2z�p�d�5��(�IZ��.�f�9 v�Li�� �`πZ�EE�Ӈ���2x�9��̈#ь�9)$��QJ��8�'sE$���1�������_�JS[k��n��L�R�'�ӼC0�v<��Q��cڨn-��x�;�mP�����q�<nǅ'���~����9����@{��,^�����Xl�q�}$ۮ%/���9n�{QԴ΃�(d��W���h�8DI�n�=D��(
Z�Wm��tŋ��$x����7�m�:��bM��^���q�d����?�;���7��ί�9�+P(t��-@1�p�y]~���<��� ��G��0e��$$hw���`=(��� �#7'��b�]����U��Qiܮ!h0͍�m4��M���wr��#DQf�d"%@��-~0UO�J:�B11�������KU�� �?�/:��cL��d�� �_!�2ǀ�At�x�����+�5�^cBp7�Z�t�����V��G%g�{"����ņ�Uj��1N���� 5���YB�����44��fL�/T���SSIyH`(� ��A���;��3Ő���#ۢ��S4�f��!hE-�I�2�qҔ6�C+�2���,�r0�g�\���;��J�+�Kf>��q�d�Er��ϴDJ���b�����)P�O��g�>I���֓�E'=��T�SG�G�B(�j��o���y�B�Ts��/����f_�~�^���+kOY�봔�z�	oD��ZSQ��h}�	�Z�֌�#�%�������R��KK��������
������\U:��,*�O�HY����G|�d"CG�!hwaף��cj@	�F���������>���Q��z��x6�FU���ӕ"j�E����_\%}6m�G�����՛t��0<���=ۋ*3BI�;����i��wP�K�x5��I��[��&���9ﶕ�d�?y�ê�<��}u *�&w[f[f��n+�`b7]pṡO��sJ�
T�jn:�����?ѦPr��=�:me0@w�r�I�Ǥ�M����dR�"�Ȓ�ځ�S����3�D�,&��s�����Gs��,�׆I�Ƒ��I#�b]ޥZ�9��:0I�zJ^��;�.����a<�~J��o���	�S�ٱ/]ة,��ɯ(DB���g&&�6�Xv!���]��7�KAQ�z_��n�0�������&�9̞j��oWo �ݚҫq�N�o�N�ɝ� �o����ɆIm����A�F��qئ�� ����#ʡj���FQ���yG���j���!�{�-3���5�H��� ��� Q�Ì�z�S�����WI./n~7y<�^�l�def�PY�t_�}���M��0�WZ���Q�8��o��C�>_��_k�}x�����A�m}����Q�aIs���B�L�q�C�j�b7ڻ�y��˼��7�[D�A���p�d�A���Cl>�iv��V�K�@S�$��,�ul�6����$�:���n�i��J�b6�+"̊;��B�ٻ��F���8W����}���������rY�Q��7�D����ݠ�.�=(6˫9	'�z���၃�x�k�����{�:�ܮj�e�e��Uѵ�Q_����Y��Q/��X��\L�ʈz�Y���4�P�S_I��pG����$'xv��t��L�����{�T�q7� �J�P�憡,JԿG��A�05Pu��y�;ȑ<�03+3x���{;e��T4a���N4� J�=gO������3������(@��:��&��ċA�����X���76�;׈,}��cw��F�g5��*]3�gE��z��F�e)�|�#\k>��Z�$���r��E��F9����*i��2(��~���|z�pͣy��vGgiMؼԚ>�h�{|�+yY�z۔�K�B7eO3�SN$>ߘ�����Mߙq�C��@��0Rt/I�K���+�RR����Y�!ܠ����D�	L�'C_U 	,$t��JX��}����>�W�.�<��5sp�
�Y��=v���k��]Pl��G�rM�^�0���ۨ����Am�J�S	x�o�_�g�v�­@'���K/��,�}�`dI��f���V�!G�/%�b���#J2��u��� �z�ʡ򌫅�c[$����ddK_���n ��/����$�����/n��!�.P/�z����y+�y	Y�I�e��[���`�� �"�	r�B�����I�'Ǆ�.�$.���3��C�xc���Դv<.�2J_!�U6� TE�Ɯr<�<u�!����,��-J�1���5-��ă,W�� �e8�j�s�-,��RǊf4�@8�'���S����@�*y��k��8K"����V�*r��l��%ibz��}�ެ�}s&!�Jn��&c>O��2M�_x�A�M'�.�z���12����
osL)�4� �q{Y��|f�omd(�x"lW0���H[��c��Άb�d�	ܫ�:���.���h*��!�x�%���b|Ϗ`Vdf�����l�fQo#jN{D�rzA4��U���J��@��~��ƃn*���h6K��q�+��$p��
'�v����(0ܕ#������kxj��9$�R�{~����3 a��,��4�tD�wv��=��}p���PcF�c����M�:���R�\��%���l�'����~�
��m+�����1d������r���l���!+�e>'�����X�g�[ɳ |y_|`�t��zW���I�ؼ1� �	�ǡ�&\�<���F&�����uOs�A$���߂`Mi���>��c'�7������V�If���Y��
�<�Q��dye<}�6�]i[���K�(��������lH,0qA�Z����#wm�׌��1�Y�����^e�_\<>�ǋx:�ř=���0��dUqP��W|\�%�s���0������8uQ:㚁�Γ�����;���{�d^#G�9�H|w��be�#4\��D�Gߔ����b�P�3^N��v��V���9ͫ���A�P
�>��aT��1���ԥb_��G�����Ӷ#�j�Z�?��� �0�=I��h+������o ʂՏs'�����m"�p�U�탬e��\94����,�����7Q��@����R��r-G��������d����'nw��y%���&*���3�i�H�L�N��eS�A��|���m�|
rKf�M��}�;�7�y����U�=wH�9
"V7E�yQH����*G/JP� �C�%�ge��f��0 ������Xx�R���bL;�r�ҍ��X�b�ҳ�� �����pt�6 �Ԭ5g�$��ڰ#0��>�?�*�.��R2e��$��iЍj��yTÙ�2q;�O~�s���i{��p {�_�n��a5�A�愾평fz���Jy�l�G�n5���$U�2f�W'�E�mQZ*��Ҁ?�9BF����0T�ߏ��c��u2L}�i�9sA��m%?��u�����C�_����	�h�LA�HfZ�H="~@`.빼Q�6N��Z]�WU�g%�	�jO�(�xIBB�`������\?�w�����q춅��d_؀n�	����H9ڵ��b;�ݜ��_(Gd�����{91����ς.])i��"�&qgW�S�AC(
��@)�f���w�y+IUۄ2��e��O8�>�2���7���������=6�?�Ca]���M�qcA�p��n���@���K�&JE*"Ĩ���M�`�� �s#��^��;ɤ�H�d@����fq&(!f����=��p,��"���zBq�k����Ç��̘ƒ>�t8���p���9���Kp��Nc�qe�[/͖�N�q�Y�?��S8��f��ȁ����y-K��@�HG:�>Z��ݵ�����:�����K�����/b����@�徬N���&HC���h�J��E��{��F{�StkQ�2�?TZ�8�}�O8�tQw*�|a+w.|�kB$�v[�eD�h�NFM��ݦ�'@�y
/֟�뉀�<s�����sm�����6�'
�[�a�|N�������U��c�vºlNY�Ʌi.&����Ŏ�1�?.���F��kX˿WY��.�����Fϵω����{!�]氪v�(��)�R�ĥ"����������{�_�iz@ֳ��N/��W��b�6��?�^��(T8��uABy�7�ш�h�_��3o��z�OK��Z���,��1���2�	4�,n~O�`TH��74`e�~��g~�v�=�r�!��煅�|��6l�9bV��*��W�-v�o�.�X�
[�e�fa��0س@���5Ъ��ΝS��̮P(��_��9�q� ��F����#"�h'�đU24��x	�E�E������t��oc�ZF��3�b�b��F`7
����#�����GN3S�B%X��&H�;��h�:[��Y��9`i!KF]=��XmE��&���x���-�A};�θ��fI��~�����U���2y�v줍����l}�8`T��pL'�|����%�;����5'��X�98����Ow�F�<+�z���ZM���&&��ys�;���]�Sl��V5����r����b�=H�*���kX��ٔ�a{��
ݔ�mW���E� ���i[���)i��{����A��p�)a�-�	[�d1)��:c���j��ˡ�$)&|� �\�Wf4@V�a�ۨ7�6���u�#���\%�J����1��	�!�s��!�Ӑ���DK��X�j�^��_1����D�nP�gi/N뙞�k�1���2��i��?4;�`%1�Z�B��֨))���!`Ɓ]Mb�c�d0@��f��l؀`�Tp2VO��I�s�dn.������<5�� ��*�*��Zt��V�-=]Gv�:ը�9$�w���!�n� �0O�\����*$T(>L�Q�%C��T��֮�%�?5"����
X@@guT�"v�ʛ%�2�����E�*�4�E�+�k�	���Ha�܌�K�j�Kr]l��1�.y�ͅ��kc�B?GG�L��7Em�������vLmWE���]Y�/�A@���lb���
���5=k��rGy��=�̶�����y�i@]�_��?�<����ߏ��j�$}�W��A����ؕmm1�f��m���y{����-$�,���o��FH��j ӝ���u"�Y���_�%�B먳N�&���@"z��a���H C�]�n�u���|��$�cv���Wl�T�39L��i#]��T��"}E|���â���NTz�x�vZ�W+��.ul��,"n1{2��<��e�4c.��=�7#��0�[�d��M�'�f�y���8ؚ<�~Cz����ەʱ8?�i����!��y�B55D�+az`�~..P-;�������2s�~*�i�:X1��5:��hb%��FD�0=t]me���ւ<N��N��Q�݊V]C� B��}9UB@�7�O fjѴ����{�j��_J�x#����S�o+tb ���@�vgy�<<�Y�f��+����B14���v���Y4��O��TP��L�҃^���y����~��Ђt�r�"_�<-`3�v��o}�d#?d&��a���!�_���٩RB>r�[u��v8���t�q���"�+|ҟ 3�æ �����~�ۅK��c��k�\Ɍ�7��I��+�Y�Bj�I~L���"d
��}Y\��CdL��}}?!NB}p}	{RJ_����h�O�mr�$'��?Y�A��G����������*�#A���1��W�E�ǆ���VT2m3 ]���UoPN+t� ����J�C��j�ĵ�[}���?XĞ�ZO���fϷ|�j�r �ϰ;�M�G�Oq��@K>8vа��ҏ�<�)F�=��!��A��D�,�6pw[y*����ΏX��k����t��,cWi��{�Bz,�����<b�:'�ϊ��@c�>�f�`�"��ϯ�M�b�!��IUx`ک-�*dW7=���v�0�d�=R�0�o!H�,�)^�x���wc�I����W��ᙆ�����^@zC����J��:'\�M[����i#�TT}g(�U9o�7E%�f^���l����)w���@`��+����jΘ��m Ga����XV2g!�<l���|D}3�5 B��$������c����3�ς$"��Y��0$��,�4��/�����Zt�D�F�IA�Eו��kS��|�4��)���СC}dyd�}OJ��߭���vN��v�47���B�HNx�k?qZd�j�w�c)���� [�	��?3��Xl��ա�V�p�5�G����������|w����!��>��ȈXC���Y���n��`��ϭ��<��{��]�2�o�B��9r���1�XاZ��F�ː��� |ū�P͇����Qԅ�U�[�&��m�СhR�S�:��xt�����Y�A&����C���Ǽ_	֯��P�1-�p"�V����iJ.��]4;v\U/Ҙ��ra���jW�11��"�`�o�?-ekn�:�"���o���D�V���L�I�A:6�;��d��R���i��ı����ޥ���o��?R�a��F����QP9�����%(����t�����1�����fC��J�hD	��HI��jH6q�[���o7d���rꕜ�S;��Lj����3���ԁj4ϪQ*�é^I�)�Ź���!�=-R�Și ����ڗ����?��{�ė�z"Kb���\>��z��9^�<^���CKn�#�A��B��o2G�K�� ����li�{7���,�R&sz<2��')a�JzY3�T��L�1T��`���ɝ�r/��l����u ��4��o̊;-J@�p��f+Bp���\���~��8{&T\E�g��e"X����9�Ҏeq(9���4an��)>m� )���+/��]߈�"����L��X�)���X�T����8H��h,D]+�ӑ
�u�]��>��y��������r��`-�D�v
O<�b2��G��
������R�8�|R�2USI*�%���pp2�ّ�p�+d��(�����/X����L*�n�s�1� 
�uKW?�뵼mf>��޽�J�������V(%VJ=�pJeN޽�f�wO�g��������f2_+��(&�<�{|ߎ^�:��υ�vz>����d3KCB��y��c�)�� 6��+MH��
D��(�؂�������THf�1ϟ�
lap�cϑ7Db�=M0)�8���D��<��:f����JP�R�cʷʯr�\��J^,?Ļ�L��F�05-FQ�5W�$h��ʭ�[��|n�1�9A��>AYo2Y���b0Y��_'��M�契p{6�~���j.�?��M5K;�6:���h�>��-š��u�~m�Qߠ�A6�_=mz#��r"�=��J�I^j���]-�f�d��;i0�dG�/a�}��&�/	���xѭ%ޱ�X��q�`3FG���-�xW�uyj����l�` �,Q�{"��
�6fU���a�B�m�ߚ�a��� %�ğ`�4��*���m~�.�}���*��W�+}fvk5�xA��dD�s���dɻ7p�;G(�a�	9�&�ͼ!Q2=��39��[\!�{*.>�=�;��� �P.X���P��B�ޥj�B��D(.f�S5��h�9mR�h�q�r�cSXD����ƷǸ�!y(�W���N�d���*�7��u�jӘۈm�T�|u�=��{�oH̤#b�1D��F�JȡC�O5.�L��;Z�z ��j/�m*�e�,������S�+lo����ƃ*Y���;5(���<>Gg�`&:M��@��Йe�x�yU�?�6���#\�P݃"Ģu����B�.�L�QK��:I-sX�����������l�ш�Q��}pA�gf;·���yr�ҫ�׼�n;�rO} ��0�椘�H���p ����AY�D����g��0QD�X:S�M���,2g����G+���������#��{)�!55�+��b����u�R��4z�ع<��N�)�@�n1&bȤ+P5��2�J��� �(�S��f�y�� {m^�<��o.��q���
����K]ʷj>�ԔZE*׍" m�+!���<O�l>�,Y�.�a]��Dw���4��WS��}�J��d��O�ݤw�����)BO=+�8��r�,>��D�W�:��)�\���9 v��u�G������
�G���Co���G��ּ�
�	�V�k��6'c�J��$�W��N��Ωp =�=�xi��� �:�E�;�vJ�VR�|�h�&T��Hy{��&�Ʉ|w`q��E�A$z�Cm�AiCh#�!�y�R������q�i�n,O��	�zG�q����)���,e�b"�/���R.��~�.�q]=���ި4{j˩_�9{�Z��V��30��z���(8�o^5�5��C������PT���u����kŤ:p���j�Y�=.A��Kl��0��{��0�s͞<Rn@�ߡ �F��,ѽ���M�$N���}�+�bW�!�S��?V���ͼ���W�Ѥ�q�׈��DJ�,9����%d��9��П��.�9b��7 �|*����7���,.��Q,Xn��H��]�B\�"U����&�v�,�zb�a��N��Ŕ�\\��Nw�n��.�[_�Ǝ��y�T�J��0Qh�Z��	^%���Qw��i|Z��X+�,�Xܧ������+���M�Q�6��� *�5䎺�*
��k��^c��YGʁ���mM�Q�7k �+�:s��<քIj�s"N5�������'����U������� ��gB85�2�O��*|�5$���_HB��DVAW�ASkVl%j���?ƠPg�T�J@ȉ���H9 K�G
٪�G�)�\����Pr�Q:��e}I5��*��%Ō��\_yvKm���7�%���N��F'���-��} 8�X�}���#��и@�f����f�ҟ0�SІ��g��=t'�ˑE�@k�����%��`C�,��7PY�_j�x�cp�� `�.=E%�d8t�`C �>����z�YH��+(��t0T�88��2�Q��{�S�XAcQ�Jׅ��1�AB�}bvl�@Lm^�=��o)
GA$�H��=m�v[���y�)���K<;�o6�>��Bwm��-��y��ñ�ӝ6�d9Z�*����-�̐6������!�1�����d�}	�	|= ��/!``�ؽj5_��V_�<:W�^:�v�-8�xTY�>����Bi�~�|O�Z۬ʄ12�Z$���f���3��X�`��D� ;���Cs@�܈x��3�>�T�vp�� <�!l��9�K-������r������tY��~����kM5W\o�^,�D
Сp4���[-�~Z0�=f�ɵ,�����hF�]jW�*��ΌM��'h�G_ߵ����'�Qo�#�4�� �Ak�|쪝� 閼w�4�k�%��U��ɣٯXHHj�:�?{���P�^� w� )ё�Ё�i/%�jLNh@1�j8_�]:�Y�w��Ͷ�Ł�Dr$^ȷ�y�e���	����3�ډ�ў ��\�'1+Ю�X-VB��Һ��$I\%�!Uzάc2V����<�����P6� +M��3�,�_��K��>G����|����2cŎ9Q@v��@z%U�&# �̚Ր��Q�Ȓ���)��ZB[��Xq&#���VY����龖�F�*��o���l͋:�ɯD�
27�S.f4���$��u��T�8��^/]5<�3�>]����T�"�1Y�01aحY�`�z�m� :�<��̠k��o�����.J?x������F|��̓�i\+�����_XlB�%/�sH=EU�o!��ƿ;N��P6�g��&�ɏ��m�5$V��\�=� q��Q|rHI��<�N80�#�b+Gh�,�jdk�VW6�3������{n�����?���Z���?E�֗�*�+�޷(����A�� "�(� �2�biH�@�G���d�!j�(�^,��j^��.�K}��d]�*�GR�+���q����B�;+�Y���:5���ʒ��v��fNd2œ�eTCG;D��zdr8Йy�g����rMvz����&L���	�*��L�Q���<��G�?!���oM��9R0%!@����.0x�3�/,���°`@񪴇*�5��R�x35�̰$�O�)�X�4�.��;Z6 �V7U��,�G��X�]~�����~́(
K� ��%��:���K�[����k�B����W�L�&2�Q��Xq�AY~rq�`�eZu�����P�>{tlBG�5���\顪��b�M�
0��,�Bdn|lS�V���^m��M�	�W�7|)EM���=�.P���.�#�0(j��'����Y�7TK����NoP`>܌	��1v��p�}r-�l�9S������<��ì�b��]G���"�|mZi����`���N(Q�P3Q
�c�m5�LU�������_�b
���&�%}�TՅ�Xi��d:K�)/+\�k�����ʷ�&D�3�3�:Ͳz�^vX����@9,�б���_r��wg�8���nt���������>��U��<�_����ܟla
O�g�-k�F*���yM��V:���&��|4e�VEbĝ�46�s�[R0㪶�9�u�����4�M"�����=r�ڮ��=Ķ.	!�8~�pM��h��j ���������o�e:�0V�k�(�V^����3G����T��� ��)A��2�)���?�7T��:[z��.��5ľ�+m�c7�=�V��q����Hʱ�<.r]�6�cƘ�''h��QO�)>8*� �j�ME��6�v|8�U�G ����t�o�|-G1��|�����8��J&��n�3�.݆�J�g��9�dv�#�n{�T���3��OT�������¢:9�Kl(��6�q��)��Ia�<}���čF]D-�����`.������$�JV;�%�񔽫�?�^4�sP�%u�`M��d���;�P��xM�yj�+�T��o�|���_���J)��_}�
g����GͱC�g�=�f�҃K��p �w�9n��&�C���]�D7�#��g���P,�!w�g3ӪiNg�H?��ĜÑ�̥���H�}���=o���~�� ��`������lw��������8��H��B�B��V*,�"�f1�쾠'A�ȍ�{D��ݷ#����i^f��XN:%.����>Xrt3=�(��CH�v �M�N�w%�{Pr�#N{{�c��������Sr��_���Yf�,� �k���@ w��8x?p���?F��7>�ć��>w�G��p��)���ks<�  �_�E^��'��8,���QR�rJ�P[ěҤ~��3��o�觪`AH�s���x:�ّPV��Q��v�ˆ����~@h'��}9{db/�`R��y��d��B�Q]sX���_"Ѓ2<3�a}~]�Fl�i��T@�j��D6�I�Vf�ɳ�D!�s]�Y-��5�;�0<Gk�;նK��g���V�#��sT�� ��	/ϸ���V���9# �����y�zC�Eu?�"�%�]�ndl�i~,)[�f^�����G$�
B���1E��,uP�ł���{���ʸ���Aa�ME	AYl�q�:����V	�	R�7 ���a@m��V��"��/�}?���:΍�`p��mL�N��$�J����������������?�/�+��cj��!��Gb<<[�Ic��@� i˴�O��+�3Ώ��N�x�ް��{0����ڌC!�q����V4�����pK>�a.���Z`5���)����w\�Q��-�V'�f=�n}l�["���eh�5�X����/����=TX��G�ȓ������k<���T���%�2����%�../�f��?�h���Fo�+=�X�䔬��	V������
�k��zr(�p1d�P�;'���	��P���|�q���+vX�:�������߃��RM��.e�t�G��=ަ7��P3F(c��~Nrh��ǸXX���H8�`^��Rn+S$ǥ� FD����i0�@a�̱�[��"K��Ngo<]��J�q���m�%���4���qg|]�X6�i�Jе��wޭ�ү��j�d� ���z� �C���]���V���}�i�#s���[�x��DJ�#x��At'�\� cr�5���[Z(
������-�S5�� J��}���+:#8)��20�
��vea�����\���Ha��jv��6 |=Ռ���~�#�����L�z�Ⱥ�i�m��?s\oy�"�3o.�Xk��*M�RO�����W}��C�>KB}M��\p`�<�Z�3'���x�dn��(���<ЪF��F[����K*���˟C���Z�1�m[�eUh=�U�sپ������#�2��~^����qe�dY;�bKH��������>��e	{�y��n���,R�o�N�����~���w ��D�`M6EW�7C=^����(B=_'J�a��SqMN�lԇ)hR���C� ����u" @ʇr�6s�F��/F��ގ�9��v�8T��Kܷb|+�ڶ�o:�8[�t��P+#�R(�۝hi��/�@���	X".@�`o�PO��=���:{Q�����d�G� V�P�oΘǲؙ�y���g+�u���@߿������u>��D>��#��^Nn'ů���b����+C�7մ6��������UxVJ��
�.�F����Q�M����'k�@ o��4�Y�'n�u��h�j���a��a�tn��]��z4~>5�-$�e#R��YY��.Á�)���� �det�BP�v]ʴ������(Ȍ�H7G���&�`��$X�}�y��������df��V�,&�Оk4�����
�߬X�%Z��ێ+�l�c	���(׆����⇈���iq��"h�c����/��!b}`%�E9Ao�� ���ŮFֽ��E����H�~X��U�}©5l�� n����t\(���5���rMD���_WB[�>�3�EX�����6H�
��'�Ks+ D�D��W�Nx���w9�԰x�&��4���Vc)���tלO�ZA���a�{��m�i(�P�X��Z#�P��oאs�S��k��y螘��9%U^��T�k�a[#��.8�j�a�������t�~�"�%���ё��T�v��u�L�=�U�,�i�7�rOHx����EG�Ö��<�h��I��0Q���zj&>�J��1/0|!�E�#�,7�=RQ�hP�\�o-���;�A�?�-�J��o�%��o��6��FclE#z:����Q�C��p���#nv��N&�J�\R���ޝ1o���?��<�B�7�QT��y][QYe�{J�~qZ�W����r��J����,���O���3�X�8\S��6��p�sR�_�z���� ��LUUiy)�y1@8,]�Jp�<x�#CJ�D>�|?[@�S�E�;�aJ�鎭:<�S�c�9k�:��[�k#ڇt7���W�~�96��z�}�9��T���*���p���m�fi�����+}��v���iW�$���� ��E�=F����Pe�Ê$�v�:��V�2a�7x��2zM��ۉ��w��+�fT��J�������k ���9k�&�����#"5�;����u��+i�^)�%r���T_{2$}�.잂m]���cqC�����'��n��~2��-�?A�l�0Rh3�}tsը�C@���s:�1�9��tnF�o�'��^�a� ���0r�sZv#=U[���g�X��ҽ�f�#��4q��q��U5�m�+���!�:��L�t|h�^y��@GH�iL_j�\��{|�6��� �F*f���[=�f��K��7e(������(e ���tf�i�F��߰K�	��$K�Ե����ǵ���#(���S�p ����%�M�T~j5R̲���%�(H��B6��eHr�"�`�N�_�
u�?kG^d�\�9I�A��,ޕU�믌�JY�I��y?��v�W��(�ۣ��Hj�]("�.O& |		O@�w�armP�w�;��}�{c�};��|� ����X���	h,��}��R�
=����܈%�r�s�B૑��A�֨{������D���!�+ǁ�#���
gΔZ�̃��Uh1OY�xA�&$q&�Y ����u��ɞ<y �gZg���'�e==|M�k�)]}&��� ێ�x��!vfA�Ya��{��x�;�6�/g�ص_��h��6�?=�20����5��h踠���شH(Z�%Ӧ�r�����%!�@�{R:P8�,}�i6/�������5���N�}������l6h��/�1yMVj�Iq�KB��H�@&o� c$��w7P�GU�Hy�"~m}��K�G!��mb��� �d�����}?gx��z[�'A�Rƌh�',��Fq_sJ?�4�5>t�W��L֣+lN�M��'��}�cV؎���R��C=d#;~"�����$��8眖��GQ��~n��PLk�.�X�3��j$jd���{X>�ʛ��]�����)� 긽+?>?tQyK����#�d���k�%��H2MJ���Mx������|��-�W��R/��2�]?p������Md���^J�$Z�p9$��2/3�*,<ݨ:>������֠�l���Û��E�O����$7L2X��ؙ�B@��٧o��C�aO�����}Ϟm"�2)6M7�
3%�#�7S�/h4��=ݼП<S�m���� ��97��
6j9(�xC˫[��ɘIU�*����p�"�<���܀,�}L�f� �*�$j��@�F]��+�b^:u+w���IL��8^�������ɧ^i�,W��s���c�%���Խ�:�������B>��?���G(� ���K~��u�#dZ�.;uM7�*��ƺ�qԥ$Ah��տP�L��Pqh������k��ܰi+��2�[�%G�3RM{F7�{L.��9=h��G�e���r>n���x�����9��ؚ�p�2��7��F�G�d� ��G�X�ih�`�͋;R!��`4�=ZuZ�֪���҈ ���\�Ji���D������W�U �'�QT�Y����YZ����R|ْ��l"
�=Y!!w�Kj�}B�8��&��5P}�ڭ� w�O�*��G��C8��s&.��k��S6��h���lOB�����R�7!1桿$!���c;��1�f^�P��sӹ}v�)k�Mc!!�am�F����#�u{.~�<�S��=�y$�}�iJ7���D@*��X\��1���^�y��qJl'P��ۛ~Zĳ�}���`�sЗr��kc� W'z�.4�5�{hs�j�_u�8n�e�	����9���9~�l\�;�v��+���Pv�A��i�]xH�u6�tM�\$d뮞��]��ښ��:ު��� Hb��Cg8�3o��ؼ��Li�;�63�����A�L}�A�Ä�1o��ܵQ��A#��9q^�m4Z�C��l����1-���$�[IUo�͹oS��s�����h���ER|I��K���֐`*Ku�E)b1:�8�QCƓ%�!�e���5�9=��ui	�J�����<�����q�ilTO���D�Zӕ�F�(� ��Nx�V�;�<�q�	���H�
���X� ,�U=U�u����z~�X���^�n�N	��̊w�=x�^[D:b�'oGt�;2�.L�x0�!Ԍݐu�J�zsgIp��`"=���cT;;~�Ƌ�m_��I��ʮ���􀙽5YJo 7fx2������P�slT�Y[��.Aq�@�0��H���*��c�a_aQ]<�¤>c���86tN8=�����4$t�}	z�vM���G�QF��]�\*~N����]���"��~�@8�߇���W���*B���p��-�;Jy�)��o��ڋ��L'ß=�R�p�k]gu�DX�MΥH��ڡvTGO@�i"��pvcYWCR	��Y�|��p"�֗A��E�3��5;9o���y*����w�_{�{x�Z�z�-PB��g�0N#��~7�k�"�ƛ�i��[BM�ѩ��	�&Ӻr�n�����d�K8��Rn�g6	.��Kգ����psZ�Q"(tKQn���M2{Z!�K�G�[�xڱW�9��7�9��:VB-�������=ś������6�W�D��A�.ϒhu��~[^|����� N&��vn�
�e���V�
M<�v�_�`��SBi�x#u衩T2�9����m>�&�
@f&�[�,*I�*���v�w,&17Y�u�k��-�?�ij�E���f���BF�����xѲ�a��=�hV�DՊ���c�'�i5�A���� �j٢+݌��Y���$f9g�M �39��@o�tL1󂁮$R�C���Y6��]���F4��ѩ׊����
�:��uU�A�n���'��ʝ��o������թs�t6 *�C�n��_-v)�g��?s�n&��<����ߙ�$*�����'N�YmϦ��I��/�ƱB�PBd�m���}�it��Y�`|���r?�1R R���Mo�_F �E��P�W*���D�����n>ut;���ΔA���Y �R<ՠ�����Gb
1�כ8[R�Siޔ�:n����W����Dg),"�}�F|�(�#�;G��O��)$C�r�	�MB�6_5L����F�R�ǡ��_�lN(�O��WvohE9-���֫6r���ց��$jz���$�<J����i^ǈ�$;Jю�	DC|��/�Ț9�+��@Iua)>���g�1��*d��x҈��|1�� ��W˓p�"I<nu1^52�H�FYBV[��F����A��'�9�9�Z�q��`2z��=�X��[��r�o�M?�C�'���+��c�\�$�p�R�us�9V��b��2��A��O��#��Λ��|��'Y�H ��ajU���#%���GD^gr�0.��X��O�s����9?�r;��]�H���y�v�5;�0���� >�+�M��������Y�� >�����Z�WW'�,�H��j1���]I~KD�"vC��W���/�������:q8W"Bn�Ju�e�������p���J�7�$ޙjm���#Xp��Js�,�s�TV�	��M��ϬpI��Q��j�Le,�1:5*Y�N��5�?������ڼ�P��V��?ηXs���+��)!�d��it�����{�Ȓ�LN'�n�Ym��?�C�8�/�b�7A���R7m��B�$ɍ��K�-�p����ؘ�c�<�#��`�T��,���:J��`�{�����ry���6��S�3��dP�~;���x,`"�}���gX'�E4��l���=����ȿXH}u7����q�)�������K����
l%��#���[�5Y{�D��u�fc�	���j��?�	�GS��%�ݬ��JIp��Q�p u�O�:�j�(��R�e�P�i>�\@(ɮ���ݡk��#�+1e�rF:�4� ?�N�b��|��#���d%��q5�\��q0/_�Kj�als�>A���P�C4Z�u(&A��V��H�F��:p��9�$����ұ�����BEu;qV��a%�&dxX�!��6��Q�.$�s�{�a&/*�7�+�J��?��Oru_�%��+�:7�� V�t��'� 4���6U�Vz����ԓ�x8	fVhy� �/��j�M1UQ����R�|eώ?�vi�I�Le���D~���F�gh��j���:���a2��1󨋄D� �K*C=�SWC��ŝGdE������l�@�������>�i�<O.ԕйb0�wVa��.�io�C7K�������6m:����R���.�ƣKF2)��?�C�ϛ�ʼ$��yeߌ�%�L��Qe�Uԭ�^sRO�S��c.�_?�R���2�kX�,���J��f�Zc�n��榛u)��{�+�M�qp��H���
~D�ꥉ`���7����J`?���rp���g��dg��dlUt`a�%�|M~�'�j�^�~��"T�j �U�����qʠ�ڛ�m��-�U`�56�H�����~a������;����P�H�H����/"��(^~ 8��<^y��ݼx٧����k4�X��h��4��&;�,ID ��;VH�p�nf#:�4�X���Je�ް[�.�[�R�@7�c���M�_���ld����8�>�9k���P"M=���eǇL=a͑�1d/�R?�}8k���T(1ݻ��KXJhg��j�ۊ]�-����'K�b:�q����5߀���#��a�H������β�N�\0Ds��lB⿙I+��:��d0�~��D����SM�z�C�EJ�Y�)���	���}�awz��ᠰ�_�c.t����m��w��bl?���Q�5�ݓw��>Q<{?�S��M���hPyM�2�Y�K&;��t\�D(�-D�;L��¹u��]E�ӛ8�^�����#�i�Q���oX�NY)Cj���D��OO��Dz���ǆ�f�D&����I�ȭ��$5�Hf/�Z��Og	0L�.��̲���w��$��s�s�l$���sdm,�<�t���<�{�~���~F���3+zRþGʣgsf�~��B��[�2Qo�	�	�=o_Ec-W&:kD���q&+p9�_|�B�!�m�`����J���ے����|��������yX��F��@%�!�99ch�.�!��&�=o���&p>�$Ga<O�a$��*G ߖ7��f����J��!�x�0{��ȫ��|�K��c��X"�T�o+�/��j��>�2��͢9X�*W�����gzC�y}�BQ��c���
q�(u M�l�B�\��Y��G�VM��^���9�n�8�l�9�pQ���O��f��e���J0���
��!Fd�%h#��i���%�W�ILB������)���J���>_��܎�v��� �"ZM��=��!y�fT:_'v�+D���j�����x��f���+��3)
�W^\�5�,7�j�f��{6���e?�D��]V_��Y����T1��A�H-���Lz��@`-lvb�@£J�6iI�Z�+Y�/� ���ι�����#�6�ϖ��#�t$�W��>*?뵙�Њb up�@�a�2��>�ɣ��Q��T:�cPQG�)�(��5|M�/r�d�c�+����8s's2]���b�k�@����+�3c�d,��:�'��z��8���̟/��Quգj���N�W���	���y�ⱈH��Zl����u�ؚ��>]���|�R�m��L �X|d���6	Q��;��P�\A s�ZD �'�M �)w�^�z�)�-R!���d?�)��B(�DNy���R%�ib����u����q�v	��wQC!��f�����B~��Wح��DNA��m.��X�͘�Z�rEu�	���iɄ�dP�_8�TF7\F�o~A)��>�:ϓnb� �yG����bY"�����7&�]���=m8,��}�s��J4rA�9e8����v}Pނ(��0���4k���b��D_VR���"��_��&ǒ�nOc�t����p�k�?��(�BcbϬ���e�Ϗ��@����>��
�O��*�l���B����#�ND��Z8����� �S2/U��)����iQ�Js���Ł C��%@��_� ��(��<-b6��*Y���3��
�>c�`@������.�h�:��>�q"�RL��9:G	�������@����ET.�a�Ġ�K$� �뻹��W����VN$8���o���_1�0ݠ+��#r�7��QM�H��������-p�)t��^6�SİX6�h���hZՈ/l�k`r���[ 4�PFF�Wm��_^���p��(�?�u!���/�.Z��͒���-F��kXb_�Y�7ƚm���3|LQ�e�O���_��7��1�N ��Y u�vi���/7 �P@�^�܅�Ę�"О/:�n���`)��������i�r�M/��2���SE�8�8{�i�2��� ����Y?�_U��W�>w�Gu�σM^o�3�n�X�$�7#��]	�ך��fe#pa ���
���H���S��qb4���T�y�N��Nϻr���C�^��x�v������CPI�^~Ǥͨ�8�5	���]�v� �$��u�%����w��d.X��`�I��M���]����>��4Ϣ;�U��o�\�LvW��0ޛ��^����oCzm����
}�D8�c\�
��*�0{�VU�K+�Z�fݦ�ݐ�
]D6������Kn-a�Đ�T0 =�l�:qo[z����w�͙�Z�Ud����Ę��R��2|��Ix�v��v���v,Z��e�t�.{0�&�@шZ}x^[\K�P�����T��6�B\� R<� A|��˾0���](�]�q?ߤq.,����Z���\z�F/���1~kҒ��ԮIs������$G�vVĸ�HcBg�G�9��^�i����'m=���
�e!5*Q�tF㔀�=����]������fU=��0��S��5����[�3z�s�.H��:=���H�Jp���R�&�
y��&�D(B�޻Śt�q�Є�I�"Ē���ff�^���HA>Z��ΆO��p�X���Pߞ�r�@��(#��*�د*�˲�J bN��B5�W_V!�.Uć� R�Yѭ����]>��1��wi�k��̣c�cÑ��_ί/
Z��6o��d�����0�'�6�mH���Q��Y�g���!�<;Խ%l9��,��\(4�/&SA�D2x(Jf�@��;��<��\�)W�p�֛lc0MJ=����N5�V"���=�������!�*X�Y2W"7�5r��w�C�m�7mo�2�^��p��N �	�0]�1vJ��?7a��Н�P�,s!P���@F�W�qL��N݀��L^tC�E�)��T;�|!3�*9����m��I~�s�'xgP7]�A��1�W}��+X�^�``��^����x�vh�P�/@��1e5rݢ=vT=��E���=dX���w٨���β@.�g��M0�G7�;t���Z������@��T�*����Oۛ���,�@>1�� Ah�Mx�n�=9
(8�GCv�X���}&�=��,�����3l��m��U��Z����CQ�l��5Bn���;�k��*LL�>?���R*�A��3��L�a��A �2�5�@���;����q���7&PE^g�V�_��$��/	E��DOtK�F\��C+�2��8�������VQ!W���P�4;#�������_��s�}p��	�����G2�uSd"�M�����s�D&�:3֜-WǵQ�����f��t�FD%pS:Dg��S��V�o3�l#^��&�eZB����ql�a�@�� ,�(��J��&f��V���]�z2���g�Ιck�����*��'�P�]�NK\j��9\O�����K����_��֋\��+���5���9��^C��:��������u���L�0�nd��Ў\oPi��U��e��hc�[T!:��6���:k3o��l��61/n���Ė�	ݼ��|7\4U���6�>�o���5���W��dm$5�Ay���j�.�'�=Ur�n2#Ɓ�+Ǫ�v�o���"y 6��A�jB�t�P��ˋ�)�=����C�Pl�%�$F��a�&0 �6�Cb֓ON�c�S��'3�#�E���N��Us~�$S䖀���Bh�bM����2��E�����@�H�+��L94�Tc���<���� J1�)�L�L�b\Y6�M� ���a{
�ϊ�{+w��$V���O%�k�W�U�Z��Ј�ɒ2*�=�5�g�I4�-`c�\�d���2���'��݀6��~$�%�%����8�<�z#�)x�s��o�p���#��w��W����}Z����쟣\�����>���Ka�<'��"�1(\^��|����%y�|��oe�Z'�{�]� ��Jb�N��]P)]��gN�0��xTXo�X��&�)��M���\�e�&��[�v�K�0��x�g�Hh$�z�9'�~�M���W:8�Nl�*�YhD�ze�;V^��!j��q{nl�j�d��t����`��!�{j�c��Bxy�� ���g�+C�E�Hwؽ��R	k�jA�
�.�\NÕ𹽒�*RB�g�
��G�7-�K(�� �T�]Aj���8�n�^�~�8�4���sN����iR1��� ʲl�E=_���ӋI7%� �""xzЕ>�rE{�鎌[���E�5��Đu�Ys�����eR������6SI��������(И�O�z*�����/�X��	s��%�?���H��z��E�	x<l�(�ƽi���Q���(8kr����;���g��������1���r�-׌E'�%�z���mܲz}�iGE�K�s���%Y��46�}K��Q�}j�4�ۘ�x^VV����f��&@2B������`��1�{I ��#����%#�<.�ݎ��E+�:?�����a�(f��)�5�!���+%:�f��ĬɮE����W�'����z*�6�LwkaMk��;���
��@��"D�ij�쾨�f���~���ڊO�\�$k�É���'����{V><uLum��M�rd ��h׼�3䫕��W�&pJ�qf������x��㧴'Q��\����"���S�n��Cʔ�P���p>��"H�%T5|����t��ȅew��υ�VQ��p�Q^�=� ��U�Փ)�ިA3�	��~Ϸ�K�U>�R���vQ)�& ��0�=��h�0�6M���z�cu�*�me���Y\,(����Z
M��"��x��l�����vK���ئEGw=���
��}m���g�Ջ�"��@˖䮓�S�.*�`K�,h������	��ZEoKt�2^WnٮY%�HӜ�"�dCA�&�-��>?uP�d���Qږ�n1��"�YaE�~�ci�\l��	���N��S�����7�$���d��d0�M�2�R&$3y@�F�b_��)�I�����`[˻ż�z�Y�����F��0��rYdX�v گT-.�F��LI�� #�՜9�d����\(�չ8���?�ˈ;�H4�Ox3r�� VM3�,d�=�P.��#
�$��z��;�Tt��X,�4�`��k���F�����[�@�{x�Ч+<��W��6��8�֋�F*���Of��A#"/#����'Yh�$���S?�{��g �*��T��}�%Jle��|:�#wq�E҄Q�?t=h#ݷ����8��`֙-_�v��4�D
�?�9Z�7���(�5A��1�����<�}D~h��1W�� ���ͳts�ǳ�t���V��<�'��~Z�N�ó���]���7>��aKy�('����<����|N|���
�Ə�oСh�C�&��.F1�*�_�����E�.�d�d�]u�>���c�_�j��v$���['���ե�����Ed<g�>��ѣ8��8!ԈG�벾��C]TS���Y�
NV���vJge��1(�$�m�S} �y����v�+�CNm���Y��?+'�T���I94��*�oa�h�Ym�q#�+M��\Ԍ�.6!o���M/h���q�B�ӞW͵;�^��� ��k�.�Mdz�SPp�Z8����5O�o�<̞~^� �}�x����r��L�T������T���i�<˧0c��ؠ��5p_D[�2�N�����/�u�u����p0'F�q;L��LO�����EN�����r��9&�=��%J���'Ѷ���S�͍}��-�|��NS^x����JOZht���w�SE=��cI��g�YX]~��W�?/��ƴkm�Ve�
>��\��ڜ�z��������ugl��ҥ�en{��"ܩRZ�����G���eX�8�w���D%��X�6�+^�:E�
M�I�4����(�|cCk6eiJ�s��=y~�Ou�ɗ7�ۆi2z�۔�W�̺��9K�%�*ۧ��������1��+��(i��mt�L	+����!m{A��:;6���D�99#��ӧ���@`�_'W�I��ΓS����V/��yRK���ϒ�n�Ź���f�}��j�O�a���@��^V>�_`3w�tF�M7`0rQ��~��W�,�7������_Ɯ^4�+�N��ï�Fqx�%th!�/ChO�q�.��kI���sY|S�3�����fqR�z՟3��B��_���F�1�Z����a�|�@�B]�Oߔ���Y�O8��1+)iZn@^��/�ꊑA��}���^LVe6#�������O�DY1������An��%wR�\����T&�+'|�m������t&2Sb܄�U���p`ֶăJ�(I�ѫ٩M�0��
`7~<��/67z.���M'�x��gQGp�n�$��1jiW|�*y����U��L@헖뛅�P_C�>�t�=��
Ynh"��s�ʂ�l'SU���K���L)�A}�w�u�l�\Kh�s�IK���1�D�Hq���몗Q\4�,�%,'��L̡yP+.��Q-�Q���O��8&�̘��>Wj��R���A��.ёB��0�ߴ�<���A��s�[C��R�F����z�n�	M��0u�8[��
^�hHHA������ mG���n�\vw����W*С��4��f�	gfU>�;s��P��`5�)8��)��m0ů@���&(�����$=X�ߌ��P��\��n�>��P��x ��_��B	q!���:-�?�Qc[T�w�� �Y�θgB�"ue��f����0,@�*�tu��hL��G�o*b�0�! %?����Irǯ�޽$�m�|�#�#�1�t0���ߨJ�2�p2��y�[�9�ZE��2��%بi��/��u�?'(	`Z�rǰ��j+ʟ��;>$���?��K���>�����Q�5�3}f��^NQ��F`��}��F R���A>�kܦvS�0-�ue��_Ԡ�é�)B�!�2��3����x��[xߘ���*��GA�v�1��X}�&(TR6��K�Uߔ��؞ �1����2���]Zĵ��q���f�~";����fa���� ��p-tYx_U��E@��H�l����[�@v8�*�J�S1kq�n�k�s�|az�7��nM��(v�[f�D�%q���ޠ�ZW�Z��J'kv�@�(v���g�o���I��B*H�Bl�����8����k���^R��N!���G�������<�?���~w�(L0�6gY7����=?�D��5��=�(�
�t6�l`�mOtLs�?�n������ͦ�ТL��v�eE菙�Z��e^iqD΂!y�~���t�Wz	0,�i����<f�GL��v��X ��y��%�~�E�D}�П!�XL��)U7o�=c��\�ɀ���z։0L����������Dp��SE �]�O���'J������΢���s�tبDH��������g�ڿ��V4���m%UȞO�D�I������z�V���G��y�����au6��O6�����`�3�q02��Z*���邽�ϥ��28���d����l��tU!�����%b��Ȋ>��}���s�m"5��wS��:�«�5fv��݆�s��T'��/��.�LOۜ�m��.��!`%%P�?��W���z�l�&U�C�$��J��2";��a����QƊH�tz\//"��E�-漾ڰ�jf�Z��PC$��;�$߄��D�ևN��"�붥1��!D!��I!x��� ��ܰi�O	�9��>Y肝d��%�o�v29�ۤ�w�-=n��K��c��!�0�a��ݜ�aoX�[Ш�k$�Á?��9�����ܶ麺�1�6K��������'a�,��
��1%���Z1Px;l��BGSڱs%�y[yǅ��-)��%����:uZ�,�c��ג�(��V��~ 4g�-��&6������+��9i�99<j}<���?,Rt�a���sK�|�	��{y�s�/��tI��j��	�Z~��6p��>2�XB��p��dф� �9 W&)���ʍ��Q.|��dĝ��	�D�5�z�.�,��>nu���Љ�) ����q�󟖋��}[�HO���P��%(��z��J�uխ�����F���.���������5}a���~��ڮG����wªcR�3)���oJ���E�qOZ�8#C=�s���3f�82QR�V�
MZ�)y���Sl��k~BVlp��|������-ns������x���u�ڦt(��G���������˪�M�rvq��A�%�q�>�'{�ƣ�vo��1��}L�����_j*��d�;�'�V`T�I��|C�]� �ق�ǽypLςr��j@��fEJ/�<��V&C�R�a�Q�3&��#k&�hrr�*=a]B�Y�7�F� :���C�z�j�{t�:�Mn-�
_�Gkw�3Kʞ�������D������f��=%��X&�3�W�8!2�	��(
�,C˅�YMdj��iC`��knA�.7��	 �ZسL�B#��b-�c3�[����ٙX;��+=6]c�!�js�mj{Ɖ���GT�(;6Lxs�8$v�w,누+yuC����N�i?V�z��
V~Sv���B��@=��^׍�h�� �X����~8�+|�L*��p�:���>�!�3J�L��<�p���j��C* ��[/*���@�醊�ÉQ ��6�t^�S*î�lI���C��4��`CAb�q��>�i���P�aB�n���Ei6����^Kh(��5@!�j��Ѽ W���+s�O/u2���^���$6`�Zq�t����l��P}�7A3��>�-��t����@NM4-�U�?���־~ۺD���HZ\F	�\��	��o��g�NJ������V.�w�R�
}���p�����gFι�]�񞽜�P���|������a�|(t�T��$���j���(s�VU�hL.BZ�L�����m]�.�E����*Cޔ{(�	��>�5՞�!�5����Дu���P���,���)�d��? ��lH^m&��طi������|ڲ#W����^(�U��c�;)��Y3�!�K�B�p|�_�~e\-r�'��lwM�G2^�J.!���.�%��u(=���q�ԮB��H�H��}FZ$0��'��W�!%?�G�Ą��Y6dG\5� �-x�tIٷ��>�6�X���鐽���A|�ڞ`�2Lq��3h��-��~a"�s[�}ɥ��,���(�͞D?��v������|����I`j�I�@�#�,>A �7�����!�0A]c���=v�o�C�Ӛ��&4���^r��k���J ���;�s¨�~寻� &[S��ڦ��}����nu
bK֖�$����l�`��2�,%��e�B���	$��\�b���!fV�d��sݎ�]o��`�=��������)܈ů[�G�(���d�E�F%GA�P�]6��rW�|��8�ڏ5��t|f$a�)�gշ����u.Y�7t;%S:*`�	�i�Yn�\��ԥ�p��Q��C|���ko ��GL�6�rž#� ��s"�"F�8����Ҧ.ܨ5��k��K8�2���U���88ރ[3����*��&�_5521W�i�S�����Fʓ�|�Ls̍6����t̽!ȼ�E/��8���F2��F�m:�����4�[_�;<.���;���+�J!�� ���w�L�L��y�c�n�l�8��p�ss�wh=�r��`�J�wi�ߕ���o�,��L١�*�$lN��O��n75��U��Юm�0��+�ɰ2����~n��E+�.2�)�m�R��Z��~�-��z�>���
�y��W#���!r��e�0;辖kɕ������ba*)q$��.����NV��G�����cg�w�s�7��$p(W�*4������V�_y(�|Bj���B����t�ű%?��C��#x��QIIF���Q���C|\�&���q�#�=��X++�r/����XA&.��D;�Zsj ��폺(�,yr�'F��f����䦋ÊvM�"���Y���-���w�@J���+����Q���g�>	aM>��[�%�L"�����Rӧ��&�
T��w�]������ �
�)�.WW��ޓ^~<Ę¶�D����*s#�sm��:"�xyq=R��B�,-�%y۾�B�N�
-�A:�dT�
W��K+gVX/���E�}��o|�	dɇa��J�D`:�9�ı,�ޯ$��k��D���Oe^�6Ґ�Q"Z�W�)�5�&ɲ��N9���AZ�7�wm-�G<��!�ʕG�+�%��II�B�J�K@r~�ºܗ��*�ZuRG]ə�r*�p�W/��O<\r�M��J�ü���Q�����;��|7\��.����r.�Cg�r���}+��U�"f�&S�>/I������1��/SF�����NfL�r^JSS�������������S2�[ �DzD��)�����#���;�;�����g�k�;ǉ&��a̕m��Yau���:����ۮޱx��u )T�v5���O���'�K�\�6�r���f> ��g�hA���&�5� 'd�R�"���{�7S�!!��Ӓ�P�zu��Z�t�Lm����f'��	WXm ��i;2cF�����Ib��Y8G��a��3)����^�7i�2��T� F�u��=�2�EF�&�������H��6���_G&@�4[��3���ߙ�b���v�1(P|��d������g�t�6�5�r��/���/4	�/uW�������Y���Q.�[�/��#),��,u�A��Pm���g��y�|>���E�9jMc4 ��*׽�.�8��z����E!e�VǉI��n����io��F=�J �� �`�*T��~�ݸ�Z�?f*cZ�tʈ0U��%��-f����)h�]j��8+��to-ѳ�u-��.�c������=�|����W
j�y!��݋���k͉X(�{��$�`�2F�ה�Ղ\(L��b�Y\��"��n��oj:���B����G�ҿ��$�k1L$�(���ðos���ݝ{��.����0T�"Du�	���(:�*)����%�j%���7����`���Dl^�ʌX��/��E��:y�=CX��m8ǥ���ZMC�M5���&	m����yBp���$z���)u0 ��gH�x+���חY�%vѨ��+{��ʂ$��ٙ� �,Bƀ�aɋ*��R3�ޫm���M�ܗ�j�4R�H�8.r5�]@r�=8�(�/����.�=�.h<m����Al+L����>�'��T�n��*�w�q��BF����]%��;�=r�,%P;���^7�۫j����J�s�s���
��n*�R9��!�/�¢�'�����@��5��_X�mn�\�����p�q��\��H�RZ�@3MB�7 |WUUt�\XtvM���k�b��{�q�L�V|?�A�:T���z \-/�JT0���g��^�+�Vep�=P�ڔ����>�q*Ǖ������/��L��'��p�7�Xd����B��M��`M�'0n}wi��� W�~�8jͨ�ǎ1Jʏ��V<,�c�Պe�:Vg�@!����[�,�'tz}�vy�N�sa���`oK�U\p�3y��ߣ�`%τ~I�D;@�D�|��	�@��������N%ϻ��D���=e��;ܖ1Y:ζqφ�p��0�����~����4@u�NsB��E/�<��L#��>��8C��B-�&p����4����� F����uS*��'\>�Z�1��X<H�-$��¾5�L��r�� �d��6�>Aʲ��k<4�tNOu	/�VK��k��:)��Q|��N0{���|�rvEd3� [��e���2X6X |���.��h�D&����"^�ޝ��f���K�a��x%>a�$p�uL����U�*�A��w��U���[W(4rۓ�juc�p3\\>@M{Y�E���p ����J���֤�◜��$��Ġ;H�j2��}�-������}��4 �M;�7��U�<���c�mmqF��k���"i,7� ���$�b-w�U�e�OR�`�C�.��B��zf�r���Rt�W&[V�d@�g.h�	�#����>nHތ��k�`SL��B��E9�Wf��>�Tes��=b=�װ�,�����e{��"渟�I�e��	����P�)�E�s��}�As��n5i%��v%��i���{�>�i)4K};���G���(��i0��^�u>�����3�T���-�ڝ܆'��pٷ��ȆH.�i֋��G�D��$��6i۷���H3�L%%�۟�.��#r2�M	������-�ߵCZ�Ȑ���pi<�L�ij\[��ҥi���Sg#OX#�~2�g��=�&��QŒV���4����O��p�aa�Nm�S0ݔ��H:���ek}�m Z �9i��3f��X�^.(m�%}��\kl����`e�B�a+Ͷ]裆��N86��� xr�,�P<gY���7�Y:؞y�N�Mqr�}���O�!�IdrUj�a#�!�'��E�G�J�m q��"�|hu�YJ���U�$_�<D�mxݭ��}o�/��q?4���1A�a� p��ةӑcP�>��6ӷ��U�M?�:�vXLw�Ar]'��>Q������� v�2�s~��Rަ랛��k���%�/.�/�)]�Oz��v���e�I�B�~�9�;i���F��_s���Ϻ�s}K#��.c֋h�`��ke�T�>��27�g�(�eO��)�g���+�����@:�w��@� �RV֑��o-Z�7����5|�r���P�����7�n,.�3�%c���o�ՇbC
E̤ݴη�Ó8a S�YXr�f�_�I�H���pE������p`�ux��_������V��7�dQcT^9��a2�+a,H���8e0Vr��w�et�c�K�+�h��Bi�?�T֋���I����3�q��;C���Ɇ��8�]����XD�N�#��ϹE���$�	�;z��Vk�ǳ#�]�!S�?��R�^S�5���R,�0j8e�1���b�۠�Qi�T�LA��k�H�n�!�L�B�<��N���2gt�	���z�٣P� R�J�`�U��K��)º�+lV�54æAu�hG;Ϊ��/a5zk;X�d����]�M�u��d�k��ut�sk�K_��y
ͳ$;��,�o;c�%���;��b\�̍�M͍:��_�/"؈��ȵ礇�����eʚ��	���-��>yW��uƳ��R������%ddY
�J�*E��%����"���v�j�G��)y �P�ji�ŝdS�� �Q�0����*���k�h�A�,���,U�^u�^�&����m��#���.�h��*c�J��v-��(?ϛ���k�l��V��A$7ôsZ��2���9r(�}U���Kw^2;����񧓒xP���]z1��VL�ο��چ'����/3��x�����̬�-�a�*��1"[z�͌U녡�R�,�$��"D�{�bX�pQ��T�v�J�������J���pL\�H�n�s���3_}��O�o�����Ag�F"���;v�pc��l��Xn]�c�J6�� ���g���^��yL�3lv�[�/r�i�}" �9��S¤K��B���h��b�f*�MOV����y\X��_wѝ
 �b�jf���3�X-�b��0��
��f�|xs�+:g�FH�O2�������>F
���t�'C��l�j��i�Qc}��$.y\űt�����0�'IG'J'w��ɶ���.�9Y�1����ϕ�I��üx�J|���:�ԅ�Id	쉝��EJ}�l��?N��e�8!�����r��Ԛ�!C�ۭ���n�.L�x�p��w�sA{����׊�i�0�Ol�����d�{���		�
�_��#�Eɘ>���k��p� ��Еv��l��iHb��U���w������e�!i4ߡ�~�~ʅ�hq��a�эw�`�^�YB�HZ8||�](�;.␖$�(�Ĝ/�J�̪��ʐ}����s��|u�n��?,em6�/�Q��z���G�IX��z�$-@��?�[*[ݹq��G�t5�i^��<�B�|�~e0\P�漘�5����1��i^�}=����h�{L)����P�xr����w�D������B�q�y�
/gAϮ���$rʕ�m��4�3>î?�~]��")˺��osnsN��Ζ:�ǔp�zD�ь��˴=[��z�L�-8�ô�������M�G�r�$@���ԗ�с�+�_	��\���]T��Y����R���S��=Ψ��s��703��ĸ9��1�+����nKI��`.����%iђQHB/�,|ߒ�>���i���E���s��	�Fo��SJ��j���1�R]��#.���/������	׉ю�bp��U2Hr� �[I���߭�D���F3n6�O��(���cU����R3O8��i�0�RJS�����?A��G
�RcO�)��oYʸ̞b���㩌)�a�X��񮖩��C����|Eo*��x�1E�8�z7
Ǡ���l��U�rV�� ۹1�	ބx�%i���_�W�C�7��b��m��"B�F���;�7�5��CVVD�-:TB
=�	�ߕ�9B�(�e@w������p��X�^;��aD�a��'o.s����R����P��!�޻�jh�ό:=���,rw�V�cm�g<iǶr!��J�2#�FS�4oHA�./o�n�3@�Dp-�S|ƭU�Q�+�x)o$��Y�;1*�Q�C������3����5U�Z�`�E�)�v�q�%���Sg�gf!@F�lg���n_C	।�H�x�[�[@�/nA���9m�N78��+Bj=�����i&}��8��56\��G�N4H���BSH$x���;~��Z}��Ԉ�ܶ/l^gͅ�b�lf"C��/5�i%$I"�~k����m^�n��L��q�EO]I�R�k �5���VK�%*��u����r������$�ʰ�+�`�}�H���D`l�z)�ҷ�2;HMz���+7�JK����BUU+�hh? �f���1��g_�U%s�T�2��69j��Ε�[��{s�hcC mF^��F��/���hS�����^�.��'�Bi�0�Y# ��
��w���9�p��G~?؏_�S67�crDԑr��nQ�@�P�?��)%}]�G6=��,
���9Tjl��5Ī�����(��[��_=����7�[?��Z!^�N�/g�28�L�0s6־{���A����6����C��Q ���k���ݜ )�j���fP�`��b�����RM@r���2��P�"}K_��Q�_�N�^���[��7�P��/�شZ�sg��	cGN9q�	�7�@�^�R��B�"�N���kqFbi�A�P$�Hl���ΛNN�G���`�HO�X՘[��ݟZ*h��	�� �с���.�eN_��U"����sӷ�����L�Ȏ�*�}��Bw�1e�X���y�ĸu�v��<ɗ=�mMV���g���P`s{G�����Cdh?3Ѯ����	^�1q"�����͆s+�������*�^�� ���Z/����k�Y�J����Ȁ�h�pX���K��8���ޡR���	s�\�m<-�ކf��K� ,���95�8�p�����W�1L�dy�f>Q<��b,`�|s#�������1�O+m`�O/�1������$�z���Է�1���A�^��B�6h�$�!#�m�tU������3��U�KAP�o��NU�.f`����H�'��D#7Q���BJʁ�z��P���������ŷ�- f��UhM�.��<X�u��X[��X,?�������p���}z[�0��:+�`Q�o��+~0�>�G �..�qJ=�`}*�����@7i�r ������3��� D3C���EX��l���������>x�x{0���#:[�����SCڇ2x�7_��L��U�4��8�3u��a
(���?�0d<�ՆQ?�O�q{�=��W��hR�4�귏�r��t.q��COT<�Ϥ�>�6w(��gʲh���lF.Uv֣h��־��f,'���+|i���G���7%�:�Ġ��!�>ak�q�5�|���D�	:���z�`� L{%��sTw�ə�H�u��-w��&�����û(\�:M����L^#U:w�fz��%����Т ��}�Y����%��q����ǯN�U\Y{��J�Cj_���(A���s�#�Գ]�YQZ�ҩ!�n�g,�pEy�Ħ1w�錁������ �v��e~T�������_�
��O������佶u���nJ�M���'��&(���N3��'�V�:�뵖�	���YLU"�q�d�̶�ZyqyIL�H�y#�U�{��e,/!���GX�nU�"�
7uZ�Hc�,ig"'��=�D��1�&0Q������9"��t�)6a��B�k�C
13#���&HR"��{��PB��w�����<N�I�ak��ـ:{��;�\�v��*1�m>�s�kx���[�E�SDq����(Z�:�^���"3�~���=��;m���\4���}s��DL"m�_��$�"��C-y���㾂WKNcYŽ���萢�e��N;���Zx/�H�&@����-�CJI��s�X�9�q�p�i*;y�$�E�҃Oڮ�V�����ɖz;�Nz�ա�==�%���麳>˩���)t�� �"�|7�ӱ��-�.�4I��o�]MĤ)���zy����4ņ�lsɡ���X�ޚ��+�=�V����밯�C9� ������1�^m��A���~��**�_�Ü�X|i37dO6�C���':q.��+�!!�Z>�G���M����X��!xM�׃s:K�B;��|Х��HmdL�ݚ�WS��Q�.Un�6�̃I^�e� @����9����Z\oY�ޡ����#0	��4��^ɚ�Z7Ա|�����b�N3_7�������YQ�B��-�������m?�9bۚ�!���,�nެN�X8�P45ܼb���9����3�R��w���2�T9�X������,h	�.lE����� �c�4��WN����}K̢�͌��v�@{��V����Of�Pn5#菠�7�G��@+�LM������p�`S���Fi��}�J��#-��y�U�K�L
+:�ښ J  ��1����>��b�/YM��H]^�۷	c����x���Y�GF>fՈ�c�m��uA���
��ƎOݣ�X�=�L�ik4���R��[���cZ����&@���:D�K1\�T?wb4��O:��U7�K/7�����=�(X
�s�A�]�5!pnEi�Ԟ�����͠�v�2�����n"��8�a#���,�����X�=�2_4�ׁW�ò	#7k���U
EIk��2.���O`i���� dd�>ެ�		��)�ع����4���Z�,�H`qF�'ಓV��)�����\��p���7F�֕}�z5� ����W���#��Io���Mxܖf{J&���>�����c�t%B6���7�|�����1I�d���iA�h ej�q��Z�'(�W5���-��%!m��RR�d���V�̿z�����r�0%/N2�-)cGf|��^���՗��%�Ꝺ������o3�Y��� ���G��E���Z��X�-���;*�2��`3�E��$4<�I0H�����6�=I��V#wG"�<�K�&#n�ĕf9U�����LP�K��"d��v��@]c��uLu�>����4��Y}5���x�H�DU����
�c�D��'Ala�Mޅ ��>�*s���
s~�`�s�n^<����B���:;s�]}� ߦm޴�[��ׁ��§C� �n9o��KAh���N�(L9�0^شp,%V'�ǹ���Գ7��F�!Y��e��KN�}�MEX�j��]0�{���1e�UT���S4�P�{N?�T�&C!-�Hݒ@Х�9�1��#lR��|�LKp%����e�`U�vFZ��u��*yY�0�e"����\����Ϭ h��o���SVS͝�?��Y�!W�#	�i�}���	�p0l[�xV��˵��5��@2�B$E�l#��O�͊o�?B�ty���sC|���>n&G�[�j��lJ�nm�T�3�
:V�-j?�� �	�IՐhu����J<,�l;�S�	�.�	�dF���A�#��K�-ӷ��?I������?l.5g�����F��*���S:3�joo�h=���ތ����ӆ!�v3�C�֪���^n���N�@�0�VO�P5�L�\t:��vu���j�[˴�̌;*��Ox��t��y��)�ET�Ù7����²�;N���׀0��Yv?�3����[�LTy$�������찫���F[��q�qw�s�I�1E���c�ﰋ=YE�!Z�6��w�Wq��R+ �a�dlv/��U�! �H�Ҷ$Tօ]���`�ڃuS��T�Ģbl�� k	�L �W�\�xզG�1��KJ�����}R��*�	>�D2��u����t���mLqn�.��`Vdc)�@$"��v�{c���j�����F3�vl�	_۸+�Y�s ��V�X�"jjt����PFb70ֽ�{�O-�H�sv="\�q���y���e�z^�!�����8h+6(��1P����-X׍������tef-�W�LW��1�y�I�\O!q��ȹ�X]��}�\�����k�:��L:_�������.9AJǱ�0�W�1�	��E� #�6ڋ�ݗ",�83�$D	��皮XP�A���'Y��z�x*_}z�w���/���A��@����s9-������lt�S��&�p�Ih�9����2�Ԉ���3/]��/�����W �I����UF(s�ߝH���ⴛ�~�dEt�>�h�{�7z�8v.쭔����)CF�M�8�9��d����ґ���R2��5��Q���VZ�[��ȨC���Är�w�`�[ �o��~�g1���U_ J�P�ʑP�0�����f(�Uߣ��j &76 �֗�$����;��Ǣ�Y�kLfu�b�yw��[±�uG�f�w����J�o2�l�ݮ���
N�_w�|,ݵWb1�{�Pl?@)�y�v��u�"o��3���*���y�8�E��t�M�h�E>�e�ʩ��9be\l�e�O$��,�Έ�i>?�+7��v�F�Hh�N���>F����C��Fp0y9��S�SÉg�o|�M�2��[�U%�G;u%�<�3
�rAҁ�A���T#g�p\lݯS�YC�b���v[xYۿ�"A^B&��aR\	�J�O�3>��|(�7x!�?�mv�܎�.�f'�X��i[��z�:��7�#
vK|��Ko�3G[��
����%�[ȹ��(�H�R��bH�d��tiu{>1��~�{��ľ�O�M��|��p��\r��J(ݛU���k��~��q���|�2�am)6�z7�5����3"�] ���?wj����?�<
b��1xQ��M�XK���~*���+���(ص����j��D�Z���_9!�K�DX��!����w���H)��/�wa��1`([C�t���^m�㤪�;�����x.!5��2�i��p��N�kE���竤E�p��j��5���~������OH���P&��d���S���L��fWR��� �����Ġa�+�eo���s�����=�l��#�S�jÕ�W0p�߼PI\�����:�V�O���?�GZس٨�Q���m����N��׆�0�������10�Kq=�~�}I�6@~Q
�U�py�(�n.��70�ɿϴN��΂������Z8ys�/F��)��yk�d���`�眶�@H�+^��@
����y��k���r{��|�$�'�kr�C�tr�\��%5�y�b�8��C+Zī�]E��i��V��>B얣)DB+Kc�����Y��r���'��[H�b��AJB'�FM����!� ��h0�x�y��C�^�z�J�mu�FB?��(�zp/kh&6����!�;��{o�Y�xHj����Y�r�{{7��,Z>�ȡ+�m�r�'�d�6~����,��|���37��|��O3m9����*���kT�	��>�*#�SN�?��Z��ZO�ږ=�$.�c��#wA볚k%O�g���ۢKÖ���b+�뽠�#0��Ś3�}`uB�5�����@ ǧ�$�͈��ŕ{M5����~���J�q��t�,���r�ڀ��vو��ւ����qwd��&uN��g8��hJ�?��um}�󰨨�Fջ�3fK�	}�QgJ.�,D\h���iC(Q�$K�A�w��w��nz���c��? �E�:�!� `�тSɓ�m���I<rY���� ��b���(��K���W5��J"������yL�O�M�9���`����*N���Cu�۝�Q?���/T����<��)���M�2p�^��ZCXP�j��T��2D��/'ӓs]�d'�z��{��^�	2⣇*����ƣfȟ�QLd�R~��v�s�D���@�=\\�T�ê����`�L��I#�;:�Q�,?b��?��/:� ��-F�2�k/x�g���H�b}=_]gja+(�����Sr��_ȿ`V�b��ִ*}�!�j�]s>W���')>�X&}�@����,9!�Wi3��^U��9y�7Pm��2��Y�}�t��;U@1�4�o.��t�;e�\�M���2��iSed%!���FmULc�u���~,�vY9�|�}'}ʯ<D�%DoJ@�3���uaw̏�V��,�����\�|9堼�+0������m�"�sj.�?����X�4x�^|g�1S��Hz�G�S�(3p.K��X�܈{����x>v������S+����=���Da#�_k�!��;��{<�3]��� ���P���ݙL�M}3m��2�����(��!4��6��q�/Y ѳ�y���as���s/�'8P���L�s ��0�� �v�����JI���+8l�gP(��2������P�����ܹfK���k]�~�l!��q=q����J<����dW�z
2M������3��i` �7�9g\N����t�8�P��6'������2i�i&�zat�u�Vͯ���B�ds�W�B�2��$��'������O�wm�D�Ev�f�F�8���o�,��/�_�v[[��9l?�d3+�׆]L-l����|;h�?����`)��n��ì��~Hh#���M����4���Z����%un�_9����UK���l�*i�����_q��',,]-�LH7!>W�T�ixh;�溬-�����������`E���]b4vR��K���3w�DCT���l���%�=N�x�Fq ��h�в���<?|�������MSGb]X"�hD�xlJ�!��{z��|%���VNƸhﹽ(Ȯ`H��mb�+
��~��MM����\%Ǭ���&��ۉj�Ւl��2�q�sSְG�������Z�5�v ������Pz�6���'�<�AVș����>{TLҧ��tw2��ٹ�&ٕ}�Ѩ�q�Dg�!1�Ŗ�Ƨ;��ja���0��U��'3�]]�E�/I6!����Ď��]n�7�>�J�:��9tI׌�mW��f}�̏kd�/ ;����M��ġ8I�0�R߃�2�ǲ��s�I��3�}~�P��w�އo �^=\Y(E=:���s�����m��^�`*c��)�7������E(�9[}H��9�K]���8Blh'��y �	a��t����hBq����ГC���tK#�fO*���9d�W�>3�邆�9B�nߦU:'lW�_��I�������L4<}��6���Q���{��א�#���n:u��/|�u5%[�V�T������Հ���*�@�(͢D�2g���^4߰YY������O�`Bru}~G�_I9�m�@ű=[�G�.k"IID��#��w`�ճ�&p�=�Gx,C��ݚ����l/������iMb�'Y�]��>����ط�9a�/!0��/8.��1c�b4f���~%���p߇b
	ʍ!PY���X�Iuj�ùf�+�Opsk���q��%�r�`��i��an�`ȸ��j �5�.j�^��v1pul��k���3���6?@T���-b]ܓ�ђ���Ϩt�ṹ�IN.��y�CG�r���)y�i����mK�-�O`�#Pߎf��<i�O�;K�X��T.�|���]�L%� �s�_ZK�O���G��Β3|is�tS����U�� �+Y;�l� uQ9.y]be��j뻬�r��ِ��#�V��7�s��W,�J�O5�9)�i�(�,Q8s��A!� ],�j6�rU��FS%)��mS~]��]P��eS\Z�!C��:��8�l���Z�Tj�zT&n���e�ma
����j�.�_@[KN�Y-q�:�b��Sc�CF����%���tE�<]N�J��=Ƙ�����E"��R�������E�ݦZ����ki5�	�|�@2!�����ɄG�{ҟ��1	f����D�{��
�[v�q��:8Xq�8�1j�dL*������PY�Tn"�OuE��sa热*�Kq>��T-1'��ʧ��5������~�����q�p3�?�����l�@�tjo�g[��� %݋���p�GdAP���G��"Cv�����K�~3)�I�8~6�ϊ8%�TV:V/#�*>0uW�&E����粭����c���䴄�I��p��L�bq �'��(2
�-)���׾p��B_��\{�R�\&u�o9��ˁb�(���1�	H]�y�#%��6FN{.�j�(iR���0����.l�~@e�"Lz;���Ʀ5n-7�wLw�
��������R�58"���)�V�� �g���Lہ��͖�=������}�o�J傆�?�'^�^�,��59\��U���/�3pgJm��E�Ȏs��)��O)оy�����QX�3lpŕ<`bEs`���[�����7�_Ꙩ��|r\3�'D>`��&�V��h&
�$�c��!�Ԯ��zB����K�*�4������C�!�9}��>�jD0�ȑ%0��u�?�Os���8M=�+&��r9��� (P"u�`�z�
H�T�՗6��Q˪i!��ig��V�Q�z�GÏg�K7Y��e����g�HD�2I����P\�V������g��O��M��/q:���
�(�xg��E+V!�߅�q�����J��@ʱ�Ф5紃�X {���������u����Guk�9���0�m1샡�_�������5 ����r9�?�1����z�1�
-�-�1Ȋ3�����i�uk&=���
k>υ�Tȏi`*,���[��]Â�C�K�ڮ,<8Ѱj��M���`-�>�c�z ��&�:~M���PU'\S�O���n�5�8^���wT�'�%�,ұ�'Z�8�:z�)0d�S�i_f��'�p�d��Hήb%���م0'?I�>��{��L�J͗���#Ѐ�������o�K�}�%띯B�Ub�8�?,������U�	ʽ.U�)�קDb���G1�\�uM�����ȯ2��z�';Q'�p�[��uOW�G�p�8dn��+�2�9Ĳ��~�R������;	����kÊ�9�1���%@7��Ӌ�h(�)<��������K]�\N��^��%����Q�]x��Y'Ό�H�<�N�b,��c:1�w�����o��[�v��j|K��ƍe���
)�i*e������h��Tpx�FC� 'S���5q���=!/!��|ua\����9P���+%��g�U�	6���O��JlS�O�����H��d	z��ʂ��5��bC)��������O���`�Q�s04[��_ҟ�g����d�2�{�lYu�q�������,|�/$���b{?4�c��곎�e|��t&�A��n ݅��T��6���P�eV"63�}���B�$��(�����֞�SE�6GU8�F=��H2�>vh�u0|��~bX	8����K�8 4IEr*����W��g�����dH�꘺G�>ۻ�_��z6%�����=m��e%⭜�����!��I�E�d�������l�Š[��D#ή���q�,�0#m��(�8H�ښ��+V�D��)#�,Ø�/�f���e�
vmķi�*�嬬���o���C��3~���W������=��)�U�&�d�h%k��ё���m5o%q�lt�M�6�R���_�ɻ��RT�ΉF�I[݌��-��b���2ԠB\�P����`46ö���b���%�k��d�s�i�A��n޺Oط�KL��ЁO�P�Wķ2ˁ<����M��?׭zTe�f�����.�ZU:@����5���������DT�
�b����}a�ȢxSF_�l��׎���־�*��z$>=E�U��
�%�z��a�k�̹�@8��zd�ܔ������q5jʟ#��&��D�/c���l�&'��D�o�A׵,�q9$�1���h�9�J��&`Esg���,�b���	)�L6�O�j�LE���n2;}���&�W ����#��,<|nyNa�vy�BO��ig���q/U�1�_�f�~AR-�,��[r�����D�$ĸrʫ�\1Od��xt�i!ݥG� �x�Z��.�ZU/�\$eu%�b��e����_�� �� ��Cw6�b/�`��iO��L�NG�[�+�S�������Ƨ��h(썎�S�fd���W���L��]X�3�-�v�����f�m���p��#:M�QZ�?�����7����.AW3D1����_^y��W��`o�f���i��Rʏ���T��W����{���(2����M_ޕ7HMY�Q7�-�+� �uz �֩��$>˜霓IAC�3fͦ��٫��J�[�Q~�F4��aR���A�v���%o����AAESr冼R�oe+�hj�d=��J�Jo�T� �x)rN H����U�F���y��㙏E���k��X�W�揿 n! P���W��2�����n����"E�ع��Y� p�Ha���Wi�0c���,���/����v�
�_^� �rqc���:ѡ=ho�>��H,l�v�g�N-�2R�����R��aW�}�j�h��D�e�n[U���nT�+�|c<6�>c�`Β��3a`�?����>.� D��P�J˛\e���9�@�ؕL_�D��ꬭY=T�=�''��,��03h �Q>̛P'�uI;��.Ǐph"i]Kh��Y+��;#L��Z國/����)^�}�{��󸔔��E`  ���Cl$֕ג�@�}����a�C�ư٪�u�8F�rm� K!e��{`K+���W��&�}�R/����@�:���ox�ڭ��S�D`fW�ԫ�֓DO��x�ҞoPi�is(���Սex�>���Q�Ⲅv^\x�7��Fj[]���Z�ʢC[�c�d�i�D>l��|6��Z�pi��}�X^I���K8���H9�w>N�|�җ#(h���6B�p#��>�%���2dxƁ��g���ԣ�3��n:��_�Y�mw\�OI��nc���Ø��F��)8�x��rm:�Lz�ȷ�HZAc�0X���CX�v��	���p��6���:/� �%6X�:Kk�tm Xe�6�?�ie��T&{��u�Ÿ+��H\�ZJ�� &kw�Tv%a=K���{3,>�=k�im��.3OV��^��.�2��+�=��Q�F��3�����	s�'i0l�B��HM2Ʒ�y�0�m ��$��Ŕj�����F���_��s:�5�z�p"�q����0O������_�E��Cì�ޫڔ�~��g���e�2��Nډ\e�%c���C �=���9F�8�&֖�B���O���rfJ�%��owƱ)HJ\B��1�C,;`�㣍��bl�E�:���0ڧH|X�{��_��zD���A+h�)����Y�F�-"�b��b�nで*�$��k/������x��x�}�5;�@�R��ZG՚�a=	����I�P[a�۹#k�~gGZ���Rc~����aN�e+�~A����|/.��$9��tV�b7h+]�9�&��sz�3bz˘;eP�;RM��߿�H���3�My�k�t~#�rM"�:Qα�9�C��XGp�Ss[�����`���S*��jq��y�dD�����BNZ:"K�Z{�}Hcg�B�AF>���s���'�O�� �	��3��|1�L�*�M�SF�+���#b�A�䧭	S�z���0��j����Ȱ:`S]�7N�5�<'0�yi����?p�s@+)��+3�?��f�u����#(R��/Ä�Z�9|��C,���E���<Ӥ��� ��72*��R�I�.�HJ1X��S}��J]��M�����AH��}����ϰ���	hR^д���a0#)-]�D`�b`�~j���M��œp<��5�I�H;���G��"�?m��he<�6��a�e���R�jF#h���5nWi��cݱyf��iX���w˨�JTȬĜ���I���b�zq��Վ�/��S&P�7I�`/I>������}`����)!�$��Y�������~���w�A"1%w��i$*�;c���*X���3��0_�Q�aw���0Vl��<�c&��m��/��lM%;H$T�mh�իc�����zpZi�5F���Rz�O֠�l-�n_�}��m��9�I�ՂP�",>�4i׫C�h��APʪ8IY|]_���T�)$����X��Z�N���� ��)�����E�d�L������>E�((Y��fS��k��1`�D0�b�:�M��HBQ�o���.׳#ә����2����5�FP[�B�S�@�d�d����SfH��ኽ	Y������Vꇭ��s�Y0�4	/�0��#֧𘐩i�SP�` 1P ��}7�C����wu�s�G��V�p�(yߙa'�Q��c����)��Y[Uf8�"��@[���D��q 6g(f�G��F<$������d�rP�&
LI�h�4����"�[�Nw_z�97���>��!X�c� �gd��H��V.ƹuٴh+�zzbFd�����s�&+��']���?���oVi�2�SIZ�^w�V2#�5�B���풘 G�aG����r���)��?k�����yϸ��I�5�_:$JL���D�gO/|�gB�8��s�y&��.�qt3�2���q��Q�Y���h�cK��ꮐK��;�WBZk����ц��%)�8�s��c�F��<h���hG�\�&A,����L�E��}�f��2^dQgt���[���+�,���4"`&y��߭p�^���=(T�� ��f�����>g;xx�X*��oA���i�ض4A� �$4�}�A�!g�Ly�ZǱ��N����]�@�8z�q\S-IM(p���P�1lͶ��q�`�@Q(�"o�S���� ��, 1�EL��FA��zD}
\�>w䮖ch�-ubCt�z�.o�H�"��LH`=�5��Y��`J��H��_��	��{0�A"O��F��S��Y
���\�Q�^>��/\>��c״Hf�D�-W$�+0�胂�u�ă�8fw�-s7�l�w�����{�=�����K���o�<l�����R��M��Q��
U��P&Sh�{��=<�
���y��Zon��N'&�&�p��s�|�q}�I��Xi}����(��6�م��D�^�[ʟ��v�����U%�A�"1:��E,�<��N�]U�u��)@m��0��	��(@��s�9;H� �uؔ�D����HP� �CD����J���k.�\Or9|i��;#y��f!�l�ڮ�0��r��vܴt����PАz9;
�ף�m �X&9���q��/�w�b��"t��iЕ�5?2��9/�f4�g/ �Z�2ו�'��ߩ�܉ؖ"u�\��aG�K���Ӗ��x���_)�E�-�x�G�������=�aE#3)��]�1���ʻ>�y�!���E��H�s�Y��k-^/\G�7�ஷ1vj��J�EG��Sn� ʾ�|�RJ}|H5�E�s�Q��^/��}V_�������%��SG�=l����5�Nur��s
�'����M�A�Y�2��A��~������hJ�V����I���]6���j!�"0n��敾kn A�N�T�Jqρ�z�ߏ=�&כ8,;y�>�t�����
�v���ď*��*���9�pe�7X��ɨ���kf�g�?a�o���&�J�T�Y�/�S}3T�6��OR����?�*�d�D&.����EO%K�Ћ�ŵ����y~K��,�������(�;�o�=�s�I5�P.c�ߖ���:��,i!�^2b�k�+�Y�� �9�ۀN��W���]����+�sD;
�ɘ�v.�uWS�W�og	�oA�~")X]jN١A���+T���c(,RR	X�·�+j,D��$ԕ�ZM�/��)n T���W3�^�j�PRiI9����8��Q��?��ɷM�G��h,���β��ZJ_��鎀f�/2T�aYHa�Ȟ�V��6<����pM�$-/�����D��'�tJ ͯeR�<'�@����=���z�y�]��	�g�3�Z���=��\AFU��ʾ�*�Ȩ�2s+n ,!�{�\@m�NϓOQ7���8���۝]W�D��c#F$��XإB��2����>lJ�`�D�L�Q�b��Q���pd����e�LRft�<jC�D$����; ���N���1�۷޷���/.�%T�G5?����︫-��ƣ��^6ԣL/��jU,��71�]YHY������*}f��.L�9o���&ߘ5���~��g�k̪���I�e�.�֘Ԑ̵�-�$�3��>]�M�/�ҩ� �rf���E@��o�V&X���~R�OCO΃�A�V���;b�ڡ�S�jA~��#�6X���y�iJ�Q�V�b��,2l���>�`"��Ri'P���h�!���L�ݖ-�L�Ї�����J`�H�	l�cQ�w�3RiőQ�b��8��=����Gv_pk�R(6ߩ�ܙMٝ#�&G肐��7�.u��i�CU3*)EU��f������Yb4�A�w���� ��hʩ��^k���e�W��m�G�'lQv��"�
��,���N�d���P`p��%|�ub̾��|�P�6x+t���T7uF�.�I?�6p�p��(����$p�t"�]��W�o���~��r����q.t���o�5�H<��  T�G+a[���1�D|�?�?�+O�m:�����W=�4P�;�p1Zk�`�A���|}�3���N�)���nf�����p�f "n+j�(����u�n�c�x�Gg�2�	�t����-3�,���{�(\�9��8]�gG{P��MCh�D0	'�ĕЇTO41B( �9��p`������ˢxqW] ���쁆=h�(��b�ڒ܂>���O�����+i�g�D�Z'	�����ߝGե��77�Y���bВI��[��,Gfe�%~��xB�x&K�h`Ww�&m%�{M��{�����?��F/�x��&G�G.1��xl�M�����,"sf%�����}��!�����{	��3�ȖC��I��)A�}Y�ɖ�����˒!�jkX��D"�y{����EX��YFr8r�Ӣ�5]�_%]^?B�������i܄A�-�I���03��ٱygZږ��$�A���'@��h\�x�$�УM�Ix�	Ԓ���۝�*aD�}�eG-���?�XI-˽��>����	�<�
"����(4��9�VڸF���ic���-��q���y���د��TQ�̖? ��  ���x{Q������]iiB��҂�[�|�!�I�n|`=��IɈ=�>��S����4Iz�8�yJB�i��e��� �r��v1>����9�{`S^T�袝�?C����I�E��ޝB���uH���(T��^y�
6XYO�J��2��*wi�z�7k�c�%g�,S��3���� ��8��/4��F[o���Y���Qop��뗝���O�f�E&�����V�08[}��63I���z�~����卫�Oû�wc>�����`�b��3��3|B���t���v^t��Z*꿃�����"$��M���	W�?�۔�*'���Qsx^�YZ�u�Z�j�I^�����P3��;/J����X�w /%��;�C�ݘ=�@j�):�
���	$&�A>&�Z����A(��e����>+�9>"��M=!�P���`<M�㰔{�E�`�}>u>{�{-��@��:��F�;^U�&�� �u<��>g�PX����rH��p��~�v&�w\��|"?d�:E��2Cy2R��a����2L���V@�Fõ/��O�����i�T'��{b� �cq�E�Z��	oh��ދ�z�<ϳ��jؠ��P������Uq�j��PaI��;�[��f{@�DDg%wC�?�߆۸#�@d���շ�Y)*�>�J��9� �j�z۾K�z���<��`'��??
��5Cª�����2��q�W�4vK�4Q�U>�/���=-@�)\�*� �$��GXU��l3�|IX�t���V+�����_۴BmA�Sj�8�/d�E:n�T
h�R؎�D/~��.ܝ���[g9��oXq�i<U?�@ܻ5 ����ߛق��&[B�uE���"�A�~g'��o�"��ъ�  R�}�� ��C���\��Ѽ*$H�h��������Y�#N*Y�N�ÔD�
�䰩5�xɣ��?�ޭP�Ś/�3q�0�c��F���i=�MpU�V;���D̞��z(]I��[U$
j%s��>
[�]AMN-�択æ���|?�i�_ڽ�k.hو���suD���*4���<�+������¥�8'������/���;���8��ۍ�=�B�u��j?8SE}�Ŕ� �Q~D`>˿�)	"�y���?iM�v���p^K6�.o�P����H_���`gЛ)[�\oo_Sz�ֻ��MK�UЭj`9�/�v��E�)՚O'#�c�t��� z�����֤$gw�X�G9w�o���]���A�)Anx��ؕ�#��&[�zD�ִ�_�����a��P׃D�hnG,䔘��R�Lf�������qu�n�ù^V�F�ʯ��2x|�i��v2\Ł��;K+�a�a�����氍*^���j�@;�_Eb6�7��-��Co)܉�6m��zRE9��������F[K_���lM|�}���"�;���#�!��RS��V�MP�/8�����TBdb�d�p�f�� �%�Z�������}��L����c۴��T��V�'�C�,<:���03|���ˉj'�>���
���C�vc\ DuA;A����¹����H�7�{�s�������<�e�A�-���Ў����=��m��W2���f��2�r1vW5�������d\Z��C��{��#k�Y3���8�ACZs @V�D��oĤv�׳��;�,=��?}>2��v]�QΣqk0z���7���M�\�qo%� ?��%�N�"�:���%�}��M-��	Bl�6���WrֱQz4���}�2�	؂���%�=y�5�l��q9�!m7B�q��v.M���>�2�eU}�+���p�߫��p����,��uZ!��2
��Ӵ8������J	�#���RѲ�7r�R!���Qxzڥ/�oϾ6J����o�FH�QRYJ�sp0[�kY2���I�� `ô=���K�"�*� *k���O���E��|<>y
r֒~1���R�)By�N]�C���#İ�}��6�0�B�5q�����C���eO��=
��tP��H��4�c\\�	��R�~�âi�BQ"����6w���ǰV�ASR�gGH��y�a��/���,����h-m�;{��"��}qÊ��5Trk�m��f[���N�>����sژ�y�#���֋��Z����G�ؖ(~g���b��6,=��EШ�5�y6cI����4�ᮌo��W
��]jP�3�U�k�"w����<�e� �U�������ѓ��\�Dފ�۱����M��H,�e���������6��i��Y���{bLAg����8�^�hZl[k�d����?�R��WO�v�qj��Qh2���uB�ܢV��>E��j��f�����ސ
���}>4}�E�Ҟ'�WD�'q�m?h�$��5B���=�,�.��zX�zQWfӏEʑ�����ѝX��������&�Y=��JˊF��mb�ާp�Ss3���L.F\���غ�$c�n������#4v�c��o�R��ȱ9J�~�F�+�\wb��Zʬ9 ��$�[C�y6n3��A$�T5�&�Iu�99ٍ�'��x�l:Xu@�J0��^�_f1�C�ۏ�6��cIc����9ӟ֏JH��9L6O�S7�הJ�F'P�Vh����*�J���LѨg.��&�epHm�kj�,h���$��bE#:Q;8�bvU�MTp�/��qL
�i1�� �@�X.���/����=��<nz�	Lt����}��Q3���}I��������"����l<70*N���鐝sy�@~ٟ?W��#~�3^���ozG^#48ʅ� û��Zd͊K[j�Z	z���Dj�����e����]a��<�gzg�Ρ��q���^�(qǼ[�vy�c��B6
.3tK��]�1�*���|����@*O�s.�(��<���[ܛq�V5�ӝn�N�UI\�je��$�LN��A��Y  ���e�UEFMz�bg��"�F����$��8��_p�fWC���ߗ�P�}~Iאjߒ�k�[�P��"ɟ�r3]y�8��w������k��]�>�}m�nsY+�~�2�`928#7�(C
��o����ب�Na�_O��q��֯�-m�z��_�X~]d���;i7^C�*�f$7@�5����^ �^�����%�ԍ�#8B�T�a��[C��=�^�Ö8�)����ƺa'IQ����4z]�n��l�g(�ׅ%TPe�6�E�E���z�74u|c�GPYM���kd�0�	iI�O�tV�t��oL��:�<Z'�D/����_Yo)����&��XN�V��Y����~c�+Q�[s��g�{>�h�;n���G�c���
1z����ᄧ�@���8=���6����5!4bv2�x	��;;:.���;��rz2�u��9�huc��/���ӣ���J�)��h�n�^��J��I�99����ZI�  �� '��3��ڝ�ة�J�e��0�hm� t�P�J�(�R�\�U�0*f|�%�aw]�3�n&8�D���"�z��D�?!g�U��{X�4!b:)O$1$�c���[|҄�`<*�,7������r��$x� :|�)K
v��_���487:/�%Ș͆?X�� >���ߙN�֬U�ɇC�J�uD���v��Ģ�&�PM�Bݼ�\薪	�ȢK���SF�+OW�Mx�v��|o\�mK��L��x�΁A�N1?�+��{��l}���2���Mt��Q���@��[�]�V�o�:an��#E792��_���s-�m�o��Y��5f
������˗�"������ �����Zɥ�At�}�p"����JZA�r 2������N^�2뛡�U� q�mARZ&�v˜y�ŕ�)B�j�y�4���*G��˒O��"�����иl#�>�F-���������iM�d�K͡�籄���=���+6X��8-��p:<,�o���Ҡ�l���y��S˄�j�0`�.a�Ǧے�U�Z~s��.5�	{_	�V�>��Yc-4��A���������޼ �ȴ�[��ұ��.��:��-r���=!/�_�{�D|��ϋ�0_���ܢU�(���o��}}�-Ϗ��U��,�΁]�Ed"�>��J9����8?9���?���K����V�)�nCP�]Ɩ"�o��%�c���3�����.�����N��^�Q�Bi���b5Z��
�"4PZ<�ë�`��D�w0$= ~фݵ	9�pփR���ڕ�B���9}�8W�_+[��%�G0��K���(͏�B���!�j�mg#H�JU�4�o�	�R%�c"��F����J0�a>ݹI��ĤGy��**�� |Y������&e��6�߂7�	��d)h�&@����č�2�!20�t	��U8v==M��(DT��`�oY�&��(6w���j(X��)�eO�q��#�jg��"9��E/dx&Ј�o�K6��q���zV�Z)��n��K�P�X*�l�8kB���{ڲ&�@�q������0���,h_R�f]5n�u���)�YݦuJe���>�ۡfZ
f�l{�8��N�L��`7|!j@���|��wQgf�|���Ml8Į^>em�}(�#t��(��P�-����遇��*�&��
�_G����=ɘ
c(����vޫ���H���zu��lGOS��/`��a%�N�l��'~6~qC�j�RB��Y]I��K�CSR�hq���iW��J��:��(?��������y��L&��@M���"h;�˛�G��������­���m~!{��*16�ֱ� �C=�D1T�6>4�y'�8ɋ��,���W����n�툏U�jP~����^p5A�j�$��)Ôf���|t�d���t�EZ�Nl�@��۔�e�5��K�3u��;�a�=゠�X.��B]^��7�JSҀ�i���)F��
�8Cn1�YRם��;W<�|�)1�~/	�K_%�[�Y�pIG�Y��!=O�'mA�x����7����C��k��xJr'MR	a��}Y2)��G���
�֕�9ghG���a+`�0����{����P�0C�}��[i�>���I��]�Z��K���4ب]`� x��t��*��a�j���/��E�RC�4���ݪ��3 �����ئ���5A��6B��A�UG���|po�ܹd={t���hd_�1��b�>�S�����wVn�����y�?ٛ@��y��]���X����X� �a'��D@f	kHع=��P�j����BVD�`Q,#H$�<<�������i�������,���5���G���$݆���;�AWm�1nX�Q�=c<�鋢�vd*��w�={��19�=jg���x�T#uK���gT"!��� N����^�����=	6�Iγ��{���&ڇ�sD�Fv �Q(�;ٜ��@�����ib����v��m���ֺm7+��5�5�̋Z���p�x�����J�5�#����2��qzG�2A"m�ޜ��=�Щ)m8S:4�JV���go���,�ebY�2�!n
`u�e0�η:G��Z����J,R�cuՔ\]��.�bz��g?L#�s�I�n�ZR�� ��m �k������D��+È����$䙿��x�E�8 d%�q��*���4�	�X
[|�v�uW�v���)w?![f��P�'a�.��iO>�\��cf���$��׃<bf4�]��nQ ��w,Ċ>���"�˦Z��T���ثE�iZ�؏�z���N��Q*�|X��*#���Je�۟��^�DFZ�YeK��B��Xk,�J�f��zY�3어���ծ��u�9�[��0_y�Q�Ƣ���R4��,1�R
]�;m�b ��Rք����ϐ�c7o�N��.y�צ(�R�R���#D�$#�*�7޹�D�q=�b������a06������s�Ywd��0I���.=�d^�aڅ�D�$��W��_ +l��^�(��I�@B7�Z���m���;I�4���S_0r!�{I���e0!�{ �o.�^�K�A��?H�m�$�=P,�I���1|�������{�v_�Z	�����p���~�5��^%��D]��@�^IҒKcĖD-rȰY˺�Ֆ��L�`��H��\c��b�M�D!�#�)�t�����sM�1���h}��	�Ȉ��G�����~ʌ��K3�MG��sy� ~̲��	�D�?j$�!�y
�3��_R��ǥ�^�
�լq���W���]��0,��~M1c��}�k^4Q���!�,�_��z'�+)@+�ۂtk����d&��P���y0���e�+�)˨���ŏmO��Mq��"j�u�+.绾����6�Z<[����7�'����M���3Qd���m�`�Q�&M� j��Z\O��C �:1̊T�XXZelQq�X��w5c�Ov]� ����x�|�ʋ	o�X�+U��s��*z������ҍ#��\�q#x�(�������T��,X�?��=ؤ�?�,&'��$�g�}�cB���~���c���p.Fc;8�������J1t�Z�f&T5��G�'�'�1e�ڷ2��[oSe	�tN1��d�!;�Ao�Ɵ7T�Lc67�6�VH�ْbs蝙T���g��O^�[v��d�ɔ��-ޝr�8��U�L�p���9�]q^���I��u;#���)���ϭaҡr�����#����(�@�59ȷ��������J����t>:�G��t�C���M+A8�8�r��>���4��M4E�	�GE�V$=�b-��ce�(EN������T�*U�L���\Z�k� δC���Hrޏ���89�鵂q�� ��C�z�C*�����r�y4�7�@q��GV�cײ�M��ז���^����&���Ŋ��"&	4��Z=醇0�rT;
��2�x��N���d���b�$O��'Ջ��������F��Z:V�U�N4L��N[������qЯ�9��!EM�o�eX$.���yS|?�<!"��dD0���O�O��ѭ�5�bDCko88�}���i��U4m��z�/^:�t�$��W�oQ�C�7���N�	�1�(���po��(L��IB/�Ь�S��XX� ��)<|=����i'��J�NJt��m��?�nxҔx����!N�Lu�S��Qz�vń�� �۩�wҮ�'��[P���TRu2��DrF�Ѝ65<��Tَ�-9��&$����B�[-Ѿ8���]���ޛ��,1HQZ|'����^�t�ly�Z�䋢^
���{U��d�\4����ڱ��N^�j�ɍȱI�-� j?�ߩ��H<�;���19h�6]���vǡ�,���]·��r�
�u�G~)��{�  0���1Ⱅ&��5u4w�-n�F�����LA4g��	d�7у��˴������o�:?�?���5�]��i���o��wzXB���^q�%S���WX��X�s8a{��@`���$����ҜY-!���"�}�.����9��`@X�U7'	v@s�g��&c]�@�{�{3���?,!�0�.��O	��m�_�d�:��������{����ܦtlu�YՍ��	֩�&9��/\l���jb6E�s��s��OD��yb��JVO9���x���?]`�-�~���Y4��n�}2��v�Z4��I@N�31B�PB�	��d�/ i�Uo�,���sn�x�n�{mX���#
?OeܟC�pbK�Qδy#���Ŏ� ��:�6���k���e�På9�����IL<t^g-�T�2��\�ƫ�>Ű\�;�O/�/�BE��(����6+�6��,@�/3<�vi��Ce�ܱI;O�ŶE�v���~�����ЉOp���Lm��aB�B<���O�@@ͽ"��5l��W�����Y�7_� �{Ù�A�F�iMHr`VPBC���5��-�S���f���r�c�`�B�oY����֓$@�Ck ��ʚ�LQ	8چ7:�
���������¿�.h�Pv�gc��R�a,�߷>̓�-CuPfи�F+��Dߞ�_@��2͇�������5�O9��j7k
t�X3rhJC�_ D��'5E�}z�Ш�6K�"��2*:�o��ޡ���`s棥�5�q�^�>�1�+�g�-��kF�iFd.���J�H-�͆J����ŬL�Kai�̳�'�<��L֤=�&v�D�"�f��hu.m}`�����H�Ni�Y��p ��fM���E�R�bG��p�7V��7_���?/Pp[�����D��ŋ��������x��嵰ŝ��c6=U�d�Eخ䞛�lsΣ9�_K��*�9���NZS�����f-C|�ld���z��4"�ҭ��9�H��ސlT�1 5(tfZ%>�&7�ې3���lB�F�?�&�r�C���b�q��1x�m�p��%������Y_D�$\3�\j7M:r� hX*���ѯ`Y+8+)���k��%�}c�܌���T;�'}�O&�f�;a��G�J;$�\d�"m���4��[5�T?'w�U�E{p�m�+a���<~�Pr�p�$sEm����'>�
2:筽��g�m�Oۣ�Z��RE�X(�;V_���2P��u'��±V�/�jBl\�(���c� �0�Mo��Q�7C!�m�C<Q�ɐ�9���uH�b��6�~�j��R����L�,���k�	^�V]V����rj���A��n�Vў9���@gH	�T<�a���:CL��2�@���#�F��j�V>Dp�7�9p�����[�#3�?�:#�$�ö���xH�?ǉp�ņ�@;Ć!�@yw9�G2�y�.����lV�4+��%�<-�Gd�P4��C�<2�~-�ͨ)귰�qe�צ���e���U� ;��Νb�g���Ȗ$잃�����Z�t4�s 8Z��?AQe,�A���2���p�~�p�m�6}ָ]<���&�\�W�s��c%Hj-|d���>.Y{`z�RR]��]*��]�		��3����uq�^	������4L-OO�)}��H��=w���:�@��YwS������Z��<9n'���ZPԂ�+|nC�}�:C�=Z��'9�$���2�%�� h��"�z�Y�-a�d�&"�YD����CI�>��`�x��"U��u��b��.��,hQ����~�8wѓ�k�����9�7��U��J��Sh-ST�����#66c<����� ����|«a$\nU�@�wn���>�%����1N��cK��������.�����X��"���02|c,��y��	S$��(���އ�a��H�J��W���E��A$'�K���?�Ǥ�F�K��6�"��B,�y��ˌc�_���C,X��+3��Z���)���ZZ��.�`}iƧ�Z����]��/��+�jLu�F#Y�hpi@��Σ�5�v
<n���*���$s*fD�8P�+��Dhr�D<�2ao!̨�qF�_���ʠ��D�/G�R/�NkA:���U@ �W����ݱ��e��umxʋ�p�+��͝�bp��ޞ=��؞����𦝨20��NHa+kr( ��d���b�fTl�[̯�%�#2o�'N���F�T�zP�.�t���������q��H�]#8/�=p�R3{P� �ؠ��y�\��;,�Z�
��<6.��tsl�sk൴絛�Ԛ"E�Č${�ʗAp	ߚ��Z��������$C-Q�i�~׶��b׈�<�����#�����X���r:�\�
���6�k�Jކ���ò��xW�?����1�3�u}��?�5*��is-ѐ���ˉ�� ��y�5u�DȬk�Y��ͳ�F>��B�i&�J�~�?��/��U*V1��}��1��-צh�����')>+�@
�����V���Q�i�����R �A���)�:;:zDɋtxZ}��:��J@P�� ��vpGc�ͳs[���O�1"FP�*<#Q�i����Wxx)l�{ˊa2�Υ�;!K�nD��M��-�ɲ%�T ��tU��@ ~��pӔ~���Y��J�i���@��@�`1��p%�N�"�e��+m2Ȅx*�D�{	ʗ��F��9�k�C�>ݻl������N$����8�F�x2w��A�,�3ְW��T�$�E:��UE�{P_t�rSw���쒎eK;C�tk���Ju�%�(~pވ_��k�J��.�y��'���y[%H����2��a2U'95e̥�ӡ�}'�x��w;�q���_�L+�8���
�u��|��0"���Y�x�\���&2RDH6�9�?�N_N9]k����O�N_(i7�PݩkV�ޒ�Q����g��S��n^M��ӂ�m�������2
\��9�#o���#L�ũC��6�х�6�c��\�+�����LZ4�y��R��1�|���[,/�����z^�u�c�UdI�êw��H�7T�۳ߖl�ժ���}p%�P&[R �P�g����%P'OЏ���%�sH���Q%�\�����S��E~4��O�
gW(���Ɉ%�;-Np��{�T幇�7�0��Q�٪��õ�DB?� �Jl����Wv�[�ia�R���s�Q��L3�͝���V�[W�vx�G�Y��4Z����.�oV��p�s	2p:�DG�G-���&�����p�>{���Q�[��4(17t	�d��
Sؔ�бf?�Y�ɸ�Y�Ji�a]�~��R���;�@�SM�׿�}ؾ<Je�'e�Foh�@��8�tp(ʪ��9Y�o���~�����}�Y�����(E<�̐����}歰�ʢQ8_KeO2
cH��0�C|=-�¹�[nS�~�6�����0�jQ�f�ݲY#6w���:��Á����k�ʛJ�Tu��@M��%���i�|0H�;�$"<uՂ�8<�߇���_�:��ɽ"���~*~~��O*S|��}�s�>F�����,���Y�'�7����5B��i>�|@ b(;��!1�c8��4�j� Į&xsJO��Y�p���� �E�$���k�dr���]��)mb��Z�z���T�Q�V ��[��k�n�ƣs�p�t΅���8� �kԁ5�J@Ⱥ*ٟ�>��*G) �5>���ײ�u���QA���9ӘU����� �����
6	 ��	�Oΐ�!n� \�?��A��4�T�z�.��0uPw�
�y��E���j}�2|��Qf�1���yNe��>��͐(�%Bg��wh�[�o�&��n�����6l#�q؋��]��p�sYYx��"���jNP��Ԧ*@��������}c��
�q�@�"�D-&>vѼ���Y#iV{@�K���h�bq�j#g��7�뉫v�r1�
7�vD-L`�ģ=��xa�Z�1��5X,p��^������fw������E�s��jH���	��W?$\�/B���ۯ�����m�#�����}R�hJl���2;GW�hQ�	��qƵW��AV���z) �*S��=��&�

�E&F�����(t�Ur��L���>-������T�OG~�!���TmIR�u�=/E�)�峹CMI��:�e6ǔxl���� �K6,�����5�@?d�V�˶G�3w���?��Igﵘ����h��-l��ߎ�/�
��c7����oz�"TX�F����^mJ4qw���)A����E5�5���T��P	��vH�k��Vge���O��{)P�E*1<0�(��t|�.\:rP�?���&�7��H��3���a�tU�*�g�E��@��e%�ff�]O��a�6�ڛ�)����oos����`���6�(�A�UeЄ��'���%[�7���b��1��R$3���a<��7�&��*g �$�
4"��M���oL]�ٿ%�y� O^�Ւ�8Ft����@���7���n���'�.ч3�d��}�����0ls�?�~��5�X��j�7�էcbp��O��3�:�6��m`�.Y��OXw 8u"��~>�>�^��Cg��3}����;w�ϧ]e��]��D��h�K��)��%��e��t��yS���i!�,��A`hक़�v�pa�Pݐ���3;Ƈ|��.�6a�7�u��T�w�hu 09ٿ���֓=պ�
�������TTY�i��X\��8�P~f�/���$�A�X(��5�]ifN��sz�s��yD
��l��K�>����椢��!簱�~)���B;���i�ʜ�:%z��Q�Y0?F�WY�W�G۔
�U���N��h�~."L�K��񛾷[��Ө�;���u��,�eT�υ���n��� m�<O��]�ذ�+�L�ڧ�΃o�E#r�ʸ�<4������rDX�C�}N���� �~(�:���*ɢ�3�pC8?���_D�^�KWCS�sl�f�P!���Z�g������psW�Pa$j��U�]�^�x�U��g������3�ێ�xY˽��"s��S��k,�<��6�����mۃ��U6�R�a���H�����@#e<.�x \���9��H���v��pڹ���a{�s��U2h?����j9�+Ǯ����mc���=V�0\�_�Vf��T�Wցx(-x��]niN�(
/ݢ�d��k��I[����N�r7��*V�V\q�e?�֪�3�	��ו�ݾ��ͤ�A�m>�R�q5j�+S�yЦ�(�GT"y�V�l<2X�A�$p�r*`�΀��| ��@���_�O 58�hvK7�o�I%�x��>�*պ�.k��^��夿��F���Gd6L�	B$~J�҆ǚE/��;Ғ�tI��-깵��^�C��0$�ZLN��K�߽q�j�������*D����?��T2�W�#閊�1Tbz���D��Hz�@��VFI6�q@-�0�9�ʘ1h<!<����Rه.��) b��99B�Zn���:_	�Ƶ�U�X�w����*�х�;^��,��Z�0z쿕�+���/ ���m��oJq���@�ph�)�=�7�=�3�2���R?D��-V��{�H#A�xm�t�N=U����64��,�C�)������E�Z>��O*�xڠ?BQLZ��5���3�7�wN��#}�oʁާhpJ���
C�1K�3�t.:4�d?g91Z�eR���b�ȧ|�;��ֆʖA����Z�/���`���t�(��Þ�Zb$ʲ��=��,v|\�t��=f���Z �p\q�FD��"��֥�@���3�։����QxY`%V��{J�����1f�^���혋�#)Qtn�Y4s�ħ#�`f�NNc�؋����Ȯ��5S�~Cf�h�(�+Gq���29v��)�d>���R����2��w�0)q��r��'�
���ɕ�`�N��(u�x~��ډ`��ӵW��9T�H93�g*5\7(�9k��I�KQ3�a~ɢ��,����k�!�[���N"��إXyp-�a�s�gP��+tl�˪��.~o���\}����U���6gU�az�u�Ia{^,�c`UWvt��vl`����[�|&uG%*a)>������e�h��d�D5�V�th!a�w���3�&F�>"�|�6J���?��×f\��ѧ�vd��V��C�(Lf:�9��T	�~�J�zy�ݐ���siޠ��z%����*s��J�Ī��
�E�����Yli�S�Hd��~9��w��o�a��QN���_�n��-�t9E�f��߿𦔞N2X��z"��Z�}1�����k߃ɏ����Z��sZb%���A����1⧏��8�Ǧ�����ｕ�ykx��d>�m���}�����s.�$���!�ꈻ��!�UwE��>an;��#	��j��&mS��χ5�x�D�y�V���������\��-z"R��[�G��9T��.�͕������zڌ�T�[��"z���L���\#�1&|�1�yՁnn8BAcQ(E-t���?q�O|��G��6ݲ����Xھ.[�kvx�g�m���a_h�L�9*3j�AЌ���D[�����rǫ��2����B�O�N�z�Q���t=c.��U�2j�CAt���b)�L�6C�i����k�ǜ�b�o��/���1)+�99z�]k~"������㸸�mٕ�<8w��݁M>��Ǯ���8�Zݷ"Rh��h���7���#�L$5�˩3�N���������s!R�*`�AD֠~`��`��t�I���n۶�=
�z�U{'�愈>��x%|R��F��KT��n}�&�]jy���[�Δ!�S����^
�a�F���AƠ����|�{��P%��i��?	�w;Gaߠ
����Ӡ®�?ov�Y�$�P����e���H���\MK��_9�W[����v���9�忻T#թ/Q�me�9|/���P��MѸ,i�ă���NJw�"<yN���sf���6	�.#�v5�Ҁ���1��q������G�8�Q]G*+������g�Q����cv��js��~Ə	�m_�:/�4��GG"��M2[F�^_F���3�� �P9��8��Wg
r����%�qc��n�L?�v�-��hщ䬤V�f3-��k.�3W;M��Wn��m?�m8��� e6Ii���^�S ���!�dϸ��Aم!�{��ӳ�_n�O�!m���DP���\l�3���H��L�&܌���@�j�ByKY�g��|p�:l��!>���"!� ��y��^k*��gR�	��l��B�
�t�c/H"n�`�<�u8�d���/�.��,[ϥ*~T73%���'58��I.H~���jL��g��*.���U����Q���}�*��u.�P,;� ]'W~P�s�4~'���6���s<b���m�L(�{sq�X����cJ��t���k�a�;qc!_�5����PRɌ������:T�����Zw�������E�N��Ȩ�����؅Am+g;oL��_k�������s���罎�p�l���)#U�#{�QFC���b~]`=��}W ifV~�폩8UV��HөM�m~�Z\h�}Ɇ�]˯ɲ��ɼ;ץi;��9*D��X����q�9]7�C���׵���N1[9��Ӽ����?���=.���p�gn�F�./~���K�-���v�.����j|eJp��Z�`�c=�>R�Z�%$a�����������W��)����Y���T%̢<�C�KA��&nO�PQ�C�W_¹�m�G����N�  ��}�����7�A'j��桛[E�&��V�E�n�`dG��\o�K��1 Y���'�Dd���;֦4�����KԗJ�ۂ1=�du0Y���6��@����qN���bտlv�u	�J�����a!3UO�*�XY4��)�{�ҍ�'�Uһ���l��@_���-JZ�L���jk�+x���>�~Γ�n��)�AШ�^�1�&���{<ڀ�{�����͝�c�e8\T�d�^Ö��H��u�=����T&m�� �:na�km��t��3y� 
�~V��B	k\�i��-0�@�=1^�/�/N�_��6��C'���c�*`����{��(#i�/8ˀ�� �������ݸ��Kc�k�歫ۺ#��=��O"4��������G�|�U��׺|�bu���X;T��8�y�ʪ��u���ٱA��������j����B��`�3/	p&Ġ���$ ]��|^]�U����W�~�-�����Z��g���㕂�K��Bbz�ìwu�x������U ��n�oG�l��55�!� 'V�X�y)���N=�d؁e�Vn�����B�v�)!����GT�`_=.�n�\� H�j  �� ��>��Z�+�@�8y~�4��M19�K����ʘHX4�cF3VI��ץyJ�t�a|�!j��F��/:>]]V1���������Y�ar�(&'��h���9>�Yֻ�r��Q�9 %���*�s����u�?_�l�A��01���P��%4�)�VN]rl�5N-����4!;��Qc���_T�t�()#��f/�I_KDg��t�)��w`���";�������D�_u��o�4sc��:zK;�<�Qy�D�L�pק� �˰�gKs:Ax���N���+R��u'�B~M$J�ɷY�Tjed�04	E�:��x��?�c)H Vr2:��S�E�uG�+	ð7�G���;̌�l���I��'A��I����e�|�=�4����SM�Zu�_��r}K~� ey�ip� h�n&{"g]�5y	ik���o�m�ح/�t���_��N��$w��a�q�9yDaOv�@i�Ÿ����=Sܼ�{�\�d�Sg�<�FF�b���;����]_ɡ��������ӯ���0��e2F�O-�
Y�<���i�EYe��0�����<Ge=�;�7�3%(�)�i|&�ҊпY��Ӗ�z�9ܼ�� c�a��Me_�rL��rTrEh��*�/(>���\I��̖�����]��[���Ί���הKǁ����{]���G���RC{>�90w,��?	���|�䲶#{��-IW�(#H����e���H�m��(�e��De�>�sW)C���k`�߇m�z�c�>���#_Y�:�$l�a��z��߽1Ķ�x��xh�!X���0&�i+	�e�nW50���p�@���X�j^{M�r��xM�"ҿ��L�y?n������q��NC���m#@c{�M���5w�y����R��&G���Ʃ*o�X��o/&}5�-mrA�����vG�����s��4�`�ި�-�w�XG����W�6 l�	��|p����c3�)�� �����V	����T��B��U�t;^å �s�n��ª��}6������<�Q�f�ˌ�7�w���|r+�������x�+�1�.���tFw�D�iQ����-�PM;��^�#Q��Fy�v�`ڗN���я��Ke��~�{d���P�/��	}�	�!f��2�nlk(W@�����#���T�К�4�;����pW�'�����������;�3�qzBhoR�.k�<�&���,�B�&.7��E�P|h�̼[b�����B����C!��WΜ.h�ٴ�Bb3Ⱦb)�^�,\_3T����7��y~G�U�)[��R����k����s5�?�x�gV�7��F�QE�=�<�ILozy�?�ʃ�!F8�(���sfq���~�{��p��̱|m(!PsŠ��S��Oř�Gb�|�u�T�X��6o"﩯�s��q�[����dj����
���7���O!<\:����������=���.T%@;�,�1��DH��k�������]�cz��]�h+�B�o�Ҁ=�0M����Z�*]�Q��w�s&�p*|w"���q�.�&[��E�B�p�o�ŬJ,- H��ǀ��?�nIu�cќ�(wef!�ȻJ��B��g|>��-�'>�A �X)�F�ؑ������q��c��we���m�`��Ֆ����㘨���\FV�lV/GNy9��k��S�h]�Q}j�m�T4� ��tn���Rn����-yp�&�Li��()]�7��^02˳!wH;��A�E<�J��&�E�����G�@�Ee�� `�/�����d@����c�|�aF�?�J�"����le�j��U��w�9��u�>l�塊q.)���g��¾uMN����ʷ��<226	���fs��V n'ne����;R
T��3~����]������9�.X�l�Ѥ����7 ���aI�Ʉ7IEmoȢ}mTf�n��U��M��t	^����jhH}�*�?X� X%�}z� ���TCp;G�rq��N�����0V��	?߸�L���.e�5�����G3AQB�O�Ti#�l��##��7*��?�c�/}f��^��<�J1JGD����\4T.T!�@&Ui�l��Q�⃃��A�V0w�D�&WF�W�X�6w��Ӛ����r����K=�7XT�P]�� ��>Hd�������~�橕hܯ O�/�ҭ��si�}�v��(f鑝��p*��l:�4g�D�W"-	��Dz���.ģLf�
�Co�B�k��˽��"O�(�#\\�����Q�t�g���zW�&]J`6`�V;�ފ��6����z����@��
�e#{f+%����;�X���?�^��ת�M�[7�/
%�X�bظ`�t<in�{`�������s��hU�Y"�Қ��X3��Ne�������/䭶`b�1��d
�6�b�i3���(-k̒�=�̘��W�������㜬?��|���;]��^W�h�7�C��`��`!��>�[�.��)�

=B��
[[\>��,�HT֖�r j�L��Ww3����5ݫ�d�N5��>�ۖ�:�iդAnn��<Rs�4%I	_��)t��2ll%�n%�^�l�#?�31��|��~��y=�0#m�u��X�BV�H�Uθ��U�!��H�z���Ϊ�����������ƣ�-cE��.��"�0�1�m)}�Ul �Ϛ�� b-4a���d�S3�������&+�����Ow④�����>�ިyH��!Z&��b��귥
$j�h�T�QG�R���c�:v}8��#ܛ����d�B�{�pu�u��j��R�ت=!wSt�;尋������^��W��G�vYF��	���|o��ev�G�L��(�A�@��b6�9YU��|NR7
W쁵�E���Z��?��(�(�?�-d?��!z؝��etC���$�+��q������ _Rcd�G�a�:y'(=�����է�#�j|�=k�4`����Y��s��?��3W�7��E݀]�7Lfϵ���[��z�2�K�M/X"*���4�b���ۍ��2�4�B�,�9򑇅&��?������{M:�6�g�ǿ��t� �!�&� H��l\_�,H�Tqܥmf\-3Ng�i���9�Dy��X�=_��g�+���t���!Q�vH��t���#=f��-��̑�-�ڠ�������;�f����V��a��N{;[���P��T�x�g�0x�q�� amV�0ڔOa��S��iPj床x�z+���}b��9�rp5�Q�/�&k��k��	(������R|`�p��$��f)"t���So(��g��`�ַ�n�:k_��h���p��J�h��O��
����m�˔r�&f0�&�R&^�U�n�Dء>��@�Ct`��� �����Ɋ��O���M����*B3�!�W�s䟞1q�?���a[s�<rܹA��.�#�6��s��~m��c���s���}A��[��,���Utť�2oQ��dF�_�����6<x�gf�W���5�H����O7�"�wO�+^��2�M}�.�����M��h_�C/j�V0F��Bm�#�s��`v�V;��
���~}S	Sg8��o���w�i`hW��Q3�b��!��pg.��]v5�	�wtY��M��� 1W���Զ�	ڑ�Q�*�8�M3�y=�}�EE�~���T����|6[n�d|\p7V�Gyw�5,� ���q;��Mfdh���݇�d��%5���AɂQ�S�N�R]
�����&-P�ڌWQ?}@?�P�9A	0�1J��/�l0�޸�ڿ�,`㒲�#�y��m�j��||zw�(7i�;XZ��
� _"�ޔvb��#g�@>�u�e�6��V���8&+l&�p�S$pj�r)�.��J�;�0F���i�Nh�A�z������^g.���[wH����ظ1f�D�W�'[M��L+�ȩ�s���jD��fZ3��@%��*r��i�k���wb��w�;��uW'�)��x,�*�ۃ�r��\���3������,�l8�����q����O�c��Y�{�}�>h[2��U��&~�sp�	[�c�>�f�@"ͫ7"\��~]\#�;2�QG�a���:�ܛ%�����m�뛱���������MOc��Q��:]��Dpm�����lJ�+��nڭ�8B�v!L%�=��'Ѕ�'.>�V;��g�D3I#cm�Q�´��	�h[��r*��TF�)r��W�?+G��I
�/ڛD�!=��PL�����G@ewV��l��\lF�d��.w���Slk�<��u�����3�lU��9ۊ?�#��'c�e���,P!W��j�ghfy�쬷��@�\LE�7|?Y�����k��Kv����=I:܊�Z��)%'t
�����&�n�΁����	ⷯa�9�+�	%�8�/�̶���&&?��٤�G^� v�e78$m�ۂ��>s���8C+T�e��.k��������v��sZB�J���gX��G�n��&�c|�P��eM�f��.װ�B_�Q�q�H��yդ��)2<h�Z����y�����š�ƾ�c�6
=�+'�XF����'o��8�mfR�h��56���}�Li	=����<��a�rt���v�X�$F���0��`ת�l��u����#3�ʒa�.�5�T]�E6��nR	(8�A�j��;�xLd!�[Y��Gэ�d��������?}���xU�v�`�/-�K]�T�����9�B��3&TDHז<Y��F����S<h���+"��B}$��1��
��Mj˒t=66�	��,3/dER;(3X��
�In����L:
|b���B7��$`�Z@mL�ꎢJ��čs�Kg��.�K�T�ySs�W��O�Y�B%�p3����$���]qF|�k�/�gȋUE]RaK��΁�c¿���97,�����v�mf��w�+��H��YO+ʛ|S�f�s@0�=�}^��1����<f,�y�^�§d�R���d�U,��a�#�c�����	).�=��f�+4\�߫ ��X8�-�8l�f�?����	������a�ъ��X�r���Z�\��|Wt	AYwpF���Mk�B{Ub�n�f\���5w@~=�2�W���H��G��F���˱��$K�z4����?�Y2��w�����U�����iG��N��LP�U`���?�q��=k����9����z��֜�Cx1O���x?<F��H�F��k��3a#����k�OyO���)EL�f[����:p-����3����P�=�4ᥡ7!��O�cA���fF�pʗ"<�[���w.90��G�fo�A��˒�����X�=:& �W�i)�k��cujX$�܇�T�ws��p�W��͸*h�ݓ�R�D���p�zʪd����JM=-f�J��?�~�	ྏmc��VO���|92?����@�6{ͧŧ���t����,I$�ik�0Y�:��╩]��x�"�2��3�	��s���AF
�a%�� �}����ef��bH�y:FO�_�&��;�5}�(��IՉA(^d;���p"\�1�`�l�e���I�ۻ����GK!�
�Dd��g��aƀ�q��d7�a��d�*�b"�ȿ�f�}�8}�k넥��Hgr9|@	7�;=@8�O[��v��p��
�ia!~I��ͦ|bN�(��j�ǈ��h�j��-E�,#��Ҿ�v�����0>�کt��	Ego� /��N����BvrRTa/�I��~D�@�����"XW�^)�*����t�p��"}�!"�[F��O�[u�>bhk�'J��J	�+k0�jJ\�	u�Ϊ�%U��	�i�s��o�7~JT�gJ��^J�V���k�v�&mO ChæK�er��)M"��<��L����*aps�l��D��>�[��M�L=@�Mо�/e�Ԛ��DWY8m.&���|�2%bw���v�����i+�bL��߰���4����SH�(�j��@�ZJҨ�/*"��������-w�c�)�,p��f�T�	u��:1��=�5/�A4">C$�L	���rj�Bt��H,�׆�C1:��� ?c�B�T�"�s+zA����\���=�%0؂�g]���;�w��y�"��񓮪����=YS�>�A�t��V�ň��L�3��d�;��g���oFy;])� �Q���vM��ߑ��%�@���߯��ｆp�`Yi��ꋋ=��"�+��	HV]��;��������f'�g�!�
�ǻ�!�R�#�i~0�n��O�����
��� *�J~�~~�,���CK}H�lmAM�E�n���HI.�p(���`��ux&��-&g�����O�	� �� ���0q�vW�x��m˹1k]�S`֊`w����`�-\ �)f	�����B����3��с#ϴ-M����t��\�����nO����Ā��FC��ߑ���;�H��*Y�A"/�O��Q������?8'_L�>��Oδ0��b6~LД,���0�WU$malm�����6���r�f㷫އ�t�وe�lY�"w�����ݮl�����r��A���z�FrG�qY���r�(Oܗ �j2)x���L%�PR!��A�Rt=Տ�s���4ԯ4�L~��A͈���;^��~K�5�;PmtːmV�ͳ���
��>�%ܢa��#���s��;X��u'���b�N� �9}��*ғ��+�TM�Z_xM3�t!Z���_+�n�<���/+�t&��m��T�O�na���po9xM����CL�/�_��J�;/k�)��gh�L{/�NB8���v¹� A���1�E||�*�������Ձ}�`s8���[h�ڹ�řᦳ	Ng�t}��oc%MI�B�(³\G��+$�R�
G�<x�;wB�(<]�	ff���brQ?�����m��㮆�w��C��bDЅ�8ࡘh �Q_�=�df�1�tv��@e�4�@`��"��1��ǽ����#�їa�Y%;S
��ub�������[p��2���@��Wd��;�֣?��?I�1Ȣ�M�+�C1�_~XջP�'1��5!J�d�.�N��������Ѷ�3��L*�bR�;���F�4_�rA_c���Ρk�wR�H�#�3��|��!6�L���t������e��V)V�Y1N�`(�[�q�'���*�%�_��]��%!�wċ͚b��!��������t��Vo��l�D-�LcΒQǎʗ� b�(���ƒ�0���F��]�^b�aR��:Kl�&�.LR�B(gp�l��1~�oN��N���)a8�z�N.�"�Qj���aJ���
�j�7�kD���|���t!Y����&i��):�ؖbqN#���<� U����/̩Ydw�����>��t������L���(�a�펹<�v��2�H-`��>>P~w0�5}(��k�8�,>Jvs'�ױu�n�?�t�w��
�n����ؐ���P�^]n�/l�}>=~T(^���7;NxvU�@���|q$��R���M��Y�uV�V~ȴ�"6���� ?�s��B�3�q�)+��u�-="�v�f��Yĕ�jԯQVA,1���uz������[��;l򯩅�x�u�c�� 2�#8	=h�ε�Hm��!%�~>�n�-RW����}���7�8����6�~�h�{����E��gB��m��x��&q�&uiq>CX��uY�S�%�PԶ�>�Ua�p��!��_`\���%-;��cW�o��_�<��vD�H,�uB���Uu_������-�ً���VPP�����`����(�V�e
^pqjN��֊}�п�]'�ź��+܇��is�T�Q_t�Pe���]���)`�r� ����+�l1��-vS�5\���@gm%�?�F��2VӻP��|��M��0!��dEEa��+��H���֧���	C����������>�������V�\�ݡzNL�\�'�E���N?j#��Mx��͐2"��,��SÑx�pr���{���SwO=���j8�r=]]�"_.�mB��᳓^
���&i�{{�S*J�+22�L�V�A�62Lc�"<Km����r�2���O2qKΘ�H�k*����9l�hݷ���8ڭ��Z��F	b��P�Z���6�O�N�i�����x�}u2�;~t��Ѧ�{��z$��:���)1u-s@q�6�gv���D����L+�1�d�x`Do<a����ؚB�Qu�U�Θ�"�A�N��>(%;;������>[vX�w��=n[���=?�veE֠�
?��UhA�w��Q�*9�%����������Ya)��f�y���̣��)8B��ɇ+$�:i�BZ0<�,q ��bih��Kz��7��T®��E@��eJ�]���߲�?����U��)x��#Q����ն�v��$�B$�#�fB��=2=j���v�V��el��I�+x��S��� 4�@a��Ok/у.
$05|��7u>?��>�'�*$�ջ�b#��W�%�]�6����/�4��4�R6E�e�"�c�'\G�Nm�lD�k�ق:��uX���r��P���!�z���k�΁#�K���J�8��yp���J?����e�(40�^�m}��	i-)�@��XR|�S��t��b{�li4j+Ru��]�U`A0o��79�kh'(}߶�V���$�Lm��ߙ��N8��R��_��f�`n����PY�s�ҝ��׹e�G�}Z�}V|��Y؛�:g0R��y(��N��.��B���Ɛ�=ƓS�6�����\5�0r�4��#�}��K�t1l�-o����t�
�]�W����Nx���S[��`�4��BV��BJ�a�wk�<�Q�O��������_�\C��U��msΝ��إ�֌��ݎ�9��;s�"a^
/�`�U������r���7�q�ݛ�m���Є��A�����ש���ȇ;d  �)>�Q�f��H;�_*���V�d�����Ć���s�J-G �ζb4����`���`"}�'vw��	q��+��Q����'Q�l��=��د�k9���3���r(q���M_X���kĐ{�x�����h���T�3��8��I4.�|�.C~���(�'���M��7��(��3����u�>�6�c�hJg��X���Q,4��)��!T́��u��ۇ�:['��C�$�� ��.����s�u������ =���8�r�I�$$�����JZ-�����NDƳ*�K��ռ�Y�NG2�+� ��]���W�Tv��v�/����.� �j_ݟ�f�'�a��(S�o-���n��ۨ��8���D�/�"�+��j�z�N���}˧������e�A�ح�|~~w��,~U��z+�)w�u��G���~Çd��b0���ں�܀�E�Zj�d�b���1S��������d�:!�ɪ�u��^+�8���J�ؓ};�u�:�Aħ�66*T��Ć&��)�'&+TB�pe�Vߪk��Py���t��vF&q��W�{O����]f�%��ff�v%�2��z�}\[\��Ǌc�n���Ael=ec��4�l<�9�{9d�_Ԏ=�&�<~Z�Ҏ)yYZe ��~��&�0=@���t�|GY�A�ְ�P\�Q���� �S�P^� WlH�y>�1���`�*�|�H�¦͒�Z�/]����	?6a��c�x��W�� e���79q�^���,�;V�V�h��A�J�ۭ���Xr!�i����B�B�u��HAH�K���R���Ias��:K��t�b�[0ɕ�Ͷ�^��k��{1ӵ��q��V�5�Ym��NrΝ����_ET�1H�`u�8���K�p��J��v��+��{q<rj���ܧh>��y�{'�=�X~ O:Sx�f�CL۾2�2��[�Mj�X����#�bB�#�`��7=sb�����ڵm���2&�e�ő�x['YF��Q�}�+�M݂?��D=��l�!��ж���O
}��_�<Y��6�0?��@Kq�P� �Լ���/�߳�SI5Y.�n/ͬ�F-�4�ؾ�MЊ��ES�F�8b�]��z'�Hڂ�+5Ec�ÿ�0T��t�A�P��S�}���L��4[޾�]8�$�S%����Ec�~B�d;0�ͳ|xf]4z�PU��r���I8�%俍�����a�)z� s���dJ
��&�*zE����V�M�lQ͊�g�r0�ۖ@<�p��t]�j�l��_�+��jρǧ0�X.�:����	J�UG�b8'��r�%�k�6�Շ�-ni ��ψ�$��f�%��8��c�C,�6 *� p�}o�|�1��E'��T���ɗ�Y�!�#��>m�����j�Iq��h^PQ	��R�bh�>���z�^���3�u�7\�����?�Sb��"K��Kˤ��,�(��\��+:Pz��ʥ�	QV������[s��"u�X�R�6�-�4͕A��s-�٤@׹~�SL��]J+[�a`��@�2D�˶�kq� tx�#%���UPd��k:�X�F�Ǧ@��K��U��{!������rߪT��'�b�9���vta�a @�����@y��_2"���Ka%�#��n�� {����w�@�_���1�ɋ��-�c^)g��	�ٍR�����_6U��:�mg���f~U�"��P� Z�;���q@�]�&l^��z أ�.�m�F&(����I��Z���3JF|傤��K�_��b*��]�q����vU�]�NI�iL�ٯj�1AԢ�C����L��L�}D��'{.�5�D-�x�p���>��p"�?#KgLA���p?	֥L�������f���?3"� ����T ����]h�
���d;��D���ע!cR�#�Z���D>��a0��e�1�)�����b)�#��,\�]_R|ҩ�5��}IKW��t�S�h���!����	���
$'r�R��Zc��$�	[�� u�\-t%�_�&3���x�ƄYb}�x�(
�Ӟ)j�|�>"�6�zѨf'�w$�s%"{�KZ�16j��7\z��?`� ��&�w��v��V4R���T��r��Z��Ν߲U��ě�6]m#����]�R��$�X�~��ϊ�sú��9��jk�L��{�="F5�pE����mVxR��{NIp)����G�j�\�y:�OOj�Eݶa��?��]ͯ��g��zO��P��?&vY���B��\ͦhf��\����8�=0~hNT�����#�]����U��d�����ZϜm�ԋ�P�O�����s���֣��Uy�J��`p�7���/=���/!O82�-ͫ�)�p�[:��e򵕌ٺ������sr����:��ٓ���C���+%����$H"�^�$�J�����	����wdr'y����Ἵ�@
�=E�0�N�ݘ%EG9,�VEu�jae�k�h�A)��T'�;�G��߀�TJ�g��f�&��)�����<R�\�,0����"W O�Y�E5a?�Jʞ��)���"���Ou(��s�F��n��U������p:��`U����'.L�ID+U�:������b�?Fo����2�A��U.�]P��2��)�4�fGcr��nn����zii��}�A�[���C���P8��Z�nR/�{4swY��OS,kQ�~��,|�jW�P_��X�ۋ�/���}N�ȯ�{�3M�r�5f��w��x��ؠZ��cqt ����a�����ͼ +�5LS ϛ	GH�9��y�O��u�*�c;d�é�p���(22�y���- ��PV~����Q���j��8���tt���+z�����B���z�`�+�(g
\{�e`�(ACٛ״j!�jY}�9�S�g�a�B��W!�¶/M/�1xZա/ǖ1f��:��Kdw��f���Ѓ�&u��xzֳ3oU >�.�ap��!p��!��7�O�S[Ü���� mw����1����]�렁``#�XV\�P�Z
�%&=�r,L1큃;�3̓'�fb>j���2��1E,%�_��aZ�Vf������ڌO�[�X_�R����׈�>;���Re��33*�'K<^A'=�?1FO�8�4m=1�t��J5k���)�g�v~H�<����V��N��C��=
[���{E�	<�n�'k���y`i��A�#1Eh{$����]�(� "��GZ��wNn4��,��Y��~��W-��� �T�D�Z��o�g�D	i�=�a�h���9s,`�g�	���I����ae����L����3��X��R��10dX���Dfs�ϕTGe27_�<Yp�V2�jKু�L�qyE}jb�S~�ɇo�R�GEN��r���PC��Vo{�Ч��Nc`豯���a�=��a~���et�8�*���WUn�i�t�^oDjZ�['��(ٶ���;}��N&j	�����q��mu07[��W��ލl������;�V�J���3C�P,F)�����g�~m=˲�D4=�筡fO�)�-�ӌ��@���j�E��Θ�#2�n��t�#��N�13����X5^��-�L̄�B�@���`��x":ag���jA*÷ݪ��A�f��z�A�,�/����3�A���?e��$��ѯ�A[���~��XKf>F�B��JXqm�σB����kB������i`��,�D�].d<b4��]�Rnp�:=�i�t��9�e5-����.v G[�,��}J��8sHQ]N|�^�d9Uɬ�D��߾�8fËz��E�0�R���2*�r/V\�FϤU�o.�a�f���8OI����>EC�Ȭ=k;��'˔�^��� ��Z]HƔ*oQo��K�����'�i�;� �4ln�zJA�����P��{9�W��v��v1��W������:��j-����#��;�/Jy(U.Td�S�ď_�莝_)<��\Md�ߒ�<=;ib�H�0C�\���0Oڑ=�8 �Q��H:\��*�b8�k������m�Rs��+��,;Ke�:��g�ZQ��4��Ӹ7���W�5C?W~M�#�AϰDe	� ��#;��4%��t�/0X��<b�X�]zh�Lf�5�Y��4��V��
j���ߐ{[�^f�h8֐7��U���Wn�h��p��t��#�~
�k�wUi�Vb}�iI\���e�3̡w8��k)M*�=  �[T�!�!4��-��tM��9��s]�ux�Tm�	4.�h����;��l��	�;����V"�ͱ�<���0�^��7fc�6�S�J:j���b/NH!�8��vB���� t���4C0h���b'�MP-w����H4��~/�J㤵��������V�7kI
)�V�#�?�� �� ��B�a������˶_��}j�ˁ��ڋEUW)G �g��Fg'RK�y--��*%��I1A��:������J��/�,lzf\�����ܶ�!������a��kA��E�c7.�L�,���KE��=����u���_��� \���6��IϷj��������^��]Z\WB���W*8��([�׈�:A�*ܵ�}��MP�n��u����Y��M����?�V�V�-��r�mİ��=I��}���¦VL���̻��,��_��x�9�ˡO�:��Y��eX��Iw1�u���.�jڀb��\��s|`�S<�c��IqR	�;�`�ىV��X�#z�ٽæp_������vc�v���"&� ->e�f���<�q"	�~⇡�k�C���	H�\0%4�+3����VtG����G�A.�/��c�e�*a�	�Z1���cU�fsd��X��8�%o#��E=�+�	o���״��%vX�����'��J�m(^�ZL}��_ ��.̳zW(8���}�qX�.�����"���[ 母���y%ˈ�%l��<�ˋ�����$�?�lx�o��d��`���g">e�)x�,BXO41xA����8(�Y9��+��=�)�[��d��ǄRmC՚�ǃ���Dʗ�T�?Mof�� Zs'��k���1�e�Yp�v̩E�zlTD&�t�=��-���&�m;�̡4� �x�K
$�ɒ~��<9�y��1p�&��;@
�<_�'pa�a��cj&���Z�?�E�H��$�w�]e#ʸ�����`x�Us�P�Ip�u�;A>������\����\UF��]���?v10���c�!�P`�/c�e �8u�Fs��o�<܏r���v�E�C���}Qhlozv�W�Ҽ� �b�Q��f6��������\���5'Kx�!�F�Y�0Y$���	�֩g��s1]Cs�+�U��i`�L��L#�.�����[��j�k�Ac\X`?u�$R�̲��j��T����ɍ�Ⱥ��1�Do���ZS�T���`�[U���VC-i7�c)��M~̽����Ӯ;��%�>ڜӍ��I�C$���u��3Jo׾+S���Y�-,Ｍ0Ҟ�.�y��f�������O�7:�
<擬d�%��D���G\�hAn������˛]'c-P�e)��'ghc��?P�ѫ���P�]$W��9r<�j�hY',�F�D���� 9p�7�����G�f|�:<q�z~�O�}z��ΐ�D	��jSf�=yY�CtE%�%Y/�������ۧN96,�E����r�1h��J���� ��N�^&���#��lOL�ω�S����M�%�z0�k:Z����(8��#Nt�"|��%��c�橒�-G@�nq?\�.���Tkg��D�
��]P���zy'��e>a���nX��i����%J��*��_+(;��vVxI����ٹtꃀ
�4L�O��}���]�*�}*J��m�]��W���O�#��;��(���1��c�o(^-�	_M���v�x��.)���?�Vy�{���w���_��ڬj�gn>z͐��
GKh��!bn��#f[��8��������
���GHkey�٦<m�՝� lO�;[�2�͡/S6������Q9V��_����2�I�}�N�sj�)��:���d���!��;t���`Ιa�t���H6Nl�q��_����������P
�d��w�ȣSfA�&tCFvf5ƽ��bP��Sr��7{�Oi��6��t��>�5�F�Y� \(*B+�N-���>�Tv��_�x��*�V���1���H���m�ɤ4�� �;���֊���&F�<�%����zrZȑR�k_%�-y.��˜��C�L��9dX�g���r^�ԇq�fQ�L����������¬�G�M�a�:x��v��
�B�UZh�N���ޛN��:ަl�r����<�w�7�ܜ���ܦ�, o��oa�����e`��=��Y�+�kj��=����Ǒr��\�_����������_�""�q�L����PM���a㹎:-VTp�di�oD�
:�{�%�
"������4`b{Ԏ[�B1��J��G�؅����c�m��X��ۛ? *8!I�\����V6����N2B��8��&c�H|_��]���EV�Q�-)���י�b_��9 ��ϊ���<�
���EgƵ�Y�� ;#,�]3�G�wt~م͠�ס�Ǥ�02E�5{�!k�U��</��A�ǚǹ�}�`�
�|p�h���3�4&(n�}o�dCv�ܓ��-�D%���i,e��ߦ�H�raVܫ�(@�����5_�,�i�������~��Z���{��`X��ھ���%2݉j���Ͻ� �c\��d�R�M����Ҋ��]7aDO�!��;g�	=	,3"��Ԑ���q��� O��֟�VS^�\p�!Y�w����}�w��=����Y�B5�>��m�+��sbܱ�W�c����1-��_�XT����
3��)"p��%c����ތ $fu�ѕ#���rcx�^:G�Ai|���Щ�M>��_�Hg���%�ް}���߃~�VWh?y>��ޭ;X2� e�CV�S� f�B�p��S#�_�����ԪĲL\u��x�U�|����r�b�/Qy �մq>0s��ӗ���,\�W	{��
�I�������w��}/���%���g:q�Z��DG,^���k{��P���^bzq>�F��!�^�S���Ef�Y;��<&�T�j$��jߛV��n�a�O�\V=��тZ�Cl���2��o�*�����5t��{�GԹ(�Jm'�O󴹳�xL��dVr�ρ���Q���kY�g*��y6�J%��(�5�$�䀁��iX��!��f8-��q�����C�
�����5}�؏�9���x�b��N/_J'��t��U�ט���
 m�q��L#C� ��˼~�:D@
}b��7��;|�Z���}���~hw7դo�s�@�e��#(n`�[2��4��M=��?����j )�E"�*�/��f����N�E���E��=���g��*@^�a?JG��������!	��_�43&�CE�!H3w"�	>�xt�0>��|@�`�����8���ޢ��&n�$!���
P����PT=�G�;T�65Iu0"�������A)����&����V��x�f�#�2�edlZ��\��҆�n9�2�T7Z�ѪIG�4�z�a����ߺY*2.y# d�X�[y��F�V�����/T�L� =h���g*���X"��z!��-�OM�67SL��>$3|��H'9ק�`(;TƖ[�Ν�xr91#�w9��� F��np����-CN�}@)�Y�"��K/ZJ��h�]�2 �ϐh�V>�f�� �4Im�,����i^\-��_�PތAd4��^�3���5C� R��^(͚R��L��R	uWѧ@ ��>�����lFk^�"����JD�}0�t�2�ɱ'*w;/zΎ��!(���޾���`\:M,�#MƬ�-y5�d�x��NH��pu�m�ڍ�Gt�HJ+]ks3�}���=�3���Ja��4L���+O��Ò�h�.��g
�����K�Q��H��,ZϾ��D���t7����q(�,4s������xI�͒W���Ԁ�'�4Yw[W9���#��b'#�&[���R[+��J��*Ԝ�9eZ+������3}�����c!AS��dg�������QcgD�2���<����l�Bef"����n�F	��g�T/FM�7�K]<��7=qu����1�������ֿl��C(B��M͖�K{�oLd���ߕ�院kZ)с�II��a�Ȗ1zNߕ_\	�{sq��N�a�:o�1}�p'�-l���B�!�hrI!ϡ�S��<�"s�b��T6�]%\D��ʦ@�{����A���K�-\#��cM�m�%��}񿶭e�X
�d��D�W�qY��O�[���:Yl�͘,��<�ֿH��椝'�T�k����"w��ז5�H_ ����R�W&��6��YAkR�eu{V��):�*2B($27QL�X)11��	��K?F�����*��Ե��Uz��ם\��~<��$�/�ٓ�,��b�'���Mi�>)W�T���������YƐ�^_��n��%���ԵA_C5*�lǹ��E��V�&�<(��ΜJ=��ޙ�����{���s��g���i�G�����8�`��|���/c�x��X~&&VTF� ^�@!(�9m����";�1�f�G�N�5��c�R��NZ�>Ɗ�p�Bw4�#���Q�Q��2د9� i%1Zb�|҈��X6��0uc<�vkM�ϵ��Y����� �<q�@߅k2��@�4���$:��Щ�f�s<Q8�>:�M���!W5�muD|�@]~=�1��r�4���Ė�n���_U�Z����WpW�w�Ug��,v�^*G�Z�k�)��\�f�ø=���) �R�+���p8���ͷ�u������iֿ���a>Z�z�ͷ]Uvhҵ��A�9�I�(�A�����U1&K�S��>;s�FxR䛨������L��$�m��\�>$La�=WS-�Ȅ���O��<`��h�$Į&]�@�쨟��|~�6I���b�c�����a��ο�s���d�y������||�o��ߙv(3��loa��u�%2��߮·G�/���v��])��T�� ��������_�$�ְ��1���3�7j�;��n`�vd��!�Cޱ�2�y&��� 3Q!�a0�IK,"<6�6�ǋ��Q����Pt�Ӭ`�3�%����WY���cJ��M�@4��@{��9��N�sCI+C�q�O{�p�����>���$d<�9��9�Zc'��oyxʁ�آ��q|f��ª�?�&jD�A�YR��,�O�4�LT"ڠJx�p�}:L5��zZ:�x����K�%Ēb�T�<b&{1�*+�B,8��|�Y�����	�.��ձO���QA�,xm�F_�>�v��id=��V�hI>�*��K�B@��\�<��`��x�$W�������}ݩ
��������`� z�y��A�W�cK��Fgʯ�V�8��>�k*�@M�w��l̖O ���{ȼ���� ���%�@��|�㖐������B|'��	�e@-?Ewp�>e���@����:��h������0
`����p@Zw%1rD� ǰG�/����H��H˔��-�~�[kv�@������>�d�D������M����7��>g��~5=�Z-9҆���v*B5G���^',fc�o�7�X�;[�ML�~H��A��)�^!�l���6��oG�w��>�D��a��B����pݏ"rxw �ѧ�o�~~<�q)�%Ƅ}iʐa6�����.��i�ǡ��n�v:aXx���|�A�f�����I��oYrY]̸�)a�����G�v0��e6yN���+"���ԅ�M�4��҆�‛X���P]9���ǫ'�۪+�(po���3@�kQ��՗T	h�4q1��#U��$���bT��5���M��;b�!v=�6:����@Oԗ��.���^���z��rwR=��o�O0"fQ<� ��x�\�xHm��7�U�A(���݋?��&^u����wSk�#�i06� #�kc�ޙ�~�V!}H9�3���.쏰E���ZC
9[5�ks�9���C��({�J�	�ʯ���A���_E� �oK�5%���̡u�fF���t�7������[�p
��0� ��)�+��Bk�AS�Ge=g�<i5��Hl<�l�}�h2*�G
C��R��Gh
G�vkf(�i�u:��O
Y�k�E���+��N�ئ��w�M��zX���R*�b4����/�+6*5x��)x�[wߓ��%=�k��K��v{��\'����x���}���mg��I�}�K]F��M�״��4wVIk����DbSs)
8n2��#)8ra��l�������u�6u�S(<��Y��J	�z��0�P2�W+�s�yGp_I���^��š\����[�>p��u�汭C�����xu��^wA�q#
�_ɤv5�gw~&
�4r��r�R��������&��`�-FK�n6�a��풲V�m�	Y'����Y�T����h∅���˅\ܣmJ\,#|m���f�#��4�N쀂���Fui��Q��`x�� Qa���+"�W��^���I�z�H��4�3����	���4m�%sƜز��u��j2)7��g=�q"9ŘC6�q͵���u^���$Ob ���^�}C'ab��+��b{^�!l�º��b.xZ�3.���4�4�b�����d��2Ӗ$aL'>�*h�u�H�D,�c$%��Z>�f,�nH���i�b�7�%@P@����&��l�>�^����J8��l�=�Iik5�H�������\�d�=���j'7�$.��Fʸi#cW��R�Q��D*�����C�s<��qUI֍>�"��c9�@�]�I���ZƘ?�9_ҲG��{%�[�e�����#�6|��:щ�bh�����V�?��~]`�������L9�C]Lz�\a�5�c�C���|�T�?��=&�⽩M 㹃E�m������$����b-�����o)�jDW��L�d��ưAK!^�ۿu�lb�3��v��=ZI���l�d���}�>�)�AS*\�и�\��ű�`L�T1��7�:��v�(�p"G~�
�	𬛹l�c���rz��.a�tOIoG��t�g��B�|�4˲���"� �{�l�<(`�w�Q���"���<1/�a���A�N����\��?�v"�K&0,�5?b�Х�Q������1�����"I����P�L��C�6�\$�a�]x�-Z�)���Ě>d��{�D�Uhk9���0��'�*�3�ʧ��2�ڪ��e�4�g��h�������5Fwk׋���`�D�����,X��eOT���������2��{!�L��ju
�^��]�-{	m����W};�;7d��o���7�	��j6˖R�['{.hc��{!�b�Ib�1�e)��Ǯ�����.n+D0�>v����%d�����F:�Ǽ��vf��zWů���93Z7�1�J)�ƙ'�(�-�-��^�*�%+�!H
To�s	m���x�`	�i���4"�:m�t�o}��\�hI˴,�mB<����{�:{��Q�J1Ov�߆��q�P�A� �fDӧ���oÖ׹��{ϝ27���/�j���˕1pf�=s�èE"����Kֈ�
_[���C��}2
P�t=n;qu��{�6�d�k��㇅ۓ��֛�%�mX��s�;��z���(���c|����?�<��������L�M��_"�~�[�q^��*~az	�V�ۜ���2��f��{D>����,$dC(4��d����>���o([wH��GW'�V��w�|����ɂ�R�
L�uMT|���[UV�,(����uB6Q�P#�&�)#U�'�h0�("��+C��(彮Q����h�P�SP��j�ޏ�*��d���-f�p"�T$fo�p}�KфC���W�B*B�W}�fv�j�b��w,_$	Kk��MpF1�2��#�@D�\��r��2�ȳ."�S�k��'!S�_�a� x,T(k ?�c�7,Ǳ#�Ϻh�M-�%��Y��o������G�_'cl�#�w/���R�]�˿3G�<�a�������/Eߝ��Y7��_��yؘ5u��`�Br;ܥD��p
�2+
x%h��_x��m�������B*��ڟ1,��+X�5���J����H	$������u�mA��7�D�kV����6?9��81�n-9����io�@�<q�U�$��a(Z�.�ӒT����~�g���b�3� 4�yz��s�_廨a���F�B��W̬%2.��w�t���
d�`/��ߟ�qj��9�y�̯�)9�l��/HeeQ�M���w��_S�m�ήNpđ��/��Τ�_��'�ہ�ҟ��^/���[�{�9Q��9��wW��.�|$<��E?@�u�/�u�.��p�h}!��E��G�S��v�A���fɡ�i8*(�̳|�N}�`ؤ�:�܊iuz�ƈ���Zm��SR\���E�,mC�>�ɗ�V���튲!�'ɏ�[�9A�s��dh��@n0�ZM��
\Vϸa�[,?�x���>��PI[��7S
�߫Se�oa���M��K3I��h�{�����v��E6X��^"�'�7�R�bw&Sa=�1S�}�oU�Y��ףqPM2���i�+�}�`}��4j���¿Z��J��zCu5u�������F�$,���=`ۻ�b?l��A�&"���<a�숅.U��$i ȉN�%L�%T$���^�]�{;]���,�o�8'��+�׵j5��(�,�k<wh9�ػ����)��>�*�}e\,�B����x��~��m�u�
H�����j7��A���篲G��w .�ݍp�O����o=�y���EZ?J��#ψsW�@�dh	��7C�rdk�ς�LK�T���a��c��l��(3�L���s�����$'a��hQT��a�XRUz�m�:������r���m%r�uX�[��X������=����z�Mc2qC��y����FTΉG�z�f�}�[q]�ȣ0�y���=j}U}�4TA��6�{Y���#��S����iW�=��x�l��ĩ�ʋ=�GS<gz�!�sc�p���y}u�{!%;��~���хQ�[��\�Ӳ���y��R)�N��i>�2h�?Y`��<���6��?���L������ց��n�%�#=s-r��\P#��S*~�s?%Q�2=���6��B�y!�K\��Љ!�	�?�������/��a��.�A4m�NZD�,���|�H^��&���@�&i5n3��dCؖ�2�,�u���O`���Q�tE�{Bn��{�����pv�lay@���W��F@Hb�3rK��/aK(
7m������������:.�U'б$s�y�;�Ez~ջ�*��%��4����ż�|�Hm�ӣ6��h�;ϡ˃ A`?�<$��.)�=��	~�j�p�m�Q�#��5���G"0��&e�9[���חd�j�P�w��`4B�ѺE��c0��ʍ��*���d�QȐ�%���:m3 C^�o���B�U���îfRg����w�_��.�w�vy�y$��?�
ϹN\�����ڦ�<��Lk��C%Jy����lR�X1B�'�c[Z�Q�5�c@��L��\p<���~<q��e6�LG�O�AO�ΰ0�`�b��H�#��M��Ӹ��E4K�\�
詪�zh	����[�L���������,5�:�%�+�R�_Q�gv��?�w�m���P�=)kr�ؘ�7�fa�N�uU>�.��O7�D��ZC�lT5�x�f� �nm7	���x��Q�>h�?g�!@v�bCַ��H̚��KgO���}�3�b� !WהU�o
������B'�'9mUe�����_d����j5
�Mf�'��9�������B�.}����Zo/�����Q1H�]�~	ZR��tG��M��|�}p5�9�(��:�zkX8}<��ihK����tk��:	�,��<���	����A�� �h����a�K�P߄R	ƗQ+�0m��% ������
Uol�M�� D9&8|ڨ�פ8�	���I�WÓeMY�%	H��W�������#+���)}�`l�7��P��p诚����gڛ��z�ݤ|t�9�n�Z�}Gh��jKÄ�X�)|��d�~��>���i3��P�N��O72�O�:F�	/7�	`g�C�+!���w5V�ĳ�]����jR�VAC�Tq�P-���CC��L0�$^���i6@Vz@���S�MSy�>��%p�(��;ԱK���/XBфW}"�V��:����NĀ�&aQ��jD��Efګ�5%�k5,�m+������kv��r���´;r a�z�J�V*
Oi	 n"`\נ#�{�����
��=;��״�����{��oR	�L�B�F��Ar;�"|���o#�E��n�c4�]s�&	ۄ�iwk�
"�*j�������E��A�Wxz�Y���\���O����+�A�%,;���؁sN�K�V�@-��|��'$��g�+���-~D��X�-����|��\_������b�dW1��&T�Z{�z��G�"�}
G|A0�E�tK��E�`�����7_qj����)��e���cI�:���NrHu��x���sD� ����(a�q��B�(�t��~���g�	�~YI��;�J��46�S�T��nBH�&��K�Hd�`w�V#Ү�<x�jaKW.���pقi��jK�d��.1�7���ćA:�4�7�:�W�-�^�^�$8�q��MU�b�� �}���H�d\�!$)�F^ƻ-S��SH�2��y����mH+�d����8!�aye��hYki��fX ��:������kUf�L`	��w{T1��RW����>���7#m_GN��^���TJ�u�L���}�����h?�QGj�Fk�wl20�U�Xw�Tg5�?#��d%�"H�b��f@~��Ao�B �w)��� �L�/H��-�h����X��t-KB���J�/��s�{��"�������7�Vӄ�ί���e��x��HO���k�$U�U��B惿���6�l�#dS��:0�J`���\%��Z�yr��]K-q�TaP�@��4Ys֗��<
}���7��1��x�K�(B��5b˩e�H�<;TNJ�ܚ�?i�h���x(ٿ 	�؃�Q�.`MG�_?�b$a��P���Jb�q�L��L~d(c*�eI�ٵy
����8�*�h"V��XXƟo0�����oI�f��S"�J[{Y|���A�0ѷ�c��Kj�?S��K�qĭ�&���^i�b�<jF;�!�۬�WW�^�m`7~��E^����G�?7��y���J|������+[����T�LR��rr�A@#��2��~ᵭ����08�bZ�����VL.��[r|b>��w�X�N��.�{[v��@���;�(;^y�)�~�h�#f�����k�{M#�I Ҕ���Q"���IU���oR;<hzWy����<�
�Z�!Ȗq�/�Ҭz��*%�Ε4h%k�&|����=(��r�(�q��l;?�h��E��yDh���ݦ�x�$u����Ť����$&z
�}�5�1۷�7I���*�K�feU�J���Oؤ�b"	2H�1���t���N;�^�	m<1��&��'��6�a!�i��8�T@(�<fL���+�f3bK���f�#�OP2�@!��V���CLN��1���v�@�v) T2�ew*𵔁u��Ki�g瘭R�!�S00K\�)xM-���:���{��/��0�l���tI�iAL��d���u��K)���:�L7e�D{�r#[��K���*�� `f+f%���Y��\W�\��!D��P���D�J's��;����T�Z,Z(���|l-3�0�����PMîo�o������c�U�d��w�< [.��沥�٘��q[CN2%���L�C(�u�����Qw��t�c�HYB$�o�"P��]2+;�=Խr.�����Z���4�_����B��G�NB��7�����mw����t"0iHb��at��<�P�[�@��)�fc�hr$(��AJ�h�"�������>�f<a΀hς��W/��ù�k�Ő��lU��q4\���o]������ =��A�Xs6br�6�Q������p|X
��������[h�w�Ԅ��ѣ��̪p��߮���P�<����'�������p,p�m�ߠ֛�cR�q+V�rr�����؆�&��rQ�(Z��ʅ���y^W�p��
����������X}h8���Ԏn`Q�#�������Qn)��Y��H?��c`�ɢ2f|�x#J{�h<}�v簑�0��՟��{{�E{QkC�ޕUah�&�׈t���n�pk�^
fp!l��V�j�GJ�`�6�����6�4X��|^�����o��� ���;�m�9K�\�4������(7rN��ĞD̰ϗ!!!���'��:��=�չ��ѳ�Ǚ���[�HBs��r_����P3��� ����ֆ��mM̚�Wύ6@.�[��ל��K]	2�8?=�K�y��2�f�z��h���g`7��q�,+�7���Gs�v]�ݱv�����?b�sڋ/����(Ǫi6�G���7��O>���eZ�@�V�)�OS��HLƃf�s������~�hA<��dS�D��w���˱��~�<|�~r��"Ƕ���4�՟��c%��ˑ���(
�q��ֱS�(�w��Ӿ̵'��KaW��h(/�v��y�J�?'b6%��.Fι㶴���J��OhZDk��'�����PJ�(�zb<���^ڵ/��f�m�?���lSS�^rpj�sD�{��?��<P7����֔�6#��T�����=HX~��j��b3�4���e�c�؇1ｮ0�`���uU]��?#/��ʥ�_���vl�w1��Y|��������x�Q��|�w����Ra�'����gOGR��\��X���܂RF�9t�zN�����v�ء�]�#���J��o�
�3�G!}�X\>␥(:�^�X�2�y�)+�p� �)o[�.���RAAj+�a��7�R�-%*$��\r4/�V��D��=Q�,_	�����*x����n�m��R:�Xp�H{�؎��J$8I���gk�h��?�l��A��A�g��2�]l��e�<�[�l�O\q��G�k|���+?��e�����?Op�-c��΢Ͻ����x�
��=�
�}���.���㎴������$�EE!�'�۩����
��q���)z#�fD�']��2�&���OV�2��;����:������ 9��L$g�B^R���ըV��m��+l�SHJě1H��\Fuo�x�����
ѽp��Ҭ@�H���K�uM��gb���`Ƀ�p@��u·Q���Qa�L�j��I��d����D���!�-A~wk��ܬ)�_N`L(6���/��<���r\0�WA�����V��qP���R<X�&y-h�X]*p�w��=�ۖ�Ki@�)ı��.�;�J~%��c�ѕ�X�#kh`F��g��4s$�u�����c����l����g�x,eŻ�M�N������� |�G�RC��%��w���}�5b%-��!kB�Ks%����n�9��R����ЀӿC���k|ڌ��8壐�,����8�pū�3��!mY���A�����	j]��=��x�m�����?���l�ϟ^_K�j�vc�������W�5`=����G�}�4a�FS����p�"�!]��~Ix|�C�[�����L!�o?n�zVҒXt��}G���Y;�䳵ZTh�(�{u�C*a�+v�<�qh�D�]V$zԽGy��)2�`�� ��D�S<p0���2.�c6�ˣ�ھ~v��uL�Z��h�ۀ�\�T��}��z���ց1u�8�F��>�n�r�j^9+�N�sW���z�Q��O�S�m��[�v��#��>��
��|�)�il=U����X��x�u!�`�F��b���#DW��3��ܿg���P��HE$=Z4��`�������T��G0����6��e�^��rp��������W�	��c�������E8Uэ9�o�32�RIp���Y��$���]�w��n�������2&Q�#���KN7��|]�^Z�1���i���r�����h�F��M�,��� �歅[:v?��_Gf	*����9L��pa��k��S�k�	��P:*���Ǭ���C(�k�x�ʢTKQ)6����Y�l��g.����d�tl�ˑЅX��T�3V���Nj0��隁���d�8G,%<��E� �b[i��C{�vg���psZ�8U3A�*���Q��[��4_�Y���k~e#L�)���8��p�T;�zOC#�?R [zc`Y�q		��f�5T�P��XOy;�c�+��9�ݝ~K��`��J[�bƃ�1�*C��#��`�$��v���:Σ�*g*'лyc�A��4*\B�+��w����k�)pJ�'�� Y܋Ә��T�=ס1'����{d��T쇾ߗ��&���C����gHy%��H�7�cd!ɧ���wi����?�%�T�������V��}m|Қ������o�=��)�;��Ź��/��@�f�ݖ*V�wރ��4�h�����(QlbZ���n��X�E�+���* t����<�#"�wO�S�#�.{VKt\�-|}�)��#L�svwɀ���P�u�(�cE���N�E�DMT[m@@��#�1+��G�j��XH�����C�i�)�C�|�?�JIr_� ![p�F��T�`��:U*q�����7��>�����	��U��:Z�g��	�v�w��q�g��	����W����I|�]��+�ޘ�{�2��
���ȸ"�[
��d�*��0���; ge�/ i�ݚ�>��MS�� ������M�o��7�mh�~�[`a9�.t����'�������
�Xl�N�����{04X+PO��4�6?����D]zN$�3e��A��հ���w���ɾ�������5r!�|��R��JL�ď�g�U��[�T��,�^u��s#���sL��h���2�:Z��E����p��.�j"��ٴ�G�3S
��*u/�i�C��Bq! S{}�Ԟ��z�������&� J�N0�.	п9:�JӘ.@(v�(�����ol�XQ5&��!`?N�~\й2�5�X�wn��#���CF�N��}�E$^�!��3��v���T���ö�����l&��{V,���Nx[�z�a���*�<��飡*���d����Q�8*Z>�����z�DA#��iv�F�O�J�t�%�����C�7+�-2���y�!e��{�ANdRV+�-�q�M*�C�@R��:�*�BI�_sa��Nd/�iPwp�T��/Yѝ{�iO�0����0��M�c�Z:�N �C�t��1+�eN&������H�@1�cFgr$F���R��r>00b�1�b���=����,Yf�"y�����꣦'əayS��Ҫ����⢉�Tl���/�"�N�2^4ڰ��8E\�]��$k)r>���޲	�2����4��
����z��D��2�/�A_�*��]^!��0���G��"4�N��R���{���U�)O��g@�{��	�e|A�T��
X^p�턁�_�_�9��϶3�E�$ �s�-ʑ�C�z�lJ�t��\$��5�y����rҦtq�h��gs�����9�m��TM�=��3��S �L�[�.(vӨ������,�O�WY�5�+�gmt�3y/>��&魭d�6wzr�a^a3T�Ayy�g"�u����5Z�^-�|/�h��5���!��✴�)�O8Dh��4"��^�=�H��g �J(�((7��b��nt(6%SC�Hݽ�hQ�x0L�4�E�z�e�_Z8��f*�Ʀ,�Cna9T�<X%��R��S�J�$�HY�?�}wU6XcϿ��Wj�φ����:dս�[��<��ࡋ3���^a��H���[��>��Jaf�(Q'cz�ʥ�]|�Np޻i��-g�N2YqV$�ɝ\���:��>11x�m�^O܌�"xbx)� ����m"������C#��̰ l�mξGbS��C֡m�=�^��؛n��j�%F����߶	ֶZ�M��Σ�0�MO�e��,zQC`x�g�10���`�C�����IL�ȱN�SK��!v�br�*w��c�f*\���fp�e�3�MŒ�#g{+^���$���y��� {�3�Kpn#�w�v
B�&�?�`�چ�( �:+~��o�i��PP�D֣HTȓ2�d���T���� ���\����?`�3]�]�4_j!��:b�3#F��N\=++g���G{�a��\�8C��NɄ�jV5*��Tnj�cO�hJ����,��$)aK|{Xӥ㳓���%�~B���v;k[�ӯ�WT�ᳪ��%���nW������ʩ6(���@Rz�l黧x�6W��"�͂�bo�7��{��x^@�T�!0�*�8駢�bn<<RZ�Q��WV�X�O��\��4�Mn������t��ݠ�e(����&l�vn�#��m�E^�B���q��凉�»X�Eu��p��@��Tt�o����u8o����o3(��u�>�a�Pџ$2��+�'�'�����R�l�]�� x~^'��g���&��|���f>��	�` 2e�`��iF?�{���~��e��2��S|��ͱt�R ��Y���Kw#�� �ʛ�9\Q��.���$Է�X��G��?w���ޑ��9uDi�c������!���6�9#�5�q>Xi��e_\��_+�$�~�>�mn<9sWT�Rj�q��r���ky�K{^M�j�(X�p&H�܌a.�A6�� �B ?�=���_S�4�a�J�J���j�ЦQ+*M��_����d��̈́�;I���f��0�DCbN"��L��h�����rPf��I \c� �I*
�:�d�u�^1���r'ѻ���]:��b ���:g	Y�Z�-,MO�:�5��/��:��!o~ĺ!.���g8�nԛ���R�9�|.+�$}�hU�|^���|K�;������9�i��|n�?���%���%�N�.��8�m�wt2jr<g$5\�f
���t�3A9�ª�o�/���Ye���e���qdm��,�$�Ξ=N �ޯp^�M�3�GXv)�!2<Cż����on�"S�'$�!�+eV)NN��y)w?�Y�-;W��������JSfs�,�i���l�i;DɶDu��l�״~<���+'����Ycٙ�U����'���z�GY�03�t���,���O��g���)�~W��8t��[�t��7�'h�k8R�z����av>sf)%��/�Mh�����i��}�|���zt���2$Ir��\6m'�'`�V��C����1�B7��,���`j��8� wâGnud��p��?���P�*�x�5dv���s>�r��$D�Q��dɎꅁ�]��u͖�
�~�ڱ�*p�B���:�H'̼`�?�%.��H'4P�XH�wߌ�����X���4-��"jc9x�"���_�pZ�?h��Ӄ#4�i�@D�	�{������(�	���?X#ʣ�[
+�����Z�����	~�|GϠ��ޓ�NQ���D�9�&��QHw��pQ^�O��hd�\'
���;�P�ޣ�3|��q�AE����q��������Q����M���݁�PXϵ�#P+l�N������r�RM��ͳ�Ԭ�wKB�x@Ͼ\2R�� ,�o�||���oŮ�sԝ�e�����yЬW�.�(�ʽ����M�`f��Xz�����`�����h��?o�((YB���\�$_ZC�|�֪HքX�t��# ���>�!�o�yru���;��
�S��b���[��x���ӄ,��"�)lKC+@A�/%"fyJ�vDj�����u�w�YVzh�`,�	L�Q�^,g���LϠ)�-*�]\F���ڲK�s��oՔϙj8��j��L��1�N_f�	e�%7� �s�Lp�	�`�V��t�`����z��8�y���>�М�oeM������G�x�> �����O%�5�ͳ���s��?#nHςxR_l�o�hUA�.:+���I=D�zvي�ٓi�(R���֊��j����hǡ�vnP��\���)%1'�~'2a��LB��.��smb�,TI����z󱩍������u���Ωa�x�F�L�y��5��d��.�ʵ��y��dՌ�<Kg88⛌�J���E
�H/0��ſƻ�C�,�	�\溸�ƻ.�?�;�<�"�Іۖ��|��Cf^�װ]���vm�"��$`�d�m@����S��eM^����B�nM�A'�;� ��}}�Oѭ��
��:��]�G]m&��c��L�!A�\���5�91�_��`�Փ���*�*,�X�3����Z�}��A%6��`��b��Ob�Iu}��B��o�K� ZV���u-��n��8u�.���Ip�L�O���F�{X֗m���xn����J��*#~Y�wP[Ӵ����хƎ\�����J�3h6-����������Z���R�$@k�ZW:�r2඲�����"�h�i���Ϥl>�ڭƼ��
���J��-�pRDn[��=�����U�J]� BO�͂$�����[����R���'�V�` q`T��ۛN�/&��`�#Y	-�fS�"�� c���(���\O�U�wr�Uڻ
T1Y*z�<B�R�\��k�:0(�*DF�H�����:�<��(5��[�qw���o)�4��u�C$��V�lݒ�O��p��5��X��o�U6�ea���(:G�M������m̴�
yt
M@�5%�>k�iA���]��ɿ���ڣ����c%�Q��ˀd�!H��]��g��t�BJ"��o[U�����'���/C\۲m�2X�r>�C�XvF��g7)'aک)���~�2;�N�ov	z!x�����m�A�� `��-�����(��Q�Y�:��ԱU��������T48U���f���j(K���V�O.#z˃�����/���U������Ƞ�v_���͆Y�����?��?���ۢ.5�A����Y�O;�?s��x)��֨��Se����v&Xr�{�m�JX��Ih)q�]b�pL�����E�]�$�{�>8 ?��
�?`���/J�i�D��H8lj�;of��w��<]�[��)ls�=�^�i�;/�E�7���.�[Ve�;����6_����$�]�D�t�(SAy��i���gqlrV��`�x�b��݁q7��#���J�1o�+�3ĳ�: 3aQ�"`o-��z���ߺ_�;����1���9�'E���h��b<���l�;����V���r*nPˁ�z���G���xv%V�*��6��vm�	Mh���)�EN-���z;NW�����3`CZ]xu��5�g�R�1���J��R7�1� uoRs����| ��m|��m۸�aw���^]ð��!�_�=*���v��Z~c�)����:�mĕ�!�x�����.�޽�/�?���/\3{o����\ꐻ���E$8���{$�����kYܱޖI�t��� P��4���2��:>QU�Ć�E�w���W��l%7	��Uc�Q���wLaTfPD<�������ku���-ФGn椾����ʮ�׵��0,K��$��{�²<��H�A�,�;w�IL몢F4��::w���M�2[)R�\	|&�B��]�I��Lt� ]��� ���5��4c��S�@(�®43�w�X�|��[���I5t�F���5Dp(`�=~Tf���.�!��<��[�`i��-�5�"��{�a(�c�`#��L�6Z�#^��*�3�ح��I�6ԕ� S#�Y�<��Rv��F�����{�6��{�z�QI����aa`�c�_#��'�A��#�p�۴��m�2�:�3{+/��0d�t0��9����E���d'/��p�[)w
������c�PrV�ʛ�q�R�gV����P}`���!�����}%������,<]k���{��v�¸��*ZE|8gk*��<�Wj��Uڐs�+-���5���l�p����Y�J��@��yt�7�B�7�A��Bh�ˮ
ػk�Gp��Щw.�z霊���(Y��"�#FH�E�6���$[�����'�Q�����h>�U���۹n�B�[)�E�6�+(�
���5X��0O��HNH�&��#B"��v�I��I�W�Amע:��.igh2(P��{}��^���08d��O_>�辪rخ��z���!�e'5 �	;�d9�����Ē�QY*�N��$��O�߹?�O#�8��C�c�\RΫ��.�	�9z���n~�E�ҋ��`HԱ?v
��"���ns �ɉ�@�ק������l�}���k߿FK7C��Ӗ(�˪P���!3��l��9���:ǌ�a�DMwZ��0�L+2�sT��U#�k�h9���� �:�Y�cN�vk����z"O����R�Rn|I}Jw�o�	���n�k���۠�a�2�ߐ��4@_���̎�?�6��`��dr	M��P��&�>�(�Z��	^�Eɴ~�ɷp1�^��НR��� �&�G��s���	acE��|�%l[.�f�H)Q>�������Lm� �23�ɡP�o��^��
*)� �sb^=�%�z��2|�.�uu{6�m�����C:����!Q+ܥ�t&����n�ZGlӃ�N�;��9U���2���3QG{�OK�����s�cAB'�Ik|��~�{��{�b�%�"��2e��P����XA��⾝�r�ڑ��4r��y�/^�3!tn�H\xn�Vnb�s�,ra�(h��կT�sgg�u����b`��Z�>�͟���b?˵�9���'^A��mXS�G�mTE��oS�~���=G��3v꺆в�ˑ��n*Io*+��5e4�CYt�T���!��>cGd���~Z5�"�_�����*��*�6b��;�{���d���L%ec�Z��/m�Y_�u�/*q��|k[�$wM�7���n=K$�|�@������E��v��J����G�/�/
^]���b���#s	لIq��*4�_�"@�w��l��\UF'�ɞ��6�)<�����,�/�ЇV1~)Ç�«d3c�1=@f!�@��ғTF�?���E�+˘���8 ���)֮w� �E�[�(�(��H����z'd3��!.T��=FY&˼ه�WB�*~�ўiµ��� %�*F��H�ԝ�C	�ʔ����C��_����x�mW�R�/^��x�p����;�3�Q��7�D�yD���,?���όb2	�	���fm���+<O�d�)�iJQ�G�q�"ѫ����e<�J#ۤ�Hɸ7(Ԟ�d
b��6�Iy 묭=u���GP�*Բ�I��Ŭ��ڽ��%*d��ѓd�b^�,����>w��}�cyڭ�{G�����! t�`CȊ�F�C����':,���|��=�k�xå^�P��� =Ğ��ˢ��Ny[Yh!%Ԧ2�.|��k}��U3��!��S�īZ�SP�Zv@b��{&�'=�n7,�v���;��L����^�}�Z�ED�Z	�ý*,�c����D �$psgӼ�%˶�ɺ�n�8҈��fQ��襤؜��	�%(A/]vP;��p>E�>��R���������F�*nc=��u���ޏ#>����"�t�!ƞ>��b?:
�\���@��c0<@�^�t4.N�b����_@Z�a�k0��!{'"�b�Hj��6쉝`�ӰN�/��9�Mt�[��ً���0�Ǫ��cԻR��	�5��[�M�8}C2�Qc����j��N��K�ȥN� ��m��S�@���f��پ>��yC�����9�u�C���d��3=��_�:PM��w�s�*�1@�Z�| �Su��3r�'��٩ewݤ�ٙ�Q#V���?��J���)�!#��=�)�<��|3��k�4	GQ�)1�u�(Ȫr�-Xx�謧/VUZ�����M1�4�DA�`Av�+�b^���sL#�<>��0!���y��	^��kȡ$z����c��)~������,?�7�,��ƃ]#�ӤV��)7��Lk/Y�MeO��]]ı)��;�،�g!̧��;�*��`��VS�d��ʗɎ��C��׀�l�����Pc҅!�Z�x[9�����7���jg؃~�e�zn���V!�z�J����R6t��l�̐����aO�	��ď[h�v�&ڵ4�@L��ڃ�A�6�XT��qB�5}Ǆc���>K�B��d���І~�~[0N!�X���%z��Y��A
��祇�\G��bk��| ���f�z���7��E� U�+}��y}�@ߟ>?���4�I�g;&����dJ�v8�}Ԭ���ѵ�\��R	�����R�����~(o.���Y/�M����*� kԴ�@�S���\h7�ޒ����:V�-wIkј���z��F�����3oe��e���	�L�zQ0BC�P�����8qՃ8�\��M 	��NE_#*g�?�-�A���s�n��J�ﭏW`iO�_��ZD��zTo٫��z1s��"RS!i$���#{�
H�l�s�6���V�(jNI����M�s��yM��P���`�u�CZ�5�VѼ}�HX�g��E����~�o���(����>^�d�����o�8x��.{���"x��ԩ�WnXa܎���0(n�n�5)`�r<��M��E�Hi1S�jZ�g��:��л�ϥQ�Ӌ��,�[�A=;b2�;�\��<[L���%���qer��pȭ�RJ&�N��Y6�����\��C�F��Ul��Tu!᫷�`�'��_�6cI0ǉ:#�!�����M沌�>E�A?��P��я־�����@������2��j:r����sGi�<X_A՞Vu��|�ab�Ζ�\0�O}�7#����.�'��Z�Ʒ�Ͻ4RK�/)&3�v���t�X!�ͥ1X�k������'q��x���E���:/�OC���m4�vԎEV�IhQ�	509/^���C���Z����qO�ø����0Q�1!X����D���I�b��gRV,z��]eoRCb�z^�@N�'��&r�����	�W��Г	��]����w�K��>]�q�VB�.�|�Z��h4ZsӲ�ǯ�#�ȠD�}1���q��j���]�nuPhB�L���fW���|���q55;��B7�K��g0'�[s��yZB��Ӿ�n�3���r�-r�sV䎆s@cS@9<��n���{
�ƹgɫ�R��/����!��hv&U.Q��0��Y4/V.U!Z���RG��
\����Yw�4��C����ځ� ������ O�T@�!\l��%�ye?�{6_��� mD��Qp��$��=y�����W����v �3�k���1� �]�Fߡ�nX��6@au'/�9���J�[��m��f��W�r�s��m�G&_jAsp�Gg� gS1���7V1�j�&��
�n��͌t�t�i���F��� 5	q�"0(3�� �HN����:���ʅ�Uq�Nt"���n�'�7����	ĵ�'w��708�U+s��~��e·x��� ��Nx�U��y{m71�>��O/떉`�!2dR�$X��P.��޷zt�N���t=��70��ʔ3�K����Vͺ�[��P ���U�@�m1�.��4�R����"s�[<�]T)��O��}��z?V:e�6���:�,��R�od���:��i�r���b�"IJF�K�a:����f~���E�)!��YʿƮ��'���Ű���I�G�(�{��d\�P
�b��UD}��2�͹�w��]'r	h��FSL�@�}�)��\VhN
�w��5���P����s�+��:�U� u%��KK�A��a�+Ɏc�ȧ~��V�j�eN�_���Ѵ@k*ʢ9��]/���B��D��B˦\�A����Ѩ��#e�8�Κ��=`�~7*T6c�2�zx+~�9�o}$�f]4[�ؒ�ݶ3����X��LK�68���i�9�4�ε�Ú�w�.]�	��R%��Ra�:+��oxE���V
s!a�?�%����n���/q�#tЀԛx(�����_��
���#5[�ȌjPORNU�+��A��Į1-�)NzJ�M^�E���@+�2U���{�!�z\�>7��/�%�%�1�;���ċG�#�Z��.�.���#�N	g����� �����5�R��Ɡ2�)ڥ1�=�'Ţw�����;g�-Q�*�B��\X�60#�5�&�o�%D ^-�w��0|�qY;���W�����>�`P�����	
�kl�֌�:�*��%����ƩSf$�39�_�~�5Y?��}p��'$�h-#��?�Wx7�x����Ǻ#�9�Ȓ�%4����_0/���ӑ�A���{��|p�@Sk�EU���B;��_�z�nm�N��~�RLld��d�d_v�G(]"���o�I��8Nꗬ�R�8Yr�9�U��Y����T>dz0~{C^�C���7�2|'���j��6Ё�oϲ\4N��a��2���_��9uT�{�F0	b�Q)m�4��i���M��M�<��t�B���o'���gW�㧍q��+0N0�3� o-h~��r�`�B���>��
ń)!��p�rk�yK��� �/"}ۄ�J��&�����;**�5���F�?7]k�˓��L����-��Źv�s�]'�VN��r
�DiG�����Ee5��;��h��,1[x�mje���މ��*#K2����+0f:M���]YNp��l�hOh��>B��$Z;��X���ϖ�-��Y&��q��Ĕ��P*W�4�MI �n��")j�K��XՇI4��[��6ۮ�D�%���9�J`��ߴ�#OX)#�:[��v;V�C!cQe>�1%�W��=ۍ"�^`�30�}��gП���[�w���� �ʯ�� e�����-E
�-��$k.��������1i�4�ɺHZ��Z����]�ޛSO��	���r�漸�uQW4��M�lQ��A�����X�SW��~�`��Ӗ>���gQ�?rL�+���ARk
(�x00���Rz8N��3��:N��Qbl@�P`*�":ַ뙶G�!$�Y<ǹU����GR0ߴQ�U+��|����V��*[�ƮB,�4"�`�2��D����A@�	�a��r�1��+r3���|�������Òuz�K����B`� �OZ�}X2�*��pڌh d�����b`	�GL���נ����\hq��woɊ�6q�T:{ 82�W.���8�)����H��ӍǴB��x��gC�]�7oB�J���MO[�|�)���q�S�
]K�Mg
�Zi(	��?�}��.�⩑K�<:#^u��&��'H,��P�I��*Vu�	��÷����G�k��y+[��F���c�"f�x1J/�d\�'�q	�YUr�	xf�U�Jw������W�����<#����p��o���k]���)Jo�R�bW*�2�X��HC>�,Q�;�p�f�JQ�<	7�9,ZN���wm�&a|n>��S�m�	;⅌<_��*���_ƭ�c�|S?pF�g���I�Gi�� 7��l4����V���c�A-��J���IG�2ɺ�/!E�t�GY^ ��mZ�����W�2&x�r�L����tZ;=�/	��n�*2E��LI�\=i'lܖ��d��a�n���K�<��M]�u�~��>��zn��H�����s����R����<�b����]�������~ʏ�̥p����)��0-�W�f�5�?}�0�'��f�z��d�J'�%�>h�"U����Z(��2`��a�{�������X����7�C�L̥�Z�DնMv$�R��Ҋ��?��l�R�6�M@n��S\��k%�+:  ń��p=�Q�9q�9ᨿR6�b��|o6q2�3�+�G3���S �J�W����Z7X 4�
�u�͙���gQ�2+�8���6�
�������--i�0�'��5�	c�0*�W�4X*'��Ik�o�
����W@쐉5��8?�ԥA�I٭J���#(�
$c~v�1�3��=m�b$��y{�����~��۽�iɶ�+��a?Dh~(}Ue��={�\}�$��`�O6t;.@�XU9�-V��D��CA#�)C.��\��1c�J,ɬ���ΰX��mR�ݝj|đI�����i��؉���(`¶�m� �Zu�_�3�>(�+Oz>���<^+-��ؽ�Ě?��=�i������#ǟzp� ��E�uA�s'�tY����V�:`q9ϖ�]���ϖ��Pa�~��Y�~%6[��<ݘ�s>���!3�l�9��{�B�#A�%M���%��~H.�u]�pl��o���V���z���i��~�l�f��H����K��U�����8 Ϥ D��O�~-[�C��!�ye�G� Tò�23  G"���?� ��5ޯQ��?�)W�e]�<W�t�.�%�=ՎO���L�R1'�L����8�����t"�>~��( �4�k��2c�	�X� �?���5�X�^��W���.�	�&���5�����+�h䓲�N�B/v ^,��68L�a-H�&��@�ÉR[0*������9a��E�ffz��ݰ��*��b��7N�I�x��ǴS}t&G�&"�xzٯwz�x��׎�� ��`d�O�5�k��j���F�)͌��ه禣zd��~��Q���1�7FD�y�ʶ�AU-Ĳ/K��ڻѿa���0 _i�T�/A��#ͅ�*�+]��ӚN�4��OڝF�Ѿ����6POL,�8.�4��sd�/c_�9�����=����E2�w,+���Ӈ�k���6�?B��&)��%i���S�ٵ]`a�P&r��[.F��mU�s�$��y�F#�\����E>,��ˎ����k,�L�k�^)�����܉�鉱ٱO"7�����YU�Qh�#������ɯ'�����l�z�	B�B#��0Ǣ�<"�Id�W7a���PƓe�T���|��!���C����~/�XHL$�2�ϸP�"y	��C<'�b���D���K4eE�m7:�Ɯ۰x���ˆ�;D\�Ie��wK�g�so���c`�,��5�!�9��*y���]��L�o��Ԛ�0&*��hE�)\��D�*!O�ݣ����V?�V
J)-Y�`�5�(.�LJW�B�Ҫ�@�Uz��7�+�}}�^��^ԛ��"M��eJ� 2���Kt��(���֪m`�s;ğ�վ�vkH��
�
B4-�m��H����3&`Ղ ��J����?/.V��������iK,7�C�`(�#j��\��YB�51D�e�NA��:\4`FO��W���g1���\�ا�� >*]E1��ɱ�@��DM�F>��ꗤ��e:�O+���b,{g�(u�ϰ����v;eCI���e8:o';���%?�w�}t��ȯP�fe#��0��'�[�=���~��wGF���{~6�*Ā�rV#n�3������s��:-��h�&p�}�=9�. g��z����̔X^\�����[���'���=�\����)��h�՟ˌB��X��L�M���1\�&������4F[\*p��4����x .���P���7�cd$?�v�u�+e<�D%�2x3�~�W�h�:l9T�����X�:�]���Y���H)-j?io0�� �����r҄�,�� ���*
ҩ=M��T긬fL�v�i�ԗ�D��9R ��S��/�`鱬�����?'�_��9]�'ޭМe+}��ߐ��3G�Ͼ����׵��7T�����^�]MX�+[/M:DC��JہTH�U1]?'g�a��i�ēZu��J(�Oi���)X!�
����m�;��%�-����֥k�&J~�A���q�Д�Ȥ6��uuƚA�Uf��`q�����pȓޮ���Fy�}�\�k��%o�������c�J@����h�-�;빛�a�P(�%/aѺ}.`�O%��(�oC�4̉e���p�H;�U�(T]h4���
�OW��Jȕ	q]���Uy���cλH���F�l�HE���Ȑ�,
�d���^s��S�5wCN��h�u>��E�r
Wc�>ƶ4��>��:�is�\�K��̢�\�F�wf'�ѕI�guzx_�(�q����9A+�7+��/O�"E_���}���:����)<�-�;d���v�Olst�M"�<j>��D��4><HH���3�ʥ�h��U�f��V�)�2[��a������M�7]ϦX�
<�*�֛v"\bQ�I=��ďBY�l6ϲ-�}�����n(�b�iH��f��=*'u
�"p�����:?�]��AF�}K����꨼�{����+�l�i&_D���r(�����xB����kL���.x	3��Dj�������E�c��T�m���᨞
��%���2�5�!�4�F��*�O�~E̮�.Ƣc����xV}�@k�<<A�ؠjjVOK�G�O�; �Dl�8��LS�i���3.��&�?�o�ȫc�����EIvV��Ȃ�nQ�l�n���%��^`ӕT,%IY���ي ����jm��/�����3��5���1�w;�Jb��Zf��*c�J�1�H�7�*=�S�� �H��-�S���M:Ƕ�c�~�)�2?��ky9Ųd���29^��L��r�NGξ�$+�,�����jm,P�*�7��e"*d["�/u��p�����_2"��a����C�}�
1$���pf�}�^ì3�v�A4���g�?�'�ξ��Jl�0ꊟY��@Qk��Ѝ~(U*-��������eL�\� �!�Q�m��
q��qkf�� Y�60���V�Jjt�=�A��1�9�n�|"�L���B5��+1�Dًo�V8o�<� ֿg���!���2>���!��?��#!M�)���<��˙���H��<���9��*[o�5~e�t����>�Z�~��6�cf��6^=�52����	t�Ġ���:�s�>��6VV<�A�|�܌�n���E݃��ܴ�|}=w���Q���~�J>�~�6�F��p�X�
�%����ϝt�u�O��D�H�18*�����9�&?"Rf^}$Qs�=cPyn���5�3���G��Z��;d��pY)�eW#G��"A-�-w�N�Τc&�����)��tHJ�s�ع�v��5=��!k�	(�k�9 V�Se���w�k���x�{�:���n���O�Ϭ�/����`���-R�<dxf2�r˸^LӺl��.��7�������ct�LUо���C[��x�'s���]�G	Z
W���b�2v�x��9R]����eQ��+�5<�x�M�;��T^c'��x��%��3�H΍���Tm�(~$��lZ�n���.������o��S]	�y+��j��P�3p5ŭ$���RXF+��� ��oyєR��ۮKZ{��XA�<6��@e�@g���X�u��i��ƈ�Z�jM�^@�F�O��s��]W�S
>�0���k�i���[-���k}T�Y��ߘ�	�%��7��d�+FL�"���@]mo3R|���;��7����*�h�-���an���1���5d�\�Zj� ��!�=��XB݆���J�_"I����I�h�2��]�o��nC�U8�4�������XI1���IX:��B]L)X����[N�㩨)�*p��SG��ϻE0�nC���GnN�̒m����&��-`��}u�"<.�;��X������T�h��s�yU�I8p	�!|����{��D�P��?c�G�by/���(y��*n�b�}�m 4ѫ11��$GO?�x�4a�b$G�K_{�<?��f�L`���9���u>`����GdBC�)W�e9/����Ӥ�ժz{���h������ݪ�"�WX�v�?�x��\~�4�ϟ�UVe�Lj�)���nʱ�b^h�?����j����^�~L�����fe��"ZB� c��I���#�<��á�B�8Y��I�����\�`|ֺ��� Q:��[�	�x��w���T�B����8AƇ��r��Z���{l��\4te^��	V�󯭀�4���:q��.��t~!��7�#z�1�_ZPv�F$��嬛�睄�!<E��JSD�8��<�Bm�m��q���l��K�=�-�M�=lC��P#@��P� l~�Uk[�D��$^��bU��V��#�o2��\%v�̀�iQ��&��*GV�O��L�QLN�g"h
a����W��G�8HJW��'r�e/�6K��zK$�2gu�T�П�|Z�Ӽd���
�y��ɜ.� �&ԹC���}e�Co�]�F�w�m8�q"�̩�#Z���@��|�+���CIZ��gH���3�
^���%�Ob�3�v��,��0��U&]�9�ڜt��
����0�����ף�܁�����yn�l����`�9�_|�)UZ%�UՈ�<����=D3T�&���RtDN_5�=ϰM�.�ϖE7Y�h� 2KЊ���c>�c���{Qp�U��G������_k��͙b��,|;��d��BmSVC��D(�d��`E��s�ö���J��:	�Ga��Z��U[�7�&����R`5�����_�3i��R�MΙٸ�>��b�D�*� ����Z2_F{	��C������A�L�4ϔ48�p�a�<
!m�7q��U��{*l.�q��	����1�"�6.jѐG���4�+��7��}pf�^k�$?�`z-D��WDth�[�j���'�����ޱ��i�p����C�/iEAlï�~w' ��@�seAk�Ro��=��Ҟ��?e1���vrP�ɽ𴷐�
9YFF��3ʔ���~pn��[^�G �iV�P 2AFT�v����}�=�D���|)��x���s��`�wf����%6ݵgu�Gv���
b�դ�ā�X;rP�_��r�4��U���o�rf�l��O���:+�+��JEyvc��c����,��. \8��&��1J5�Xo7��"y��>J��]X[|�LrWR��y����
TO��,�����.e�a\�˭>��4���z��Ο�.��Ե���Օ�> �V��.+�Gj�b��Ax���,W��F$�44(�9�K�	���j���<ے1��-D�B�ӵ�T�@�T��үو'\� Z3݀�*<��X��~;m'm���),0���pɟ}�㌕��M{tT����UD<����*��s#�g�GT!�糘�icOjK�6�lx���4ե����||��0�j���P[�4��U�Z�1}kG����'O���<���0���&3�����
����& �{�"����h�i	�`L�|���J<GK��0x^�(�u���&��A�ABuʚ���h&�=:��(;X���ڴ�sW���%ܷ�#�P�N6OA�{�+`5�������&�Y$��3����̋Ab�hGϭCa�i�2B���%��L�OЯ���Ǎ��*�=�SC���s-�ʕ����wv8��$OQ4�n��P|�3@R*)��x7N*��#_�ӳ�7V\:����y����N�WON�gR�^;�T�6_��D�ĩ߄���z GL&�,0��s{?��g�a�7K��L:�~�K�f�z*0�˱�Ӿ�}/17���=�a�KY�F�ۓ�|�����as%�w�`��zk7%k{\8H������-�I�!���&��WO��5���G|-� �N�J��ia8xlT�IY��_��r��0��mo3�k����$$��yf
	0�)����U���x�����Wc�+�HK���#NW��c��u���ۼ�XV���U_����(�=���`�;�7i��&a6n|�׊J)z��l�������/��n?����j�$����&4�cH�j.��=��m�!\�� X�6�Ti�y>2��~���UC��!�=�Q!x�g���q]��M�em.�\F����g-�%��$���B�-�y����?����P�%#�']�*��$WK��K�s�A��+SQD�������g`�)��YFA= B�IG�l�K��VHڝ%��,�bO������T�w`FXጉ�+�m���v��x���0�[�(e<���'P��h�sob���������==�g��EF�ZȍL\�ۘ��n�3ɿD�T�$���b䝝&-V�*f��(4V�L2��Fse��5@L~FJ�f��}lE�Eե�Z�h�z����Vo#�bھ��Rw��֭n ��W��Ȝ����t��0^R�'!O�����^�8pG<���?V�Ŵ/xƼ32LOX%�p���p�d��i���2cIz7__���	8G� ��l��4#D�gý��S�1)�nR7��G��d~N��'q�
�O���V�T�?귄�z�n4�Fv�vOB��Y�3�C�=̃��7*�ʗ��S��YAAk�X����\����^�m��E5Z@F�
|���f�6�"�qҸ� �1~�~�	(����K�:�b�b��/�Cn9�vSg��P(��X&k���BC�O�[��E���,G���yPۢ?�����W��T� �Ɉ��d�f�U�^]�w<�xO���^kQ����y���?٣�'>���}�{af�ť����06�+݇ER�E\���&_�Q��8U���6�%� @��Z�' p� T��	�t��(�l�hNk�y���Y��/~�qG!����+K�W��Վj:U�Y�,'�F�h�Pp�؊]��Z��o'�����dXƫJ��Rv{��8����*�rj�g]=�y�d�����1��U|�D �<N\��С�jĠ]ow^�1ʠ�_#/�x^���-������!�Fe�~-��%0�s۳ǅ�4������B���F��W���r�����ֱD��� ����u:v9al��"gBX���q匹W</V�Fmw�M����i���5Y�����\D��:'�!�fs~����)�Wp���R}o��	/�B�B���	P,:+�|�X��4�or�H��X�ؚ�L��Y����c�G���z ��(u��t�oٱb<4�����D���V=�2kZ�aϩc�l� I�'�u���y�q�����ݘϮ���X��_;6W5�U\��f{Kp���<Ξ����l��/��W8��E�Sr�*�" �Gڀ��nbn��!�t������'[c���D%�8���U�]�~���He����W~G�@a%��֞�<]|+k����:�}tn�uɸ�޼]�Ҽ��"�����0�;�C���l�m��yB��8�Rr!s��r�c�ɐ���_�W/"D�2�[��Z�Ϲ�U<1d�tŕ�D��3��|N���X�W�J`'+�f���GK������n�UA_�r����A��|��5�v'ӈ:�7�9���%�k���oY�r��X�\f�?�����~��8��;���~�q�>y����Kߑ���z�P��{(GG����@���=y�1��9���m��\�(&���h�	�y��O3�n�a�AiKZxw�^�/߸lq���cn�X��Y#�rV#	�����˒N�
��hLf�t���-�����N���C�q"�Cz��5H��e)�d�N�
��&��r�!�o\{�N��`��l
���E�W������''ڏh��]�yꛨ&ې����T��3�`�DO��mY��j>B���)�������+��=}d�ZNr��eAr~�P~��0��v쟥�⋚0���e����굒W�f�N��i��ow�=D������6���5�	i�N�ݼ�#���\���Lo�� ����GS_ݚ>�/y6:�Kz����~}7pÅ+���>Ѩk��a˻Y�9P���8�;[��QɨMCZ�/�\�?��e-uO�(�\�ס��+^E��е����A	��q!��Î�����6����LE�t����0�~�4jW.�夶����7���K 0�ܗfHt�UCڧ\M���W�s��ZU��̎ek��ޥ�)k%-���)Fi|��Tn�$0���UE�e\63%@Ӵ�ʍ+m���J��x��s�7�Ń:�sF����%f8��y�Lbq �%ꛨ�pC�[qu|q3"	n�(���o?�Fdm��ZJ�cB'D����@���Y��)�$
W�ZQ�t����æ��yB����'�Φ	�rqQ1|7 ����'�;`"܀���9V���I����aN)�����U\|j3
l�j���H�
��7%��|;3�
��yTJ��؀Բ�^N���oX�߸�`qc�p�����R������*~tD/���^�nHkN�gؾ��kx�Uo�뙐�<%oG4S���6��t<���F{�:��5W�Za~p��q�y�3����t���!M�-QI���!V�"|WKVyl�� ��hhW1��F���v7�¤�se�C�_�>��{����bjX����T��1q�������%:.���s�S�f��������ҳ.�v�z������άП|���<�
1�T1K��{��)�}�B���D�ٿx�XS{������k/3�<h<-Z{\��G�����\ �MaoLY���K��-{����D�Ҏ'���Bk��P�����?6�w��l%1��{��uW
���a��/��O�a��
~h_����)���'�i����]�]n�\�m<_U�#L�𗔷#oU�N�[�e-d��W*gr5t���[�kc|馌4�X:��Ӑ����n	υ<g����Vp���x��#=����]~�p*�yW��3��[Ɲms�$�E��q��H��-���Q�H�=X� KN�:�	)G�`G�RIؾ�wdp�4�h�'z��*��ޫ�f�B�Ow_���ǵ�H/����X�4Z6��#^�Ac�;ʔ�r�m�	T��TϾo�Q�/�j���ݠ��_0��*��a_%c�+�K4�z�M��WȖg� ��X'� �<���%�$L�R햚K�D�0�l� ܞ��7��r��I/�v۾�s�����y`v�`�
n���,���|���չ��&|` �`߼�2_K>�
+i�����fr�>�!��>���!�e�"���5�g���)���8Zg	*���`$�Y;����[�K�$y��i��2I�g���{�b�����T#h����M+�c>�T"��]�Ud�?��z�\�0�Lћ�3='�KI�X��f�l�ϻ�9�	MNV_YZ���D˭��˱#`,�ϛ���X��F�o��x�r�}E(������8,�~^��*�ʪ�F��B����[S�),��G=�N��3F/#عj�����X%_��+�)<U��^�w�e���MP,��j�˫N��P3�}q�ey\)�y���3�����v�|F�=e�4��rv�؁~���4�kR�%��ש�v��R�空�Yi���6r�4��D�3K���a��8����R4�4sw�C�s���X�����׼�uI3��0��n��']�W!DAj�����A����ck-Ѓ��=�_(O��}$e�j7�	rv�+�ͧF}��_�>��K�N
ԇBD��I�+C^y:x�v3 �<8Ij؂�r��g��[�'��ʑ!1okx�;���ٞ7�j�yM�<�#��6袳�_oӉ�B�y�{���[S'�2h����O�q�P��º��k�6�&ԁ�Y�>0ĄF�=.4c��u�	f�,X$�A�b*Mq%`��[�d�_Et}EBv�nA���o� ��R�O��v�Z^	0���K���޵Pܻ�O�LTn#�dmh1�HϽe�7����R,�Պ�͘�]9������o�$p�`f�W0E�*,^��o���@�lI����h{�ET��@㬍}A��lX��}"��u���X��ɹ3�4��hKx�J�aU��W%ķ	��H�p�HhH�t��ؕ���C0�貢w���76G�RR�r�&�K�9�w�����Ճ!�0Z��G�,�L�, �8%|�|�Ô�E�zF�c��2H}�㉓�m� ��y����K��5��$.X3\v��~hD�iL�2.xߝ�V����@Cs�4�.
^%K/m� !Tv�<�
�<B�R*?O~�Jˮ'��N����Sl�c��l�.|�:K�i���j
������������uVNfk�z��t�=���$�̙$i�\�*����R��^�K�1���C3za~� �����`�=�u;Z��mL�
�t�C� �N7��Un"<�H}��۠�'�|靎�D�W�R�9��U°ޜkf{���q/�1m9c2PÆ��N��1k?��Ǣn�����,���} ��9���6n,l_�?3�}�ǽ�d7����`�H!rq����F�d�m#��R^ڥm�ې��L
��6e����(3M��^�
��Ɖ���d�_�ə�y)B�<Y�((�b���[��P�G㏓�F4gs��4�;6|J廸���|}���� �O)�L���9���7S�){�a�=��mHh�}��-YOq�=�)~�A�4F��]�fL���dƅ/7��ڗ���sd��B�_V-����~P��E�"��LZ*�AH"�c�U��elfqm�����R���zs
"��Ͳ'�����;��g]���r�d_�4F�-�������'w&����=	�ƒ�����0H��K)G����v�d4�ŶWL�Y����Vsm�d�hR��&�
U+p�K��Y��G;?�qV�/l(װ6B�'�_5h)/�l�jXD�`��&*�V�~[���-N��]���O�C���
�"d���l�����jӦq�ϣ���W��]U�uJ �;b4^����ڽ��T4�f�??p�b���N�]=6Cf��ZR�ѓ�I/�_]?�cB�!��y�Wӭ6����j��Ƚ9	� 2n�mo�I�ߊ=O�ci��~qn�+g��m�m�F���������sz�$��(��ӏ�!
���!>VI�	�3s�]I�x��x���3�2nu�^;\f7���UKcp6@�a,z����Zz,�t����3k�w���U'��Q,r2ܫsB�!1�0;��7��1��8�lj��K�K�h��92�&l�#�����oc���U��h$�a��DE�/Vb]E���1�E�2�h�/M0T�8R�m� ����ۈ>y�����#Y�2Fd
�;a��a<�#{��x_��Qb�Py��3��	C�1.!Á]�o+D�t���8��_pG\�1�f��*{�*5\�Ŏ/PdU���d�r4�ͨ�Z���A��vpA��|�G`v]�0�GD������8:eiM�йe�Ƽ|�M��m�)�O������ȧGt'�>�������0$�6��%�}ic��J����] �>V���a�C�-�Q�K/���A8N. ��M����e2�9˓�̶�5=QM������H������K=�S!�ƞQK�%d�ǗUL���dj	�9�j��:A�H]�n���t��{s���I#��/4�6��I�z�ӒZ57��]����
�.��i]A����Ki�uԞ�n<f�������'Ť���\������y�{d\l�ì@����y�T��c�,7�x@^��4OՑf�%�x���;�YE�Ӣ�о����Տl`�H�?Bբ���sGfC�[��"����S���O���U���k�װ/�ѿ�{z�A�M�}��%!y�)'�q���։�K��x"�n�γ�e4� ��0����%�0\�Њ�q�~�b��B��2�s'�:I�+��}�����R���ฅ3��VY�g3:����`�����u-G��������cB��"	b�2hwK���$����WI��EM���f�^i���z(g>��t�l��iL���M�-��N ;�ɋ�v��jŞՖP8?�ە��$���K�Pp\�X��� �X���A���2K�,A	�7^Hi�;VC��e���rͧ,��{	��)'��o�d�s=k�e��"LIfBP$G��-}��D0'��U����_�g$[{�,3K_v�Ec%R�L��`q��=����^���O�$���ź�D&�+��kѫ۩����ź&�%�(�m�.����ƨaQU)��d�,~F������g�KI&�E�F����~ׁ���pmׯ�I�W�����D�JJk�\| ~�$��B׌�<}F�Y(��=�����6&�L��+Q���Jx_a�~|�V�̍�E�M,H ��hV�[aeV���3rdU����si���&��"1���4O����!�F\���T���v��m!�x���:�S���;̓-�<pr������7F�� :�Wo!O߰�/��p��};7��Θhjfzi�ۈ䦙���	�]3DA[����%�.0J�u�oA@ w���Cm��+��h[̆'�I5z =���8��p�J:��䷽�)�Ɋ�țތq~���C���e�lQi���Lk���k���198�I�0�����2�.��+#>kSa��:�n���X>���H.�ձ�u���v���5�ze*D��5��t6���`ad����a�����4��C\7���I�F��c�!����10�RG>0�F�7����S���Q�v���,�}+A�����"{���1e߸ ͠�Җ�%������{+����������+��3��y/��[��H�52g����v���Ӣݼ^��\y,�_�P%��V�t��)��)9�g�Z���6h	V�\sX&�Hyk4e�bi`�%9lu�Bp<n�5�;��x��o��u䨋ma����HS"*U2�?�����qZ2�;c���51ժ�xbmas��P�]r��b�x�:��9�Dvr�rUՌ�k&X����R�f%�RS���ã���U40�#Wj"a�X-4|��ƀr2F��s{b�۔n��e)�3��2ym���n��Q٘`�[P��da���v�%�C��X%Π�����	B7�Wܼ��{�,,u6���'�����`���;��C},m'2Ҙ�9�r�.8iҵ ��J�
hu�~��@o�H�u}�����U�К6'�}��y�ͳi/z����Nl�����C6�<9���L#r*-�+Fle�)kWv���lV�.x�יğ��k�aj_�ǩ����ٌ�ea�� ��Ѹ�*����@S�������R�M�I�ñ��mT�_� �k@Q9FhHq��*h ͦ��1���N=3Y�3c��]��6�lR�SY�i�� K�G��5��u�(\���(���)Ϊ�ʙu��7B�]��d�t(�k����aD�kద
���R^t ޺ʏ��Z��_�b�̹�]��ɬ	�_��:�3�ȫɄ�������1�N�aiM'Jg;�e�%p	����>M�(�Q� N{�	��"�4s㳓櫒7�\_.�Qͮj`-����o����W%>�w�����
S2�l�T���3�����k�2�/a|��w�*�ǔ�6U�a=�Ӊ�kI��lNAiZatgȖ>|�����0
o��^�!�@�~�;S�P�z�Ry��+�\��d(���$y6]T�`=�0����Jf�}`=�S�)�ÚZe �%�<�\F�^��aB-����c͊$sX��
�[��{TsT��Ln���ri)�1�L�FM�bH@Zė���jQ/QA�Q�bş���Y�*.�%D+��P-�����rXd�KO2�{ڿw�����G*^�.}�*�t)�Q}ݵ��|ap"�g2��q����vf]x=�M��(�J0ʢ}_NJ:�Yu��#�2�B) ���ZԢ��	���eajx�k̵���������Uԁ�oi��q�P^�1!I������B��U��f}m}�i�{���-�U���K����_^}��0�b��6����/�כN.�'s�S�ކ�r(�	[hU�	�VS��4���JY;���i���;�e����g�����)�SǾk�U�3b{�[����q9�ߒ�_��iA�2��O��V��øO�����O��h�{^�2f�����huE�P3*�5WB�թ�K�/8!ޔ'e��s_j\������<��˗���?c���l���9p
s�����(PZE��!w'u]'r$A�YLe�U7J\�������ZM�aB[Lp����~��`�Dy�*�r�%�����<�s�X�֔�$N������ם�0Q����Cۀ�U�8�!zbQG eI]E�yT�rש!A �.[U~�����OvPn�9i�� �����2�"�&�$�*\� gt�$����Z��e�`�dk��η����s/�5Zmٓ�Q�NT7>��2�F-�Y)Y�i�;�A2_�%�*_�tA�Q���-U�.�����=j���Iʒ�q,:�Qc����A�H�RcjxrU�B�p��Z.w�G�X�^l	3�*�@�p_,�p�LV�f�s�r9ʱ\H��Kl9��P��G�p�]�X����X�`�B��f�:K�J5�g�����'� W_&��x��*q7�H6Y�P�w��H�^YE1ךl�`B|�f����1nxfER��r�]9X_����;��O�jgoTWl!����>خ��\�Ԭ�$6���ή������vCSL>f��-Ҁ�a6
�Ix��\��5�v3�W}t��w���_�7BY7V�6��Qh����UjUш���Km��:Y�ɤ��2��)n&U�h
#½CJA�u=�t+	(�	�{��C��bQ\�Roswb)��r�4�j��?UR����5�[��_�u���!Z�g�DR
���l���r��)�M��|B%��
�h,��դ���섓�@#�T��I�d$0П)O���s�!�B��[(���՛����`�[b��;����&�����r�'7g��)g�y�!lH��_�:�¥��M1$IF�ޖPy��_F�U�����ϖ���_S�\N�U���p�����ڬ���VlB192����r�%�����k�!e�!Q( �&Ν��`6�ho�>����C+��s��E�u+;�C��F���h��)��|��ţ�E)�l��%IY�7�����U-$�����8"@����+1��L4J�59H�y4�aX@.�,�a���t�.�@�qǷw�k��H8�
zԠ�I���? ��ꘟG�[Kw��MP�^x'�[�܀�i����~v��Yg�$+���(��$�v���$ey�gK��)��.:c=U*`�c"���e�/���LɊ��]��voPT�!P�r�u>N��T���F�}�j�3h����wi�)v=�94(V�).����CՇ&[�u-�z���� ��Ur9������u����(��oIuR�����W(h�&�}�>Z��v��]VP]�N�'���,�X�⁚#i�)��k�.OY�A��k�_R�@I&q�a#����)�+z��+�+%$���P���b��\��'$�t����Va�"��C�ҝ�K��@�Fd�����F��!�).�y749��H���-ЪA�P���V59�xz��<T��X���	��d� U�8O�IbX���q)���,��IgkZ~ߙW�C�U�mV"6?�-�R(8�R����n���n���lqt�kx�H�
VM�wz���^��[�r�8}6h���"�Y��q&fW�M�9�|ƌ����`g������&��_M]��V0͑(�H.��ߕ���gv\Ъ~�?�sg&���<�ۗ�)��}?��c[��=�7�i�Ơ�8R�OU�yE]S)��|@���7�e�|���=��	a[|쟚'cy���Q?���	UD:v�0��f爍�c1Y� ahu�c:l'��-J���J���u��<M���ܺ���XG2������e�M�b��(H��PFw�ָM��x�a�YaD���/n�߇h�:�$��2�cw�B��]�i�	�S��%p�S���P���m������P7F�6]�Jm�Z���<��e��k���$���V�8$Բ{{Ro������%i�Hk�*ނ�vH!L#��A_��^I��6�_}��~�~�dL)�R����ԚK+5aZ��E{����.B���$��کm>ы�Pt��Rm���t����۝���)#~ R^4�r��G��c�֦�l#'��vY��V�J]b۰L��B���p��	�c���Gz
>�W�1YTaYf���/�X昴���́���[��OȖR����A~����?���S�(���v˲��I:˃U8��h�P����TF0Qy?ι��8�V?R�_<�y&	�=�8����D�rX"Hd��-r�G��u�٨�8�ao,�V�M���]�<{j7e��'�3�KJa�&��A'�5�F�
������z��Bj&�@��@eE��$	ښT6'���*�l*��}��j!$W5j����'�35/���5w�L�r�X�b��?J2r��9����}��SF�-2{��7�1��t�a���Ѕqڸ'͎�����ODI��>�DC;r<����"���c- ���[,R~����8[:���b���$��zX!��s����b�߭nC�.�H�T�u��؋�Z�φ)��O���O����B���{N�|rhN��UˏX�%Ozt}���(�-tF˪AT��,�[U����n �����L�w�3��t?"�e�UB� �����/�P���4	t��K���itT͆�_����.M�W�+�CJh�km[7�3\�ٝҜu�J�C�+ɝF[��N�RKʌ�P>��oھ�[�B�b:�Jh_�c��)�U�5~m0�g�� ��U+LkR���~߫w�*L@�L,����ۑ��?1���i��Q�AY��p�n�%2Lp�/%���.7�[s�?ն��.�d?Dn"�?��S ,.�yƔ4�c�W]�w�u*��\�jv>���ơx>�X��3d��sf�듐^�ͽ"o=�RZ��Z	nH`#F*�v<g�Ԃ6]���*8i�}�#�p��w�m�ĞE�.ε5�"2��5y�/�j~S��aYC��O3V�<������FU=��T����B�k�
��[2���n�J7�b�B������.�?v>������L9�9�EU!ױ���Ķ��}�~�JI�A�J��0��ы�}/L����]]�?}�'&�G�XZt��NZ�!P>�����Cq��Rh��E�Qq�+%6+?����=C��$Cc��\�)=�w�[�L�'�v�2��[ݞ�DL�D7j��%Z?h��u�3hʸ��@J��m�YWv�Fo��!'���{��s�o�`j�w@K��#O����r�7�κSWCi��@h	�üJ��E^����/�Wc�*����o��y۪ځXcl��l�� W�՛�� �A	��Y���E����p*���vᣱk-��+L|��#��Ї�������NT�F�����Zmڗ�"N hO���Ɩ��|2'�Z��r��5Z���I7�{��n�e�G#Ǹ�[��?��|���p�l'���b����a��_a՛�s_����Cu��~��M��<�̓�XW)�ފ~\id据�g|�m�����#��W�2R&�W�6>H��I��w-OC2��㨭
+���}OI�ùL�r	.��v79'u~��
Q;ˬ���ᕚ.��A��g۠��.��p�)������|���%%�B����h��Q;Č%R>d����ُ�X.Tl�"ivAX��n� ��%�ﺿ���5�� �W{L:u��p:�f�n�q�a�+�-���_���b�}�y���CǌV�.��ǋ~2�����b<8�׊d.^��8��F��0�_�.����e�<q�`n0,��?�L�Ҭ��>TH��f\�e����;=A����>l��b�Q8�B�w��ʺaDap�>��@�R|N��N�� %{1�<t������k"�kz!ֵ�+����6�����(���ᜅ}0��'KK�DS^?e�m�)\_O-���Mz:9��˺g�	o�!*�X��_0 ɻ�q��|��)�;8#e��T�����'��	�ǽn_�7*�}�9�<��[��K�����G�~�1H�����_�%x���}�yhK��]�?s	)��n��OӖ+����I6K�{�u/����[h]?Su�=-W��>�"7	��ݛ��1D7(O�G)kN��m}�a�:�DnA8������.^d.A_��70��y;^%} 7�E���FOlU��ǵ��aG#��:�]7����I�dCd�8@���GOG�Ǝ�;��A(jʜ
{w�T�"-�#nk�K_��C��(�����bs��B�,�a46�t����(�.]�ѵ'��+���ֵ<���_��p٩�Yئ����󲮃s/~"���pϞ)��$Mh�[�=������x?$�|�]H|���N������w���Uˎ�U���j�؏�-���*�G���Tޖ��'�3q?T�Q f�ʽi_��t��mZ��]�o��c�����!����?�@�˓=�;&:�Q��	��&�NѴN˩���X�����߁��,�a��| ���߭�U���Cײ7u�%w��:}�]ꆐ
��U}�lٶc�IK	�5zA��~ �+�$��][��:Y<����gN�^�R����
���Լ'R F�b�j-�g��܅#g���b���%�Zg�fk�x�\+,�P�7��H7{�#`vxL�=���1S��U��ښD`v0�ŧ�;�`�� :ˑ��X*�v*��Y�#�"�V�q���D�8U�qN�kV�oM%6xgT0Z9�5v}�q�qV0����7�khp�&5��-u���	;�1u{�	�N�N02�,5���		͞+Z/A�:�gJǕ�����- ��Vڛ��c�FgƸ���	<DG��y���ŕ#�ۀ�^�xV��~5�:6֟�^$�#bBq\�OOiZK��Gd
��?��VxN"�P��îW������^$�� ��u���B�g!��2��1�W� Q�8��[;T�kꅆ���9��>����m�nˠ
1H��ʬ^>�Lj���e~�䵅n	�,�˱����ZT�V�Y~���b\2[R`�oΈmU�wUy'�2�M�VL���A�g��	ꪌ�J��(����+-f�,�k���q��U��7������e��BߥT_GS�HV����Rƽ*,a��;jƁc�������N;:�a�}��8�N��ZH��d�"3�3�V�����v/���hy����IKWY�������7�CۚF��6�{�&��Ȭ���R �9��X>�\*��P�t���
�C���k'�o
+<rd��y�]ʁI��b}. &,��:`/x	qU?,ܟ��������rh�|���Gx��~xE�ϭ�]|j��W���x����!��@���}�)({���m�7v���Yv��h07<�g�%{I�h�1�W��>W �3.������kB,�����E�`p)3���"c�§B]s[�)���"�����uR�x_R�5�h�}"6��`:�	�Q��BC�V%\�����Q��JI� 9��]�G�(�g��(L�1��es^'���Di�M��ם$���U!%��3Ro�k���ljT�3��g���%��[m֌u�~�]�x�5�QEJ�9�N��@ܛ��ad7B��Q>�FsЫ�v����%��>L�@��*!ה���.���5�,�#c����O��X�

AM��9X�Ma�Ĺs�}r�ҟ����[��Dx��[&!-��JG���Z	��������������!�Gf�Qi��I'�B1؅_��P7���$VL���+}z���eQ��scpd��+�7\<|ws� Mw3b��9&ξ�1GXAs���"�v�����R��a���Y-��r52 ]Z��q�Q��b5ׂ�r~J�s%�}	+2���mSb#V�ŵ�����A��*�_�T��d���-�F1�O[,ȃ�~���􌐻�c�U�N@�ix�P��0�`6� '�o?XQh{���ln�\f�U�Ӯ�ڙ��<FtԞz����0>���m��h������������3�=�
�J�u�_m�q�nC��Ğ1��.q�yK���.�1)��9��x(E�F>��!��h���ٓ��r�������-�b:��C��U��J�-�����WG��_��́�E�/;0h�7�|9��V^kO�>��y��OZ��Ni��r��^*]6��*��^�,.H�e�As`��s8ʅM�T�������ǽ#/�Z������*����sc���t�k,�,�mPޞ�ܼ���Vp�5��>T��#��}{��~���I�'��u?yuYn�<�L2��,�~{���v�wo��ie���<��SF�T��x#�(��r�)r����[�_�y�/7	�_,��J�Z�IAP{��G�M��K��wR��`�DU~�%o`j2�����.��	�G�y�(;�J����`,� �^�r�K�E��>GsH!����H��4~xN�h���a.�k�p���6D��:��׃EiTk��t�I*U4ݠTtBk̬M=+d��}%X�%�'Ǝ�ڲ,��z��V#^�������N������8%�`�����鍶��{�Lwڂ�rU��=f������C{�y[}�B��HVd�|?	�oQ�Wa�
�V<�Y7�R繞���6+$�КI�E`�m)����cY�q�ݏ��B��: 	�s��ݙ*V��i�����̄l��h*�y.�a�Y�`��IQ��"5f
v��+���Y����ѹ�R�R�G��]U��@S�OZ"M׉�\lb�.�AtēH��pI���KG< �ǿ����a ��0�������wԅ3b����W
�Jf?f,?'�"�ۖ�jc6���X�ڐ6���������0�ݗ���u,T_""��V�J5�����y�P��4lz%�cN)�W������ |��嗌K��,�L��}��e/�R�����\�\z�������n�D������:�ɬ���� 3g�)�o-�zK�ֽ��P�x-����EĹ�<��ʒ(��s	�t`M�%����y��\�*�`D����`�J�-� ń)OUb������ d �5p)h|ɧU�ҘI������f��Т��m���FJ�1_@�U�Q��j�����F݀�L$;�{� ���@|�N��l������!���F*�eS�c���N�\#����Sy�
��w/45C��~ߊ�6�ClP�ȥ��]Cm�z�Z={��/ɂD��^��o�+����~F��9�w�ٔ$�ׇg���&�;�$�"0B�B<J�T���e�1ql�N��
B�)J��4���K�EQeg���50���9vE{��u"����/�D7���1/�c�ή-�bFm
@�l��;���W����ִ�:���V��؞PS��)?0ě�J�p3&�[����rШ��i�/?��#��=�ʄ�inb��L��u����0~&=_hu%��4�琞��%�8@�����Å�QZ�P�ՈE=,w\�y#�����1�G� C�����BT�CuJ�� Z����)�k4g(��՗k���[ł�\l�I7⛳�_6d�)p�����7}�Y}��s�����(��1�O3S��bAmDЌ���S���5�#�������Q��쀴�Mh�"Z"�7�gL�U�Fbu��/�`zH�� {c�&ۇu"b�Śr�N��A=ƪŴ����Cp�a�Y�+��d��:�b�� �����6���;|uT���Dץ�.t�z6�3AJ��׼e��K�K�k�y&�pS亨»icB�iO1��7�3шhh,�<��'#���˝�S�z�b�`{�[��U(U��|�PMJ�
���J��`0�+�:%-�h�9r2: ��`�<|��B���(S�*W���
_�Q����Pg���SQ�k��hcDސYϱ�w{���T��H�qy$ ^�G����jѳ�?��(�@]��~�dA���O&͜���g��i���-|��Ш�)���$7	!E��|{�l���%�{�j��S�����r_e�$T���b�6�0�/
��"2����@֮���X+�B��X�$�)�����K�8([nB
 V>��*<�ːЉ0j%,��O�Q5��4�@\&ݽp�s�Af&�+n����!|�X�O��e$���yZ�ӧq������À7?0�ukC#�
Xe��AeB�y=|��� �E�������n��jw�¡ڿ���<ôyb`>�S�K��Pl��m��1���{��tI��M�Eh�"�	Y �6�".�%E�KZ�D�zx�p�r���#B;�q@Q��^M�[�0r"$�s+�uU�!K�Ј.�ߣ�(����9[>��+���8e�I�&Z�[���H�@7�J�`Q苠�@v�6|�Hގ��e�O�HE|�L����a{�Z���0E])I�t�wò�ٺ�O�k/q�Y-����Гc����z����_[K�H؛��7���EQb�ۈ 4S)�7 ����%���G��,�	C)�D�ĥX �w@@0����������ݾڂ?O��2]K�����L��+��}l��Y���-�A��#�H��ȆֆO����ȸ?�>�+����D[n=��V�����g�^�`���i\26E��B��Cr��$p�f��"I�6T�Y��☚T�\�䕥T��]uk��58BV���G9�?�@	�Y���Q����\i��{N�V, �J�d�$ľ@6B�O��LA�aaqN�k�H�[��D�n�g9EH�d+����؜5�k�uC�y���̱���ݷ���Ry)�����攒���mg�X�v��i��_���O��m����.7 ��ě{=��z)́!4�
ß���n�Lh.D�$�q0�lf1@�t���i'�����Js&)ߛOX�Nt=��^M���o�8+�x�lk��tP�9=��"��/'�4���g�s�J�<>whg�W!�1ktI�}�k�{�7�9a���~p�YP��[ =!]2�ş��)Q}�)Wo�/�P���9��M�]l���A�M]i�Ԋ�n�8e�m�%3�^�3��!�f���<Y���$��(to�]�1��1�ҫ %���q6�C���5�	� ̽�z���QY�O��z�})N����=�~:�,Th��ئ�UrZH%ǥ�n[��]\J�����YX�����|:��O[Yi�;�[�Vڸ��X_����`�ǈ�/"����Kdmf�#e| ��:ҺfC�	o)|̰���_�c�[����"y��~���6�Y�u�'��zN��,��{�hb��oCo:M`�F��ygm5��c�0�H�^ڽ�^�lul��x�5t�8{�MG�o�L����H*�4�$~�C��1#��h��/�̞`��uI�j�sp�l��^�-�}���`�E^���r��Ԧ�6��DO�q����-:����	cW|GJ��xQ�,���4�Y杙B+�nM��
��"�,�Q���'ZoTê�����I�+PIiK�Q-?�O�к:\F�b��p���aFE.�>�Տ%��6���w���i6��c�*c�b���L�T-|(��#=i8޴���\g8��`��֘[��S���"�à�hn`r��_m>ȩ&Z�MGk[�(��ǯ3x%�l\
�#��:8P��蟛���V�bR
-�I�
ƌ��$���K}�ϻ�T�j����t4+�P�B�r�J�-������X��Y��I��
�&�s��t8���<����� �S��mۮ�Y��h�/��8hBGջ켒�FG�[ñ4b��3�j�&~�6�ݤ��.P7�����t�ʕ}�G��Ge��*�g��]�בۺI\�ˍzA�w��.�N�0����/k;��d\��u�w�� ፇA��~��j���������J@W�}Ҳ��p�X�D����ݮ�3M�f89<�׈�k]ĩ���]c�K��.�� 1˰!��X7~��I`
�^Y��A�����\�oѳZ�-�ׇ����ZN����{���*H��`({w� �S�?�/=�W�����|J�����4�� k3a���Z��Q�^1�Ƭnh�<�7 �)���o80�p�29_u�Wܓ�h���|��1B
Y��(�tԅLB��6A�Qu�#��HE��r��k��c��)��Ǭ�:y��(-,ՂJ�#�	�b[季�H��T��)������4��}�n2
G�̔���A�.R���1'G%7Td]�=�F,�!f�9�l�b�O?@@�<[�O3�ŷ�on"�Aӽ�
<��3�Ȟ�ςb����Vo��
&7�y.�P5Z\]A��D ���A1�z�f�/B4�k��Bź魉�8�A�ΟP���w;c�.��̃�/F��z 7#��r�d�������bn�����f� N�3�����M+�o�E,V6ح�StNe�au8$��>9�}�͍�C���i���Z/�v��5�RUWAp��	��5ξ�7t����
�ux���1�+�J�Jd5����l;���7صf'�*�T$��HM�֒
F���{۴�^eJ�J'aL���nM[
c�ma��M��i�jJ�~V�3�ۗ�����L8 �/C��{�MFj��F�¼��'��/�`�Jd��<:�!(<�j���w�a3;�T��{)'$zdD�[�s䊃���y��?�7!O+�*mٙf���9�Ǩ�dɣ~����+��s��H���":#�@�K�;�>�T�a�y���)���&���"�_e���@�9��dqHM'�F�e*\I���+3v W(�]c�\��<[F�R�H�;��~��W�AE��D��.�A,=y��$㒲���9L��擗'�s�&��e���R��$���C��ϋ�	��&vy8>�' ��B@�텥�����ccЂ(��hZ��4�V��]�����{��C�pk�k��Bf�.��_�ۅ>&�k���v��i��^]N���b0m��5ч�vH�Г�4UPA�����=�)�E�� ��i�^l�������԰P����zn�k�I���n����
�m�H�nwS�W�O��A���C��P�Y�<E��x�5�sN ��^H�?�gᇆ�sO��'"؈�!�kl�ʉ~�g�xK�����p�q^B�1�C��@>�Q���o�����DϬ@����g�UOY0�p� ������[s��z_��k~>�,�pavt1���Ђx�0�*�*�H�c��p�S�� Nв���Jvخ��5\j)�!��.)���5�i��Pi?����5ԛ�]iBZ�.wSR�����E�y��� =[�T0�0�9�~���Q���Z�����6fV�KؔZ+�����0��mq�R�nT��0:_�tb�H~k2��5ۃy��n{HưG�
� ���q
�l���B�5���Ų�����l���p~5�j�Oƽ��kP�G��i"9@����~@�M����??X���t�������O_��s�_-
!9�<@U��1����5/P����Aa+�C�'v$��qN�!��d��A`��A,l�"� ��n�����V'������X��A�g���ywq*ل�S�zz��Pe��`DSs��\T�^��۱�K}6�o˥Y��;}��UG��˂�4�]*刉H���.�V�Q{��\�Q�OeRy�SG`��R�M�׶u6�������/|Z�o�?7�;��=T�����7��1�d��w����S��]6x�ݣT�A�Y��Ȱ3�ٻ�0Ǩ�{�5.���`�#]U9�Z�i��m�����~�"맯Si�m�-լ�
��0=�	�=V��>(�򞙼��vxq��=D\��u��9�4j��k���T�[�c�ґ�<Ƿh�D�Ьa�|U6&��NAk���q���0
Y�@o�_�"�Dࠒ����Ѡ�;p����p#����V\$����|��l�D�S�Sbڐ��m��mF�m�p3�0�A���(ey���%^k]x}h��L�
�:ij���j�H5��Q��[,�pu�fGM�HFƢi*'u�3���m��v�v��_7�7$eL:c	O����� 8$�����îY���`C'qE���*���%u@#�qo_�^�&��`.����U�X��SH �H�/�g3����y�HV��a:���όXծ~l~؁���1�b{+k� �v�����W���NYx3����|dzFH�/�ѩ���K��\�>M4�M�M|g�/�ف��y^����C�1H� �_��ׄl���8���"��V�*H��!�d�V�.�c@�}���qo�'/���a�2�&H	GyN$ƀ�=��xm�<�p��Y��K���SKt2� �4���7��Ʊ�j�N$y�$�Ao�n�aK'b����J3p���n���e6�ݐy�c�N %G��=�-x����xྚ�}y��27|+o^��ޅ����^�f�4[]-��;�I�,-���ܵGk�L��_�:�|S7���
�:H�b\r����Ϳ
s�uRԔ����e�_�o��V����㛋H�R"L����g"�ʴ|��d���ajZ��T$�C�عE�=���U��g��a��|�>i��5�`ˈ(gQ��+!}�ND���r����j+�MŔ�֤�;�!�8#������M����������zm���,�y��{C,��h5�_�kT�9�����>���a�[`��~�:Zijm"��1��>����ʨ١+h�%�}Kʓ�%WpʋSC/:�)W�Z%��pɅ�d�~��X~�0ة�ī�ݐ7�^�}�m�{���K�q}W1�E�.��H��( �/8su�y�_�Wlf{4v̚1��uʮDd��ES�b���,��[��e�-��v1U/�����	جBC8эT��O��2�	J�f���w�Ф%z�8(md������Dt�Ik��k�M x��V��w�Fy��ZJ�*,%߇�������ahh�[O����d�]����n�b�)�X{a�R������5��Ӗ�>����l���{O��%fKQ|(Me8��!��ء����I�|R�VHZUϏђc6�V��ҽO��^�uQ�C`��2�̪(m���XE��ݚis�몦]����\�$ɪ�@�Bg�N��$����������+i$���$;�|��0���f�J_9O���o4O���|g��A;8�~}v�c`Pv�j���G����&�2�8ҏߑ��N(�N��c���Yl_Ι�8��$gY� ��$W��P#1��j�ֽe#�:p�,Q5w2܋f���	�a�/��UfFa������t߷�|��M�Lhh��k�q
Aa�nۇ��/��5�b�}��8�8=�<��A�8X#���kZ�$º�l�wJ��M- :�hq��E�Z�wW��~����@�G�]Y�*��JTR��߼pI\���G�u��'Ϙ�i����b���%�_NN���N H1��Z}�'n����@8g�)�i�u3���"�Q}��Fbma��PP4u�өCa�:L� �V�����jf-U�D��+1�FE�1 ��A�9�
ޏ�h�sTЈ1ښ����~�Z��W)�_-�b~+
R���C~��?�
#0�briq\h�RY��Z�
�S�Bq�2M�K�����`j�qⶡ2x�D�Rӏ�n�T^
;��Ks���\_�g����O��M#҉��yI�F�C/`�u8�ӽ���V�����[��~���ͺ���	�i��u���z���=x����F]&�X$���.�O�N�8f��%x��Bnv��2;��h1���L�[F��c��vyyx�2�=��|��R�D)>�?�r��W�
��T=���.9���z1N8����E�iv�i��b �h[��F�ح,�|6+so�{�k�N�=~�挭�o^�)'*R�+�|���4\�|V���H�v�GU�>/�u�~�d�}�\n��x8�"N��.����j80�p�Q$�!7�`���Q ������W!��8�g� �:��$ǎ���[�Q���v|U8N�4��wt��ŞF��$�m<A9��Yп~K�Ց�F�?�`b�ɾ�(�~Zs�1 78�m���"Zs�,���ԃB��!Q�C%��.$��;%�߮�M�n���2,t.��;4f7�l��e�B~i���ϣ�B�PG��:��%@H#�~��xAEu�J�K��<fz��pJ'���m+���I�)Qk.(f3Й��X��OSɺ�2������l���ҡ�/ˤ���Y��^"�W�8�K�&LG�T·�r8K��~+�(+Q�2�Ip��j0׮EN���(��.�B�ѓ���yG��;Q�DB1yW��q`�
)]Z��\i
��(E4�,GE�]�s�4���5�G��mC\`3�D&���B����zy�-S�&�������o����*֫{�jJ�9��K�B�3݌��n����Vk��?9����+,����R�ԝ����x�`�p����<���>�6 P:����8�@�~�x�o�lB�2��flj)?���c��V.�Y�R86�����u�}5zrT��c�\8�mpr�%� g�>��T�A;��bjo���fGF��&��=�B0
�9
Б�]k��w�$�_C�(ɏ���`�9%a����J��7qno�6F:��I�`<�:RE��PO􇂸�v�pq��*)��<�dw��C�F:�t��%�AF$����_񿘩Eʙ����B0�b{� �>?����_�Yp�+�!R�mc���Kz�u�� ��Dd46@5oj�[K�)��UH��m�/��⾄��9��f3�eL�N��v1o�G�;��B��*�dY�|�P�J��H�bv��>?d*_?.}�(�ʞu=C�z���%��ػ��?�K���fW�\T�����h�Rt��o��Q]=g�rl�HP�:C����z"���c��$^�<Ͽ�gޘ~'�5¬�T���E�7�_���R�%Gg洒� �~˩ Փ��P�o�(r䰴��e�kiE�� <��C�q���	��r苁}c(��g٩�� 7��E��1�4����Sd�Q�j^�p�#���e�68/�ۭ+];f�������!���ʅ��)Li����y-�?L1�`��Wo��z1�m���k��ױ3.�ǟe��F��u	�)?�C�����[7�f��"B����0�a�V��О����j��\�ă�j��o��3.銃�
���p�%�:��ۜm�_"A!q�l�"7�a�X�K"!Q��K�F�`��;X�4�w���F�F���1X/�����yV��q#���^fR�9��+f��7W���Q|- ���݆z�"b�c��H}���F;ҥ����'�������[r?����ic����^v���\n�qNq�u�`$NMkes���Iә;�M2F7���}�D�xl"#2vj�zt��0����c�Q [!;qWg[\��bpp�s��������N�(�M*���(i7���{��Hm��U(�ө�
G#��TD*�#yc}�0變ɜ�o��S
ǍP@��M�0� �X��{��Hr����g��ͭ�aӡ)�}Z�I���|�d��}%�.c�U�D�8"	�C�~U�,�?��ݟ��Bfgn�U�����;�"��y ��6����-�
O��/7ɛ�VUfE�ij6C�^K�]��|*�J%K�go��W�i�-�������Ȧ	JX�R���>� /�euu��(���.�����zZ�-�Kj�[�6���|��)q
�t
zj_����eQSA�����HTc�\�(8D��xح%>C�KM>2�'7�b'������6l]�Ɉ1WsX]�Աߦ6(�E��M�9!��1�x"��E: �7e��TO���<��&;��������
�\��?:2��'RD�HQ���
�>������#����?T��%>��'���������*������X�f����+�j �^ۀe:7��7>�y�찗˭�&{3w�ě}=�`��G 0�"6lC9�#��dZ����H͙*�g1�8��#�9�mg>SX�uCf�rU��r��RB� ��:���?�J��r����%�K̐%�v�A.Cv�Z�מ�~�'N&=�����QO2.]�5V��Ĩ��WP�%_�8�4�ƁW)*���3�[�w$����mR������^$�a�㳐���0��Y�i���{�"y�2����"О[f���ϩ����x���n!R�¶dկ��r)��K��>WH@
B��x�����e$m�f�,c>Ug�$�@�r*�z�B�"jWs[��۞�re�Gr���I���'ߵŬ���E^���o������$<�9W���;,�"�z��?�7#����n}U:�*�D��tUz�B�)�\�t�L�uc-	U	xC��˵��j
���ǖ���~��3�����-m"{�v�u�)b�"=�u�KKS����Їu���x6�V,cE��R�rNk�������6\�l3�%m`������#f�n86O@^&�2y�@m�+J������-�>~]H�)���s�n{�濇ab�9Rv͎��N��;�~E�Z��M�C�} �x����de@�QC�/���a3}7gy����1��s�!Z(� ����>�gSm97O��]��K\Qɓ��\G��I�שA�TʳO�X:i�#��%�t9���~t��m_b�0��9~Q����C���7ă��]#���'��(-i���ױ5�]���F�l�#w�'Fm���0`�΁`�dF'���E�ﴡ֝oڌ#��KI��5�K�I�`ɊBf�����1%-
�]34_HlKq�S}����˫}X$K:��"ç%'ۨy�y�Ҡ�2Od��n\);�<G�0��Z}eacm��ݑ�~�J�bt���l�)Q*+����HS�CȌ�hV+K�.�%M�b�^�d�1��I���<�&�|�'�F��H�|��i����	!�-'�Qr��d+S��Y�fl���j�-��[Ϡ�L�����V���Ҝ���~!�Ir��3$��s��f��1�}�%���]��.��x�I�)���3(������~.2`�W�&���I�Epw�Zc�5�,�nJ,���'�Y�NJ� �k�+��8H+�m+�^[��poo�+�U�t�~�38�?Y�[i�@��^���A��z��Dt��M�3b��G��wv�a����9�??����\m���a�T^��#g~�M�A��Yz���||��u���|W0��hy	ݷ���.Z��D���V*�É���w���쒷g8�\_6	-=�/E�&P����$��Ut�8F�6�ǖ�R=�!�R��ٹ�'ޕ�c��56�EUJu���g� t��҃Ə0)�9��� ��G���L?8�l��kvչ	�j4�=��7u�ս
��)ll�Kl�6'&�́��I�l���\��K������=9�J�|��z-P����Y�䱔W�N�]bYyǎ+3̲N�-�S�>�{��w<�[��/N)E�[�Sj�:��!sGfVx|`�nv5���ǎ�M��Tw��4�{�&���;���/N���� n��B`����5<S��~l��By*�KD%�(.Ur<E���H.�y�z�>�,��lE.�/�F��]���EF�
�,v����ͫ<j���|$�e���]w���ˌe��6��Pʗ+�	�{ %8��V���)���a��Fh��_�[���z�h`Zw�5.��X�Y�s�R"O�â]V(���q�&�=��pe�dX��Z�"��	��D�N4���,2Y�cy'd'��I�@ᣙ�	�DNg��	MJ�{<ޯ�5o:���>�����W 0��$o�J����	o��w�����ܭ*a�,����b�=ĪTi�'8�T�7�%:��- �����hJL�E4{�e0�T=�q?A�z����0)C�(+R�&#�������$����Y���`L��C6��1C;D�5�����D�l��Μ�B�,�R�Zg�����3+|m�����#�]p �Z�����Z�N���l��`Ѫ$�������B��lo��y �wE"�*9�����*����I��
"�@zf�oj�u���pC�Ź�V�)�d�V���h�)����\�j�0�m��/�4:P`}y~��.�G�+9�er�s��R�Ą�|���(9��,1s9������l�Ř�����ze���������֐�Ai�b(��Ѳ�"��#��Di��0�Yk�������D~;�Aq�����I3t0L�l��O[\`X��PZ{I��`zě�t4��4A��a���kXm�0*oW��R�vIoɥ��*��ی����E��� {�Զ�CY��)��N�m����#%c�T���$Ո��EB�;O΃L-�ǥ~��t��t�b�+˔�V@D������ӥ:�M:�2Ƽ�j75z���t/_C���*��VyiWH�� �G"\��7��z��ޭ홟)�dB���A��CT���L໊�)��CZ�k$r�ccnʁ5�b([��A���`*^�{��Q<�;v�F#ɴ��*���^����e�[��Mn
ɒj����N������)ޔ��w�4!
�}r$�d���+� �VS%�8�.K���&%��T���J�~��۽��_ϐ'�Q҂#�:g<j�N R��~���m�5i��0���X���G�^xEZ��R�:��_rs��C�*N��Z�?��<	5w~b��E�ᔎ�r�����=��V!)ϯ��^XF4��-pe#��t�|#�1���3!hI{�l6��>8M��Q�X��f���v��04XK0|�=Y"{��?�́�{�B3�t{^_*�Y���M��!��<#H��$_����3s�#�0㪶B'
���=��jP�a�	�>�Y�b/�Se�[S| �T����]G�n {�<��L:�"��D_8���[��+�x�X��Rq��>�l�d]j��~���*����?m�d3��9Z��h���?�v"�n�6I$s���'x{{*����@i��9J����'�+��w�m�w�oS��#� �n �M��Q,D�qꫩx����"�;�s��"��'��<%����aG�ш%/X����H�ޠ%����F׫�B��ԯ�	X���T�ʉE�Q� h "�����d9�>�ōe��KV�b�i�dv�[�,׭�����<�N��2�0�Z��l4��xöڒ��^Ss�:8��.�a&�M)�]z�����JK��Ru�z0�����r9���VN<�oFg朇)��Q���=b�뢂*�@[���=M0߰��v礆Ŗ��P��E������ohe�~��QcU*x�G���+У)Y�]��^�Q|�
�JC*���%�ջ�d��2��NG�A�6ڤ2���w>�o�l߿��(�;��!j�y��\�����T�
�	�K����bf��2ƴ��a�ʯL�_�J�����^�c2�j���a|%Kq�ذ���w�r��O��ޭ��	��)4��U,��� R����)̲�4t
��� ܾ*e�ܴs^����$S��ZY�޻|�G��B�Ɗ|Aa�~�b2��,3JS1�	�e�
�.�L�i���-����� �����M��g<���� �Ex��]�q3Շk��P���+ p��W9泂�P� ~~p�멉-�
����@q���5>P���F$���Zc�v�_S�P�>@]ح�O�D�L�D�� �]X �G_��@u����ȏ�hw�˒
L%��Mek���ke�A���s�V��>�W�0V|�w��>V�6R�H�6�(���X��V�VÓ��hڐ��6 pe�=
U^ ���?�t�P����T�P�9#X޵Û������ZbZ*�'������>�E[9&(H� �\���fS^`F�bb�jV4��u%l}v���;b���*�@	�<v4��ݝ"�kX�;����>=�U^y����.�~�K .'��L(k)@�.�e�T�����BU�AP��M6.ؤCȩ��zu���'�`Qr�P
��o�
���à�ٲ��}es�����?#6��8�ۡ�rY��E�zU�Tt�7$�8R���VT�r���鳦8��W�E;b)N��i�D=$� Э`u�e>�����D�N��Ǩӟ��o���r6�����~��9���+���`�s_�4�ܳ[���1��j'�<��.���uHpb�4-�Ba�H����S����:��
�g?�C`������$y+Z�|T���0����;�f&Sj��%���"W,���/ͭ��B[�'���\"�s�@af�<���qw_�����
�UM
�\.**x��#/Y1'�R���C���/�D�udT��=��ܱ�43�X�����J��b����t� |���?gl�(��H����j@�[���N�f*z<��c�;e	�h��_�$�7nܖ�ۡ�g�U���ww^���?x���&y��T!k9�3V~����e�?	�R��A�؇cJ�.����\�ܗdk��S,?�4<�9aߨDIX{0q; o1�q�1�Ă�x�YxWL%��$'?uI�����%ܦ��ҷ�P*P�}����m	��w���5~�\�3Pj H�#P! �|�\m�^E�U���,�.�^I'�vݗ�C�5_o�9&KA+k�2�b
/�^9�0J&�ǅ_�͏���77��un���D ~w��o���tB��/t��m�6J  �'��\���Y�<Q�E4���H�ۍz~��4)��9$Ei�-)7@����,덞0���&��g��&� �����Wy��������#��9��8�O��2E�����4�З8�T]gt
h���B_�N��*+�[T(�-B�%�,���>݀f�|�ۓѬ� ��e���I/x���h2{�p�}���],�y8�/�ʐ�gJQ�m�✵��e�_�*�:a��9��Ay�4�������c�����/s(�;���!�x��o`)�Ȫ�E�r�]�c���w?g�Ƚ��WP����7�W%vv��d�$�%0�x(���ӾoNm���������z�����T#N�M��4�m���Ŋ�M|U�"m]H�Z���s���hw �>�9��=T
�5�?ao�ߒ�d`���I>��Wõ�"���8UC�������2�����#�\-%\F�څ�˛8,��$}�Z|L�N�g��C�;�������8tb�a:UB*���/����xW�:�i�CP�$��7������ZH$��j��P�6�7�#�(��1�o�xn�E�(l�]r�l4gk�*@�>hWd��0L7`����=����ڂT�Þc��l���8���\"��}�3s����}���s��R��!�p5ڧ5V� *�;�Jtoշ/��~fF���Q�p,��ԖP��_�q�]���*	5��� ���)���@�sw�9�ic�y�����$B��8,I�=
��Tk���)���-�W⿦��34'��D�+�	�b�P#��ql���:35Yu�� �$��v`V*�b����'gu&���E2�Vjh���à`�&R)�_OK�#*だ����JXR��FWwWq��Dt�4�=��1��]x�#�WWV)���K.bFw `�m'=s�7Ɣ�%�A�n�I�	іI���.�9y�]tE@�г�nGf<�=�om��}h��\�������u{�G���� ԄW"��`G82��mF��(E�/����׆�w~�W��&ҙ��Q����o v��]�ҴQ!�"˖ǐ�:6��4��hޔJ��j���!�Y���Y���*o�����D�P~PVj��h���h���q�L��w�Y�AUt��ۥW��o޵�v�Z$X�BY+$*=h��)�VZ��^�f����K�GS����sX��(�A�~X^�$�Po���ܔ��+N���ȹ���vx����O\��ѝXd>f1�cb�1ɕVG��n^��nB�ȨRV�6S�	o�?�D����CAm0	>�_�^i^ߤ��(I���9�́�s�oSeUw�D�Y�4,`'��夸��)F�$����N��п$#�X��x�h��q�gyk���M�3�yC1�L�P�{9�П&n` `t_&�O	T�O��' ��|�b����E� "������/��݁]p�����:�p��tpK�Nh�P*����;h�o�+Jb�/S(g�T��%ʣc8�s��(��ޜm�*���"������fj��.ZA�,�r�v@V�qv:Q1bn,teZ���������4v[Ű}��|\�%���g�������rIIf�h����й�܃^�܏��#OuH72�[W���qo\iJP����l�ky0)Cn��!�t6kJ��~�V�q
P�N�iZk�ۿx��녃����g����U2甒� ]�=�7�Y��z^�\��[T1�_�b}��L0��r���x�Gj?��������=(u��Sè��uV���'�O�$���j�=�W�'/�َ�Ћ�<�톦��2��-�spv��<$��*�b�X�w*Dޝ�-�K\ǒpb��F59�-J������&����҃/��i�&�9V4�����F�uJn�b�۴���5��AT�����{����F��C5�T�rklE���ui��$�2�G�31Bh�N�5��֙m�#w�,gG�� ~d�W�X5�.��P��"<�P�e�@s��:�^+��G+9�"����3��[��
ڨ�B�0��Z�N@�c&s�_�4�T�Iq���g5a��z�_D�(��Q3#ھ��Y�%����/QA��/W��p�$��jDC�8GI� e�jʹ�`>��{�Danˎȳ�KB���K=�>ھ�LNp#�����>�D�|������K���nC2�?��ӹ�p�x���Dg�D��DW5�coM)Q�M��V���Q��p	�#�bR�
������fJN����m:�J���_�#/ �����r��2G����r��?��:���c�U#�/�l4g��M����.��42��1��%?�9�,9ԥ�b�;OI!NQ���^��/�o�+5�5�7�]���8�4VH���ƙX��lV�<�xlk��\�;��;0�?�Hi�s٭G���$��M���v�x��g�)�X)ǂ���B��V�����?���CWy���Jc6i8�d�<A������U�%�݇/{�C:6bs��6��S$ ��wHP�,�]���jzY;h�iQBT,����	,����)]Edn �zі��JS��l���A��Jۡ���3$�H1e�Z>@P��+B}�$��<�k�n���d���b,��[��D��������gǿ���`� ��U���	'�u��h?�69f���c���M�?g�������e� ѹ?~a�a��d�oB;h�)Q�}�M�+>�i�Tp��Li��l��~�-�(Lvyc>��i#��q�NM���ý���XW�G�_�V%|��F�6�;hm�z%�(n(yKxqk6��̼<��{� � �^�"�"�BJt�}(6�Mr+m��Cj�uc.;T#�1+@�buz5�%���i�˳x�q�`^�>j���8��4R��� NKA���<.�ч�%�<�wCy���Ġp�s���<�0���L�%j([�JM��G.̫�ꖚ�����D��>�@6��1e[��rv�W'�F��R*(�X� �ǋA��۾�cY��a!ӭx�!6�=�A�+O#(�CA��,�˭]��0}��2�孠T�gG��H�6�x��L�د�45).rB�`�)�0J\��J���>���LR�kF��d����G���
�����?�[&v�h��E�qr��[ťZ�Ų�N�1f<x��6��xRY	�\�F2E�Ӌ��a�(_�hz����]��0f����(4+P����:3E0�u�=S�u(�ڢqc�l'b+LG����W����8_���n�'��l{C��X,1Ra_�j�m�Y���}�R���4��1�?šr��{!}��7W�M Ő���--%.o7Qo�s��eΑu �0�Fx��M�(��o��1?V�S�c���䔷�c1�m;#o�Ÿ���\ ��PL���,��|d�a�����q��X^�&��(]���ͮ;���I�-ch�_��2����9R�8ئ\v83Ǒ�r]_����j���jZ%��OI�O���vB{6��!�꓏{�u���yj��%x"(�����`�Y�$���6��W�6�3��5�Q�$Ñ��E!�l�ڕ�i����~���K>b������d��6ck��[������WZ���M)+<⠹UN0p%�X�����EX�5���xῇ�C�YJL=�M:o��H!C��NL���l[����K��*N1M]
���+��߿�2(��RP>(fE�n�Nf+���j8�9˳�<ub�l�n���3�\-��������?��~�4��p��1���z}��-���<b~�/����sLd�k3(���_@��Um{w�<����
_��su�w��N��{�c����D;��s��zh���[��4怽k7'0�`б��s���<j堏���Oc�X�� �^k*���(
h�O�	�{�>�jh%�SnĞ#��k�5�����m�h�F�#�(F�ɨ�{�z^�e�`%?z������kѻ!�а>vD��i�!�.�C�BdU�<�\�K�FƬRMqh�xՉ�N���E�`�O	��G�(�n���rG�R�i�8���$���L��� 4��E���ayk7�Z=.f��	��I��*�ٿh|��!�e��o�R�k��䴛�	�D��"�LoVE��]�cy�W@����rh����m���m���v��;��ߴ"�����S�:J�P�M��Nc0L�ߚ�>��ɇ#lT�ڲ��)C�¦����P-�T-�r5B���xI����EiT����\���Yeł�q��^5�C^{|��US?a��/��<�r�2)3�RU�{m*7X�?cES�e�|u����ǽ�޴�~Ac�5ʳM9�\�[qoRw�X���V�6m�躍e-�t��^�<����N��f����,�&�.�XzH/f͟��Z.����gq�����@��p��X/��K���!���}�]���iFِ�����>ONz�w �� s�����F�I�2R���0^�54(��U�{Vɮ��sj͍��"�_}&�Q2�����ݷg�wPz������W�"�����h�������9~xڏ�t��K�~�V?�d��$)���rV����봄TK����%�b%��W��*x�Z/f@���p�]
����l-���M"v/-��m̚ʨ��
����s,�h-D�`�MHS�p����W��s���EQ�]���kt�g�����K�rN��F����k�-��߯�����||�fBG��3)Ps�:iR8�8��/>X�=�cMz��/��u(OG�췀�U�="��7=<+\`aU%}~2�)����;߁H}'�����^q|߰g)���(�3)W�iQ��P��kҷ������i5���@b��>s��qS̱��@�����L�?��V�,�X�"d�-}��Fܷ磵ı�џ ����.噢�S�#� �\�FGE�����"�#����/CnK_8�(]U�\��ku��L�q�T�%{�#f�lw`$<Au��j~�O����v�r�������������0��{�''�hV���Pۇ�|Z~o���s��-`��.�����q�u�q��Wts��Ӡ��/���[X�?eAG*f��Hx�5mĬ.z�R��h��&��5��kO��%L��)̄6#��U��Q`�8ζ9ARX�1޲���&��v��t��u\[f�s��k�+���Eb8�ǖ�[�4/�dpd�����[j�	)������G	(͔�bi��TP���Y�g�"�;"��o-cG��#��M�K�6.��"���>�$����)x��記l��/m�-��e�wN?��`O��?d�ns�eG~�T�܋���:Q[�g ������~�xE1?�3s �����U<c��qq�Gr! w��Н�	�J٬�u(��0�pz]6��g��8������A�l{�e;��C?�����*%�x�E� z�d����~?$����T��A���굛�ۖ?������SB��evޔ���P_��z�<�E��֥5p��{�A���%�dCo�d�����B�>�tt*ş�=A�-��6,sc�_R��|\�l/c��ٙ(CyQ��b+nd�-���~�vW0�P�h���,"��{�(�.Rjfo �l\�ٵ�d²�6�A��Iw�(��O�	��E}#�u#��_{���k�Qeuɬ|ȵ$/Q�?ۉ֭�Ƹ�ә�J� E�}��/j&�1V64�g�7�!�z������/�-�/F� z�ex�Z��*d�'iN�K���N_�]󩚜�S�Ϗ�T�\�4��� ������:�d����BG����b�cx�U^��8��}��W���5�{�z�9�=�ҾtO;���"�>���%�/\@k�$�����`,�
��@N�����n�&��0��a�/7|14�DF1`�
C0d��Ш�ȘI��aT�Q=`����fV��I��i��J����(�/��U~1'��ʣ�L{8SI�g¼�< �S��SFr6���P��R[^����ml����y,m�]����8ퟧ��P�[�~��6��w�Gl\0����턛WZb��y�M�]���/��6�Q'Ǎ����Q�F�9�/:��,߇��<��<����H6�:�@Fju�O~��A_�缴C�V'(HtMv���E�AY �SU�1�}��\bZ~U3L��a@���R/�y�%ޝ������T��/W�t�� �j��}�ܰ���5�/��	t�nRU�;�2�;�ܦ��w)�4&�Cύ�΁r]�C�`�ق��i"�+������x���br�:�5�p��}���r�2���d��t+�4a����H�EUl�RX���W��P��pUb�n%d3ˆ����}P�w��"!I�e��ឪ^X��Ѓ?����9��!�U��C�P�U��RM�Ѕ�@���zc瓯iK���ȡ%z�̇�������x0�M��*I	2V}��A���Q��ёf��tR~�K%�/���|�A�Ѯ�H��m�!�1�GC��q:l�乺#�Bt��z�Z�e!хc��k=�b83ȏ����_U#����b��"z1��cA�@��>��"v� ��F�e>{���c�sI�<@�B̳L�w����/��!�uq)�3_�;�.x<�|�LϟE��H��8�_��x\��OL>O=@:�$�����?_��E��QKv���r��z�r|Z��^�?n�9�of��A���rT����t��z�'��6�&齴$�h���ɐm�����K�̘Tk��jX��Z�0��<��My�L�_*�=�"�v�n��Y;����(27[HM�գNQg=ra�k����ו�^��.�0u�aKt��"��w�Q�OMm����T�2u�����
�S�1k$)�|�O8ߍ����&5à�U!(�A�o>hә �-�����HҼg{�ˌ����Y�ٴP�
4� 4A#�)i�E�I�w�L~�+��µ;��5�cB��r��E��x����(ف��n�஡�e~�B�N�� �`���q�v刢!��E�O&�#݆1;"b/��PպdV?r_vb��*���-D_݆�"n�Cf�M�N��$~�ʍktȋ	@��p��|E��Og&s����c��H�ۀ���y���c�+�º�.$��ƮC����P�[w>�3��@5���٘Y4a�*����#����m4��`�E6DI�[M��HE����<���o����[waŒ�����đ���Gf�YO���E5�ӷ���%Rx����} 0�>����ǝ���P�ݎ&��.���.=�l��� ���֕G�ƎF�2K��sH����Rb
���;���x�S��BZNV!�on@vbU�!�(��V�"jɓQ�	|�$��ds�ٕZ�WQ��^n��Gp;��+�'$�y��K���:J�>5�ͬ��V�G��O�����ْ}�aQؼ����U��m�7�]�W���S��XvL����]�t�,Dk8����8N�
�����Dv��ݷc]0�	:��-%֍��W������7����u6�C�T������Qʏ��_*gp1�_��;r��"����F���J}���D ��IOL���p��"U�,IS�  X@FX$�D��?{t�^�J+������D���ʈ�:ʯ��i1XF��rY�^��ks�I�08���<�~�3U۪�9���I�<8��pܻ�m2������/�N��sE���RHDw'��2q��)�{�G�P�F��G��l�}��9���v�nƦu�!>�n����sos�?â������$�7�d o� �{`	f�Z�,k㻃�%I�kL�6�%1Ձjn�7���=y��àل�X�D,D�Ǫ�ڟçfo�����j�VϿ��)��w7�CjԷ�BmG�A:�DR��JK1����֑E/P����R���v$ܗ�Iը�wʥ����l�l]�afQ�Ru��\V�E��eq|L�E����Թ|�T��7䒤�~7��{A���#��H7�<W��K6W�j�H��D�$��:�����W!{��O9��\K���D���j�����$�"y?B9�X�����#x`ۏ��>G'�Su�|{j��9Wl���L��9 ���s�vb������:~	3�=��-����Y�@o�2��INGʕ�̋&Pb��H��ª��WSG����Ð�a]��l;����(�+NZ<��v+�Z����Er*���P��.j�h�>�r�3O��h�m�}��FX�Z�w|�l�Ϯ����Fb^�>l}~	K�ˤ,��0O	{�D��TL�r�FEF�^���r��;*�6+��� ��jV)@�����?zA�%tưk�6�DZ%�Nq���������k;�$���=�ڐ)-�G�#-,���G�YE��؍�����Xo��u�#���~��X�Բ��t/�oQNg 8��~�}��W�J�X�G�ɘ�W�q�{�^�)�15>�׀*�i��I$�>�v'�b������aBf��*�m��IT��C�.��k�n��-�4e?*�������%��s֍Í���M�r�X�2띩�����r���5X�a�����5Z�G�b�Џ࿰�k������;9�W�`A��'�;N�ޞCP�v���7��X�CΎ�z�i��R}����r��o)e)}8]����m��$�H�#�= ��ȭE�H1X��q���kv�?e��9�5�R�>�8m��X��nT�^� 7n���{\��Ȥx=�Ǭb�t� 5b�g�_bVA�X儚)6k��t]F�Z�ϑA��ٷ��HL�Y�dW1n�WN�=�T��А�e�gwr�k��z�=fC&k+�۫����VD���p
���9�M\>OYՋ�,�jn�o��M�%%C��͜O9q'e�ny�2ե���%A� ~閽N�5�D2?[��_������nŒO ��bx�d�4�ҝȗ-�Gʄ�{$�[���pP� ��hb�{���I��	�+�h�=������]��i_����@j�y�J���)jJ
�_�(#���o3��c��u�<�b.�!�C,��ؠJ�獇C�-yw(�J�i5}7]m9�"���n<�-,�M]��9^�r�����Ǆ�z����vŁHv���K�P�HҎ�XWLG�1���-��7��$�*�H�F@����������I{�W��ZC��� V� D�4���./��!�8Σ�1��`4L��(����(;3�Y�wm���ߧ��L�N+g
��b��3�&\�,�ћ@t�G4���6$��x�c�~�a�}KG�q�ą��_F�9=�����;,�B9��;f�x�ԗb���[#�0�%h�/�������&��C|����o���E��>�̫�	^�A	�@0:}T��&���z1�H
������ߘ�E��['q�~���U�.�a�Q�� ]	�\T��*qI������ds�^NL��{�J�������3�p��w.p��^�U�H�ъ9��� �܏G�Z�n�7	����Zi��סX�b^l���V�3d���f���j���xff���#��,浥��>(y�b�M���^QE�2ݧ�"(ڮ����d���L�I���79�"�a�0H�kt%��a�UBL�yW��I-MY�'��E�`s�Lf���m��^H�ɝ�{`e�&s���G8����#�=����S	�*��Ѷ/i�e��U�؞ذ�K]~�xS��J���x0X$�z�(��1q���A��"B,pK��ԗr��<f���I������S��d�hN�T9KZ)���&M~�~4#@��2IQ*Aޓiض����6`
� J����,��& ��1� Xͨ�]���:�f	՗�֓y��1p��з��gt����"θ�"����0��*�?\9��;g�I��*��B=a��^̩�6<W�3;���F.8N�S�K���H� �ͫ�pS]����#���M^��Ћ�I5%� 	<�����ymoA:q�H�i�u�Y�h�i�4�l���Pzw�P������[�W��5yZqk��k�T�
?�>&ʥ��ٝn�jI'��]b��l�ڪ*�is�l��v�c��.��mn7�����ո�
�~�tM�v�ǵ|K}^�(��`�]�(6�Ƃ��J�ysF�U+��c��5�,��@�X8%~w���M#��V��# -4�R�E�ri_��]�.�#�v�3vE?x������̀�-��P�Ñ�cހHk�Ӈ� ��ň���r�Y�R7_՗U��!\fp��	�yto~4�(�
��C�d�!ySԭ�C�D#�9��+X�X�R��=���A����?+H���磒?j�o���D㥪	*PI 8��I��IG�ԅgM��������n�\���*�fܠc��:$�O�22���]ۋ�����]c(��T��Q� �����ל�G��~��<�z��*�r�^�X�3sg���s�)ň��K�e*߿�ȚH�y�o(/�=67�Z[��,���g:�cH�8`�b���.�܈č1YQ�a�ᒯ�����S�݉���Xa�=E¦��&_� ���A�"�7Scd�6�>>R�}t�&ؿ܈�
�Ĭ�����*͐��K�9����9��3��U�
�v���	%׸�:�D��=Pj~��l�׳�_K�f&�}Tyۮ��?��y�����.�Ay�;8�[b��S�`0S�dH�D��C(���� �杦BT+��An��1�0�����	����6��֭���T��)P���}di�;Z��!�������O����d��{<qpU�̷'�=�T�\�4��;\��}�s���B��)��K"��q&RF�0��GV0�Tuь{x�^��;ޯ	��l����8��s���y����(p�PiA3�;���enka �T�f�K)�+}��:����@�4uy�x��&� �+�J�oʼ��޻��%V�s����d��mfӑyٕ`��:��0w'c����|�RXH%X�$�C%�HK|��N����>g^C��5u������K
Ew���B�':�+��(��|�]�e��E:��Ǫ�w5�4\BMw��� ����U��TzqzS�^��f�-��7Wc�ف�5~m�Sݺ�k1����M6*Q�a�ղ���$pb��}���3�Wz9~%.VF���| ޱMrOx��,��tB��vC�b%�y���C�M8��%wr���_���[��|)'�5�т�;g#���2��>ݷ$�~��_�U�až���h�	v��g�\�V�:��J	��#��Ng�f�%�N��l�3f3��Op�	�_+�T���Am�M�u���/�p+�*O[TA���]J@�a�w��=��Vog8�f�������u�.lm8Bt*��YגRGCᚊ��x0�Z�<B�@L߶r�:�h���Y]�N)��n��Mv�b� ķ|Y	U�Lz���f��,o䚡�ƫ���Kp���wF�.�~��i����l約�lp�EG�I�	��
ʎ-2Ӏ�$&2����(@T�<��q��6��9R�Q~(D�uc��F����J��^5�@�ʜ�ES몼�&A�(�P�G�-A�C�?�	��n�}	>�P�R������+VH��{9��W&1�+&�H�^��B8�X�"TU)��#��Kb�*�4���zēo�/b"���N�����s�� d�M�����s	S�V�J���N�"J�W��?,���ݒ��1��JU���G�8Hy+{���L��S�1�,��@�}8��_��/q��~!�������oy���
ߚԵ�A�W)^�#ã��X�p<\�5��U0N�������q4	'9�PI\vLp�q�O8�| ��<2�z�4y���d�}�~�[!0�����W[��h&k����[�K�,���,���}�z�@�Ac�M�C�̜t�	�Ɖ����C���$l����� )
z�S���� #�X�5���}_�1�y�hƵǳ�Ԝ(ow�=��q�
OrP���h� �YhgI�~Rӣ[2�ǿ�p��hx��gp������L�қ��:��ԒD'(�=q�և�9��WD����#0~?p5�����i�Q\�ɰ�U�/����?f�wka�2eg�վ��tO��{�QJ�޳S"�IN�'-=@ۊ�x��"-�s�c���3��KU��>m��g��-�e>�����]�?J:;%�	҉9X��,�g`������7	 Jgz�^hs�����!�x���i�O5���E^5�+�# �0�L��n �I������F8O�@dȑat�ٯ���P�q��Z����<����d��b��W7�w�nʆ�?za�(�}P����|8sQar}��9�d����<X�� �ĉs�=��c���h���Fx-ް�����a8ҁ�j�W��iN�,�n8n�����L՝^���=��u�=��H��p4�D{���b�x�����O����HX�Usa��l�h��qaiM3����@"��m��@�8gU�3nQ{��U2�ΩB����ET{��&Ao�
.��g��#S�\J��
Q~��D&�;cuJi�4�	T�^�������؇����R|K���yև�5̻����ݲ酧�IYR��a0�<C12�5ߥ�l-%��Yp�8������+�^ֶe�r7Tsܫ~�/�
C<��B�Xrr|�E����ٸ5/��g����]	/^E��1��5�JP+f#�\I��`�e�+����F�Kiz�l��a+TY|pQ�k�+��-���+�b��V�28�Q9���~�澟\|����}6� /��#2��v�/œM5�^�W���ӻx�Ken(�8Ei1{D R�9�!<�pam{�ƞ�W[
ٕ(��We#�ycU��B`������'8�3��eD�(9��� ��ɒ����$�M�g^nl��@��<lo1j�S�7³!o{�l�ʵ'�T�SR�{<������c&��O�"ða[��NO`�l/4Xo}=��Z�@�y���.!,�y��^/��C|ݓkpa��3��#K�2�?p4�eg��g���@)�}[���͋�e���M��o���&1X]0�k� ^�Fa�\ F�&Y�#�iUM8��4�|�2�ae �e��9�?�iɭQm������b�k5MC���`oNp���ܥ0��F�g����W��Z�>ɸ@�{��7jɊ����<�2 K��o�x�|���������X�k���)�\7})u�p~T)�Nq�c��t,̻��T�����	?�b*T��>���09�0��d���K�V}���KS���=��	/vou����]<ca ��6�CT��ZMC�:��&K:�~R$A�~?��5�q���&��qZj�ў�jo&�l�Jd)nV.cP���g�FG�����+��E�Ʌ�J�U9��0_��C+����=�7��s���t�=��@�6�3�%o@J#��PdJΖd���而zQ�׃�ɟ�{����*�<���!��8;D�K�)->�Sb(5��g[Ar�]8�+L�(��ܯ��,�;���%S������^;�w�Y�}�Y���؂�@�Ҝ�#8�k���v<�ѯ��A�y����(�6�Sx8�i!�|R�`����^�!P��z߲�X���U*!C�:B���9Vҏ$]�i
rnh�����*��JK�J5+��ɖYy�Zxk 0{�2�`��u++�!Le��b��]�N7���I��$��Z�o��	�C!��T��O���6�4��[�ڶg=!`�y�g�#ޙ�XdNL�&u�R�!�&J5!��"�o}����e� PRO�*m/%�Nqt��	���ݬ.s<��O�>�غ��Q��0/u���-�Q�DFDM��A��:B4�S~M�څ�~fn�}į|�2t�T9�(A~�n*�(]7��<�xw�7���tkeB��X��B0o!�æ���ANoƛ��@����Ɍ��ҟ�'����B�U�C�:ʡa��rnc��p`Dvm�V��h��o
�Z���b��ig+_�])�[X��&_X)Q��;�����x(}�����ˌ�v1��u��Jbh�Yng�(%O'�v��k�V��r�6h_@���i~��>HI�un]�$�lD?	�~����aƑp�͑'�E�U
G&�ȯ�hqm�-� .Ԣ��=Fe�!X����}a ?��jI�zvsv�d�b!||p��}�U�d���DC|��H���Q/�n������\&��?u/����B��Ö$F�	:��~e�Pf�J�s?��llU���3�o�~������'	���[ݮƠla�N��e��B&�O/)��i����[���"�{5#{��3���`c�]i8�����ȕ��{��}�ܳ֕��q�Ś�ukv��N���7!낾�_G
���e܀`*t%�~�d����Q�x���A�W�-�t�o��^�zx�G>_�����Do}�3��P��^iw�����s�I�i_U�'Cx��lC4�U]R�;��"c���o��\,�(HC����a���N����%71B�'���h�nb��3_��]���P7��$�a�"w�'fp�:�Do����[�K��)�j����O.���Fih�S��cM��y3�EA�v�翚`>���\��!�4BaJAa;B9m��J�ֽ\fj��_��3����z5A����y��8�����.#�mȉ���H���O�$���m�XD���!��*[ /����>cK�Q[�M?{C7��0��mi��5'g�ڷ
ӑ2� :�拲��/ ��RgG�s5M���as�`����Ah(t򈀛ٜ>Z�Bm)�sX��ܘ��5����@Dt#W�j�F��ϼ�c�
WSg��vK}�n��܀shq���ӡ�CΎ�οي���� ���L-�b�@�)��|���r!�"���k�T�5w+�[?9X#���/z���� ��.������,�e����z���۽TCde�>��Y[m �*�'������G���6i�q>��U
�i�+�77�E�*�^�@���� 9}n����)|*c�#.�@�	����<���p8Į0�!B�"<x���T*�d}w�4N�����Δ注��D��Z�5u���7��Q޴�q�R?$f�;�0��h�K6� r�/�WB��`����^��~�|�(�EH�Ay�>dO1.��� uLo�%U�,DNrھM2|XET� W;'��cV�C��'D:.�x����G	Ou�>�a΂>v򣢇r����Ý�H;��j�R���Ξ�唤��s�f)N�i<#Nh�g�5X��N��u�-�}"���2;Uw'����,��}�'�G��h�#���mU��~.�X�
z�7����\�ق�ީ�_m���}�'�mC7Z�4�k����X�3�����L�0�=P�����f�/7h1Bx"5�e�8n����L>�P޻Ԧ�����$��w۫��B��]��®�a ��ڗL֞AZj/��%�������0� a-����:�0�Zb]L�.� d��1lV�M�$B�Ä�\Gx!-�6J�6Ua�k��!A^s�-/����\�Qs�Ys9g8�:+�*k��jc[p�WIby��8t }{ڜ,!|cg��V�LdO�.X����+6+�B�z�������.�G`q-T����%oȑ3��'��5�Tlvq���ă��5|�@y*��:g��i�w��^l�� �O)��l���ص�>L�M�~)�;?}Հ���=3=*�Y~KXe)��B��8,X�洵E��gm�1�~i�%X�$K����_#�J񛺰}���(�R1����
:u���w��P�����y�&�}��'2"UuN���,���r�s�HHx[�ZYҿ! ��r��j����F8�^ucޯyQ���~�ٔ"�xEX�߼v���I���!�26 �#��
;��jh``��a��M���m��`J{�+��vܳ.V=+��xu�A'�id��]� 8I�l��{��*S�5�fe�*�2cz�l�3�&ss6�� 	V��T���k]�æI�"���+���g�o$9U0l�>�xxL�٭0����3$��>2�}�W���x�1Պ
"�.���q���>8����������q�EƯ>�o�K1�>O�����/ƚ�F?��r�@2�&|:a�b��H�}&�7���hv�0���x��@W�� ��Yi�=���
�sR\Ɨ�P\�h��3�5,'��Gʹ -�5�����ϥ �H('���z���0�:�F��t/;�C9�����	8+4j�]�t��0�#A&�A>�����vqJ��n2��x�T��M��5G2�^����v$P�Orb `|X�\'(���Qմ?��p�:W�9dk�,�m-�@-�
���:��7�_�on��q���^�,7\��?�~g$�����B�:�I����o�;l���F����n9��*���|�l���}���Q뾀|㖻B��]�4�SU��Gk�|c1�����R�H@�PF��R�����u�Hm����6c�[��mӘ�L�����ކ�����z���\rx�3l��:o�j���-*{���*/�,ʨj�J0�SgęF�ȇ+��9n��4�V�\���8�|,w�s$�L��gf��RL�W@PG�='gn��M�B=ߙ����r]���_˦]��\��@q� ��X������փH~��`�=�;E%��i�ƕxcV��>�O�v4��M��R�B��>AT���?����T�No�2a�|���<�F��݉	8?�-�-�Z��ew7��>����E��c�CEؕ�O�N������9@�z|�"�������5H�_�9��4��ϛ|E�j��ww���G@o���Y!�+���%%3��>n=T;���/��[�6�� �:�(ӣ�����*p�=��1�ňx3�t��c������R+7\49�E����lKx>�T���������`�]�������Y�Q�b �;-��w��0H�Wd�v��?b��%m�i����8��Uo��0`�xˬ���O�&G��λ�"������r`����>�gg�'~I���9s��MB����۠�h�s�v�dg<c;wU��p��H��FQ�bϻ�>�ٓ��U�>�wOL[z
RY��fu�
j�����F��1�g:Cҹl,�=|���.E��*z��DyY�����B7K�x���+�j��qXL�+����
���� �ϻEe%K1	�,�:~��2� ׄ�*Q�LG"��^�ȓ��Pz��!�����F��^	_0�_���'s̞W��AWQav��EU�?[����W����tl����Ov��������u.ͭ�������V!4BUbz�Q�rV|�~_0Gi��/G��߯�K� XCJ��'���R��$�A����Rpm�<V�\��
c�V�V�U?踏l;;/D���qv,v�t�{c���͔�����N
��}ܫ�)K�K��K����׵E@r�����2�w�+c�ouƊy�c4j�q@\TaUߨ�ǝ����}��m�p�v��F`���8�X�؇���Α�j4�åqn{�:�w�5��ƭG � +�)���.Nl͋�x�
�)��{�,���kb���p���:���`6ine�ڋ˰�,����J�<
�7Ȋ �$6�¾;Ⱦ�D����P��H'[�=[���Qx$����|� ۞R�dc�z�p�Ac<rK+;2\���	a�~"#��O֏�(A�b���ؔj�wTKSP�ì*3��3b� ��,i���e���Pe_!Ё�/��a����}M��V ��~� 5&�V����Y�t�[��p�;�,����_L��ѳ�4#؞@еM]�	�"���v� �_��w�8S�ԩ��35�y���.Z�111����<W4v��p���5@[u���_b��k����"�ɶ"��������Ʈ�k��/��Sѐ�&C��Y@���7�ӉQ�I�w��0R�(���ɩ�~x7
>�,U�4�UЯ�A@�����t��U�%�gPڂ4&	��Q�2����0��B����RW�w��jËa�'	���J�ƀg��� � L׭;����p�ϽKgXk�&�ĺ��]~}�Y~�O>��K���f�]yG���ג%+�"�V�b�M�J{�&˗+<wW �ϭN.�U�R*��(a�)q.\O������"�������D)��;S7)�c
@_@b�[�*x�S�Ҁ\z)�sz�����cg&�qZ��f~"�i�cz��"�E��m"~�oauA�vi�ྼ�8��6Zײ,�6`Mn�*���iGy��VF-΃��y��)�Z�����e ��ҁ;�5vL�h���;����E-�8��0���}y�� :����'�[_8.hj<a;�Rwٕxի^Fg3oTu�
non��qp(�7���E�xڍ� TE٧��^C,�4_�VT��8|�3/t�96�I�ù����b�X�^V��Tx��?+׮b�Aq7:�t��e�`�l$�Z�o�tp6�j�Q^��?�4�w��ߑ�j{P7��nTru	����
Zӓf��������m� ��&�y�I&�K
 ��+���n���E>�(��o��K9����^�/��%"ٟ$����+�0�����-�C,izm!���2:�K/�;��b@�b^��?��(�Ap�*@.5ɇX����;�Z�,� ����"�Fޒ��+��u�=�^��9'��� M�f2(H!��)KiQ�J�{ ���� �H�k���'N�{��rA�|�I��,��\�d��g��$�CD�N݁����Ii��p剐0]z#�B�}��^s�IZN]Q�
�^�~g�y{VRI�4��N���}�s(/�6V������޾���\q������lY�r�.�q�z������R+��\Z���H�����*����q48\f�&yb�.1�Ӆ�9�,>����c+Rq�B���c�$w��b�g����	�o����n�9:�ʠp�"�M��8�?u�+İ[��`jc8츎�xpXŌ�������E�o���g�k�H���g�B�U�Q�A�`� ��鏤NJ�8��&YsH�^r'XPz�5�Kq��!���%: (g�6*����F�'$�E���q��Kw��j��|t���P�bx�ՉjDr�\S���p7�K";J0���&�#'B��4Jѫ��v]��M�����d8�W$Zӂ6Z8�*�Z�F�}��==���5��Z�EB9�[>(�n����q��khD�����[cXӼ-VEE���Z��N'	�� ���y��xا �u��u�@v�2($����/d��[~<؛����h?~,��,_o�Q����NaM���U?�ݯ�?	�4�,�6@(o�]Yy/�A�|Mi��:�>��N,�p"�������,@��l�Ѻf������ VZ�:�Eӽ-�]�;�a���ٹ�3q����m<yO�g�qD��!��������<�!eY�����]�\��;�m��ӌ��$�;E�B^���{O�
!�T���>�N?S�n��{T¨�4���"��g/	�����'�.�'Є��J�W���B��>���$���3 5z��WN����E�ap ���TK��;������bo�\��g^�_L��{���q92+W�ģ(�]�}=z�b�GBk�N�������b{wt��'�6�(
�Y�۹���#�u=�$`_� ��l��?~���#o����<��Dr��a�B���+Kp}������@N��w���牃���KZ 1��	���m�Ǭ�>��@+��q_��Q���u˚�O����&�s\F�����e&2�7�.!�16 �\T�^�v?℺R���c����M�~��@��2�����ߛl���#��r=�9�� �Q!�:��y�W�K��cO3��w�r0}/S�oӬ���-�$ch�{+)�`�L���(p 2��֪�q���7�%��ը�H�;DL�lty���	�H�ν��mۇ�@/s��*7���b*DX}�1抟e�0}���m����U%)/P��8��U�֗�������a��>L�ݺj�bD��lk���&��l)2t�\|U�Gu�eWw]�I��.@���Pu��9�@�6��2QS�+��?�!N������2>`�b��m]��р��1�Qøa�����&������Ѐ�ͽ�'Jq�k�+�'�rA*��÷R�L�\fW? �奍�k�p\�3Tx�߱�	���N�1x2�\���dj��9sRH��/VHv��u7o�U���u'�O��k
�n��k2>7KY���g!t�oE�4��֋���E��-�{��F����gS���q��ҏ ���juuVn�8v��"��H�WZ�J6�i���� ���$e1������%��3�̉$k��������|wάfla��:}�,G5d˜�ɒh�Z��C7�m�<��(oY���`�dr���S���A�v�Q�ZКՖ`��	�Z��Tl��P�8�z���.6��Y�f˂)4�F�N+�/D�.-�CD���kHA(�������p�X��"��f��L��*M���$ټ��G���ZS�!�8�ƕ���X
���'���INb��`*JBBG�}�:#�Sh(�xwH��%��/x�=�9Z0��1�Vۉ����E�K��Ƶ�,x�gV� Qi�P]o}�bsq�C¾=~lC�
�ԙ��}��� �w�T!�5��=R��>:�P%3�d�bB�qP��u�&�D>��&2N���z'3����DL��U�t� �����	M���SA�!�[
��%
ٖqԗ��VSQ�BJ��>��+������3�/��D�lFꪠmw����>~+�4�%�8h��(K���� ;��p��|���N�Y�����'l��E����&��2�E�U���D���#����N�G<V��VdKshަW�ǪS�y��w	\�Թ���,�0)#�UA�"����Ӷ?
����ú���,�?��a'O�r�i/8�� 1�Z�TRK���Ռ0&@�|=�%?��(��sQ]�Oܟ���Z����̳a/��:�B��hL��W
�]��g&e��Vg�]�4CQta6tRtw�e�.�3�-��A2��`׻����q���cS>(7'��P����w����g:1u�.���v2	9��H����Ž���|��A�F����$o�A��|�-�	�����d8���w�S�v�#��$h
D?��Lao�I�M8�!�PG��X��2�`Y�A�(G��Q�-J�M��D�	�ud���	1�����Ax���q�g9k��C9'߾M9�~��-ɐrwQ~�	�F��5M.�ک������3�X��/�T.z_%�U�M���������;�ѷ�9I���3l\���$����
��j�I]�*��QO�	n
�
3���H�J�&�8�	�-��Y��2r����fE���RQy|+X��� 4=��x�<��sm�D��@ߨQO�	 �4��
���R�����f!��k�$̓�O���t���V?�]���I/�?M���P�&����3߶��]�b�� �����[�]��}����TK碙I����N�J���+��3�fQ^~�|��q�F���B����*W�|
cI��gw̬�6E�Q����B�+\;�7|�ڽ'oL��'x�o�ȅmw��D v���R����r��Sa��8��V9�έ�$?)rA�Fn�I���o���3	@���%��V����5fl�7�F�5��Gn�e�a0�Ώ'�A7<�Gq+����	g�����"����wp}����PV��?3xf��((��mZ���L{���o7(�*�I�G	=�Y��B�t���͍Ka�o��:��&�*IS�Yc/�Y+z���Gl��XWΉ�њ"	%�)نpLntK�}�c:g����Z*k��yk®̌���y�QR�ɳor�����#����˿��}��5�1V������1Ov9��P�	���8>{dCF�JK��~��)`�0�f�.�
�	 �� �����$^�ip�,��{�b����ټQl���w����d�^�_��J(�~v�΅�ڎH�:Ѷ@ ��̸��,����8L����� J���>��x`3<�튊c:�p�Yۄ	t)��rg@�������Ҷ�M�+��C4�����@�52.�N�ߏ�WX�:���F��W�҉������s��rI�T��\F#���<#�����_��^��{��Gu�̝ـ����@w��)�#��<������i��Fa�To�O5|"��Ca�����,,:Aό��f{o� Jf\l�����I�"~�p ��Ɂ/�3^�1[��e�d낁�Ra��xxЋ�Y�Ez�d�'\D���l,ϕw��
��s�����~?�T1���جoΧ�ǉx����Djkz M�n:x7��RG.���~��ؾ����s���փ�btߨ�`s�P�#�6IDp[��C�]X�'0��H���+�d�W!@���##�C,���~6a�����Z=E9��,�~����f<�Ħr�(۶~F��ڗ-�2b���-s����ˊ=9�kkk��W-ĀQO~�˖�U����Ml��qpFn�W�\��AK������	I^��v�D��[���ʥ�˛�D"�Z���6�hܷ�ˑ&*@��G����y���AM|Ґc�\r	�m�%t����������lr���y.Wq���C��V$*��AI�	�D7t���œ�
n	���:2� S%���g��F�d-S�ޥ�l*n��UrrE����`�����D�\�yV�g0�e_��D+x}/����B /2k�m��1����}��͐d�ˌ��i�	�q�H�Z��q9�����f�\*2���iv�v���]NL��l����1��2 l���jU^���
a��OKG��.�	ԕ<�	u���'�ԏE���8�/!Mo�̻MA���߭�jp��s~LK� �J?��������ɳ�^qa5�R+�S��k!����tc���;\L��fe���!T1.�9D-0�/-�������]ݯ�}J`���׍ �/�Ƴi@�P�H��MM��|��1,��}��Эvg~�P(�JRj[�ac%V�N��^}�U����2�k]X��O�NW4�J��p�S��Ҥ�,����;�4�� �*51�=�cE��[h��8k�L� z"!�6�`�hd�Ju��a'��}>i�C:�O�rU�si�%|��G�\�?�8Y�˾���Elb� �FjqR{:�����ܜ���W�}Kg���z��ؿ������)�[/!��u��(�涠�s5i�d؊�����o#;f�K��T���ۅ��`���_C�lƢ��M�W�#�~@�Us�c�������s�(�T�_V�i4��"����}%��Zf JR���w��6ݷ/����H��x�'\,��tS��:�0�����A�o�0<3s�(f�ʡ���.}NαY�{���&�P��8��J�<`�}���'�Bǅ����M0�{[x*D��A�x��Xz�X[�����(Ӵ��h�Ƹ��������w��g�/��Y�����~�lWQ�tD��W�cﯼ�ٚ��s+o�s� �%��Y����3r�ةG�R�㪧ㇲ�%��y��P��͖�Q'��1�Q��c,+nf��OuD�*P��MF��3�����A���l⏠�F�UTNqE��c�u[}���M:�/�(���L��n�_Qc�'�)}����!�-]�k�AP���M����|�`��W=�ó�r5�a����?�%���-(c�2���1p�����:�NF/+�nG5?�3��J[����h����J�.��g
�P	��9���٦����4p�0e�������y����u?!?�1�P���2��`�9\ƣ�n�3�.|M�������v����Zo7�;جņ����j��a�
^��o����G5�%���Go�o���U�Ҽ�AF%��Qo&9�bdֱn������FV'�&�a�M��\i�����%�A�f�`[6��c��F�w��9A��'�Br
Gb11�J;x�0y��.�k�M/w�v����H>+Zxru5�9�g����ha���9Udg��iL\��./����vq��]�{;���H�v�����.����K|�ґ&Me�yY�k@zt�;�ʸ�/~K�;B;g�pz�Jz,͈��"�!ۺ�F���	�k�h�A�U�p��Q3����pj��pAH�5o#�"�9�	�XL���m�=�[���3
$o3K@×�Q�R۶���]b�-?k��9.	"�m� �s9e��ˀ�����k�@���y�H�/ѨF�~Gtg���Q^ks�T�����i۠y]}�p�Z8ۆ^te ���Ҡ|\�x�/�2}�<���n�w�x��۴��WO�d�{v�y��DEߨ�r��t���f��j�0Ʀ�Mqf�����/�\�d���r���i�]�PҸ
X�tq��myaWF�of�ݛ�w���d��8:�a�s���܇,��C,3�=S�V�A��P��)&�h��<"؞�Q���VJ�i��l�D�����M@���8�U��hp[ 5�g!���@���k����VN��@zD��'4GSF:����ϰ,N���ݢ �ZNe��r�Y�ס�F/6`��W_���$i�'�у�y߃	5o Myq(�RIr-Â�[rCuF��7+�PFS�CX����;":��h���}"h��@�%"�U�<��d��I7��{�-k��_��]�#�-����-��	�<�y!�1�)���%�IWW�'>E��S�h {�c�D
txl3�t��B�T�V�e�5r$sݥ���Dv�{ё�W(.��U�q���v�(�1N_yJ��]	c]b�Q$|�l�ƧP`��26��z��fY�ㄟ/�6���f�K�[�����D�����?lMO��/_�֘Z�i%�����*��֌Rܖ�=���1�10��'g6O�����D����1�GDz�+FM�
6��$5�v,9f�tT3��XAW%S��]�����e�6����'��7�`���9"~�⨂p\f�gRV�2Bčoc��[N�<d����Yf$��u gh�� Q��\jA������CC���#�H	T��[�VMQ"�~��Ľ�`׶p����FF^4jA���3��rz1��4��M�D��dId����<?�����f}�xa�� H���{QPU�����Ve�}X\�.>���.�|[c*�i��3��5n����fCx1^&�� 5J��⯧�~��њ��E��ԕ|��л�괅�<��,|\T�35~��Y�~�,ϰ鍦��G�#�|O"���H0E�Q+�ǝ�z"Z��h$���u���z2�U���i�����(Z
R�駜�<��`շƽj�J�����'��%s:�9)��I��k\����ÏPa;�A����F,别�:���`լ��T��*���c@�X��Y҇�:�ܡ�:�^�1W�u.#�����h>w�b����
W���y��	�I���\z����2�F/T�q�M�3��oj5�~�����(�ka�����3�ȷ�ʄ��w�u��	V��Q}@X:���8�x���5�Fv@\K)��=��8n���:MO�6��cS�G���e�Q*��+	��!ׯ��;k�G��ﵢ\l��������	\l�A��G֧�g70��MO�L��gw�X:�c60ah'7#X4S�����%�7�ݭԭ-�cxq��}���)��$��km�䃡�f�U��*�>�@.�6��2��0�#[/��D��P'Sp���1r{��Z���Bu
D��]Q�a��ܺ葝V���qLV�L��=�7-�4���S��l�?I���-�]��`���:y����Hر�b��dNW���$���ꂳ�v�_eW��%>��9�2˥�!���i�o����B" �l S*���\ے�5�/d�,��RYXB��#�y6nX˹n�q�4SX����-�0t����П�S�;���Cf�;Ru<n��f�D�":ş�Y��=��*^��`���}+�� ��, S��>���MA���0����V>��uH�F�@"ֈѼQE%^��e������`���N&��B`H�Y7�{j%�}b�v.G����[1�������H�4�ك {ݙ�*��1���B����7Wb��\���:}������H�f�q�_
�|hW�z��ߺ�X��ɦM���;�9��yNv:H�ҕ�ϧ�o¶p׷���273����\��"Zz>YBJc`�<J�$*�י	Tq~�8���k[eiTk�N�J����?^�q��{L����פ�*����W��┯Hy���d�D��	�'�R06|>dV/zz�����0�z��B�8�'ؖukVAU��C���&�����!s�7L��@b���#�%����
 ���G�7��!lҜe��v��cDNZf�S�9�x�C��,	�8w�����A�|	\y�fk9E;�t[�o���>� z�ȍ�Q��V*�����/օqцq�k���.����i�W4�M_I�B�,l(L<�v�x���l��	<�J	���s�46�A\�`�����#3s%G9�P����x��;�=`$��� P���?�S
U����Ad����n5,�4�7�ͤ'��ၲ��tf��G���S�!��@�8]�d��ʢ�o�.e����q�+ )	�a���{��}8�p�b�D����؀9�!����tq{	�1�y[���[���������y�l.;T!�,6l"���e��J���QF�hh�@��g픚��mFB�ը���D���vG��
ˠ�\&�L}>!G\ew�Ya��P��(/�Ux�Uw��#�0���P��p��w{���܌=���h�c�7}�Q���=,4���rj�;d��J�,~mS\ⶖ�8j�w;u�܃�Dq���7^�.+�(���ۘ��+��Y$�h��O�tOP+��Fí� �ݛې\T3����Z15�4"sǸ�����4-@�����f�х��`˿�a�7t�zg�U���a`-�|߱�'��Y	�i0QJЈ�@X!��j� �ԕSr� �.���EӕW
�,�1T��;T1�25��'��4 ��B�|��ǩ�;��6ì�%�hʡ$X�/QCNxw��n�ަe���N`���lDV�*����΁/
7�!zY#
/����?M�x�i��6aB)���ܟ�0��oO�=8xb`�Y �i,6Ե㭮Ԟ��_���B}6;I3�"��e�A�.�2�����fr݆t<��ii��{2�tp�rq��B�T��BlѨ4�J��2���ڜJ��=CP� \�0���hE���h��O�]��]J7����ua��B�B���Ky�u@�S��Lx�(����ĥ��Y|�Lݢ��H!\���E���f\�u&�@c)މۣb �EY� ��� �l��'��Kd9n^b�:�I�6^�e�Q.C3f.��ET�?P'n$���n����4v������|E�p�� �}u6 ���~����p�p�Ѧ"a��k�*���<���>�CU;�ޯ>vLM?m���VV�:U�@��e65��gpB�h�p}���R�.�����BP�����ym���nIU��!F7�����E�����&��HM�CM�F��
 H���T��HQ@u�����l9\�ȥH��̙%��f���En7���F1���'�^����=���W�]��O&0K��KoV�o�F���\1T�''W���Ü�<��R��͟�A�t�I�C�t��^�qj��������Wd�!��47�e�#1d��23ǽ���"9����o|5�%gXp��c.³�"2�X���M����	���Ծ!\n�Ͻf�O�W��������*��s'9�H?8E��k窐��t�z̓����7	�2�癯K�<�8�2#�7�����$��c��=_xJ!����d�<G:T�
|.Qٴ�T��ޢ�N<(�a-!�+?�����	T�Ĵ�����9���%`��y��P���aN՜���^l�(�u{J������U�}M�����/Б��|�ݍ�#x�r���P��#����Ω#w�ԈJ)L������Vc!�Y�����Vds�ቒ�w�1n��ݑ���%��?iK�_��\��Һ���7N���3�����+��o�Rp�
�w3���̱�~�;}���s�u��Eؽ��O(\L�@��u��x��~��%3�.
���v��-C���c���2�}��J�l=�،��n���<��!L�bj5*6K|BFv������0~�w�&�����v���e2L�u�?2
���H������ׄ�9�����x�3���&��rta�8���eCN�,�s[9��3]�P��$�&�ʇ��K)Y���UX�^��Y�X�~���Ʃ��B�+�95jQ Z3�<U��{�ؔx���k�sA���R��n#��C�\>��T�'���:B+T ��su�x�:���I����z�<FZ�`zٕ�|b�^w�&Hvu#L��B��&�$&!"b�}�/f�t�����a7{T��a��)6PR`�x)qK�^*�$��V�X��lY	���9�&�ad�/��+��Cı��{uds��zp�YGZ�S�{v^�(�-įǹ���;Iv�~Ii�T�n�@ly�Ii�}��R�X����Y�C��_p���)�C���S��gx�韾����օ7j�׹n�Z�Gt5>%��zf��^u��! c�~a`و�%���^u�����:t̮��+�uå�I;uFQ��h��&�W�^ߙ��7˖��B�C"���ojd1�m��;,Fu�CU�Mʧ}Vv�CB�M�X�YQ��P2���� _Ր�����a
+}闩�o������	�V�����MuQ¤_�zbǸ
�?S�[��:/K����V�we�/�H��KȮ̪l��m���^��N��d�Ҁ;[�UnBHe�70a��."5�2�E�0^�KMl�(�2]�Y����t#-�uV�T*��E�S�|x��n2�{��U3�X�Yc��߳�+�(�g_X��u����E\4!�`�KY��D5Zy���B5r �fqF[	��	t1����,1�jv��ZK��)�ho���@�	�Q:�z�8Y�[�}=�������/�ɕ4��0�ϲ5�XVAW��m�-^��}�]7V���Nn*���y��kj��/5�a��o��{8q�H�9j.�`y���湮�@��r�_Y}�Mux@ ��v���b1�Sn�w��`�w�V��6�8q�`W���G���"����;���[bvw�RI���9�H�c�<|�����M� �z��S�?!���1W]`~0�6�`��+��`x�F�ۧ1<�+�����%����]덶i~#ϺSӵYV ����+a�*�rȉ�P?���.��;J��QLݠ�{j�٬Oe4�n�2[~�Z� ���Q��쁎���Z+�T�	xi~~+��H�a�?��P��t
��X��X*�U���W	Nc��c=,/�`S�8J�F
�82�0d��5��I�i(��V#�J��t�9�8v�._YmP���(?
fo|��r��-�:����Yf��#�4��=T4&j�u�H/���N�X��.a(���		#���-6�w̆|F�����&$^3����7�N�2��4wd��h��*d���cf8�� M�Z���LAE�D,+�E��Y�&���~�b�_��̖���e;+������u�SԶ�2JS�We�K j@%��Ά������I�4��V�R.n�:�_��p6�QW��{j�$<�b�Ms�Ǖr|�(ᤶ.�v�F�?>��e�BF$#;�"�=FI|���J51nG"�� V@1wZ�pu���_�eZ㣅fi�� ��Vh��	���4����(�=��B��]��H����G3;�)J���$:7��I��@U�#�Q��$��cZ�#R9�OQ��c/�>q֫ѫ�D�9���J�
�����bz�@��	��vy�23�X#'8��	�8��� �+f�v�'��>��YU�K;�܈k�)l��ټ�^4�`�$+��S�`�e"Ǉ9��V��۪�r�����o3 ��n
$���|�i81�������e�[u�in�ӱI�'d��Rx*�<V�暑�rĿ�R�A�q� *ʧ5��g�(����#0paO�VJ*!<}�zǭ�����a�)�[�X���@�#�.4�v��%�M�J�Ft=kv(YE��p�B��&:�D'󳀬��RHM��K���<���5bx\�"m�E'J�l���2"���fWMۺ�i.�/���Fnկ����u�a�\q*9�ƃv��1b?m�b��'�X��E
Hsԟ飻�cւ��e�U�Wh$��Q�9�Y0�W���K|舉�,�kt%F2��v�C�%��V�_DB�l� �>� �����Ij ��i��D�%����9��*c�ü��I	mDN"����&���E�=aa�V�+�f�u�e�-�m�FM�1^�)���D����xu�0r� M���@7��	i��s�~��J���`��*��,�������E�4������V�I��r���9�W�����FX� !d2N^4�é����+7���{KH��\����R���?.y.�<�"��q={츮t���2j�r=$qھ�����,w�[�K`WM�!�5��0�#`�µ,���/Vx�&��*�|~�͎&�+Ĥ>OG�����ӺJ%F�+j�U
�"#��xn�go���������d/�>FAM�����4֑8b+ؙ�j�ub���<2�Q�dώ��g�Q���n�ڎ�ܜ��q�P�����F��E��m]��RR�%�\����5��r-��Eٴ@!{�����;B�T1A�̳<�Ŏ��W�
�����z�	M����J9ZmC�u��)�����[M����6��P}�S��I����D�,�w�n����n�5�P�piw@��/ӂR��l.��q��EZ�էK�X&L�;���*�ef��6Zg�P&cO�����@���R	Zn��6Fc\@=�e�:�pت���׺�A\�ء��gBA����is[#���	���Bo��f��G��<ǃDH �2�N�&��t�t)�3���&R��41DJ��F�W��71NF�O��p���8G�u����'���U	*�ɒxB������ѱ�o��3��t��O_'��9�U�v��|������O5��Y�_�Ԕ�+��{��8��9T��x�P���0 (b��졦߻����ot�W��؞���"	%����g���=$n0��%��T
�AG��qOfl�2\��3q��R�<��7?�N�Y��H"i��V�B��Ʉ�g�3���y��u�xD�|&����|Y��S�cK&�;���B�(�k�<M��eUf�8���\L\�A�2jd�=P��L��7�(B��:��_K�Qm\���i�a����]Er��lF�U�-'B3x�!.Bh���}lG���h�ǅ,ӞJεD!�\�#=��h7y�����f�G���d~�����-�DϽ��Ƽ����9�E�;	φR����� ���=�W䇤f7�$P��s]-q�3�@�I1C�dNKUڏ�o��X�,�o��<�p�R�#���]!��lڦ1�6�J�KFK�L�;N`]��TR0!m�(�e"0�W[��7��!�#+�@Zv�3�M`����X���	j��n��Ef�k`�~���:��a�[��(��;f7�����g�!�&@�F� ^d��ݯ�]C��X��azl��^�Z������|
K
���AX�%N���h/p�#�4���v�{��/gp��U����{W����}����6ue�zi�a!qy$����V>^C��^A��{���*�k��G� �R5F�N챬!3�DWn���<}�s0H����ᙰt���xeщ�e�P,�g�҉����F{df"
��DD/m���f`b���(�)�P\|�Gh<�hw49�Nh��7ç�9�f�{�P�b���`�Z�,�B
��&2��;{i1V�F��0,���s#�/Ɉ��� �p��Sx�7�������(�Mh���YY���Z�%GK\�6WR���3q��E�#,ʯh]��Y�B�r�Mp �+{�R��geo�pE�Fy�&����J��B4��w�G}8�O�%m�N�Ψ�����o�f-���@H����fu�n��!�5�]��1AHgV����f����v���[`q��E������<+96��x1jE��6T�o1E��<T�+2{!�Z�����r��܎�'�W�kε��7���N���!�\�eJ��vV&����P�w��d
���bfF�Bf�I��D��?�O���	  �V�=y��ؤz�+<;,�/�G�C�}�	����H���Z=9�*����o�29����9�|���.=l|\VW#A"��1��fߡ���ݪ�0��t7��D���FJ�!���G��D+�b��^��Q������}"�}X���-R��3�T�[�kZ�Z�2D�N����-���1�>�A�_����]2��ܝ���s>��>(�$���0���@咮+ ;���W�an���!{WR��D�6�9p=N�G}���i�\��V�Hi��n'��M���:,q=Ԇ�s�pɌ��f_�L��`d��7���g���T��^Y��"�	,�,�����&��z���V翔ѯG/GU�l9�c!\��8�d ���c�O�f!>���PmY�b,
�AE��k{�+v�lf��;�ՠb��;��vg��O�TP����ů43��H�#��k�N��)�(�:y~�ፇ��|�Ri�񦧴&�W��j�0�ݝt�!f�U&�c=�#�����m/��f[�^�Q��_ÖjٽۭU P~�;WJ"uҕL����eX�����N�I9s#�}ȣg9;?�Mص���&�_Xm>]PQ���Q,�6�|���e�eq��@22}�����4E��G���>ޔ���B/g��#49�/l�G$]'Ɲ~DȈ��������b�WN�!뻊A�/K��=l��}?�$tla�s����8?.32�NH�'h�uY�,G�[挘!L����I^f�g�7�v1�����������wV˩r�WH�&��H,sJ�}�-�-�8�6�ӱ��BMf�+Qy[tWrg;0=@��e�$�G�eK%�l��:�G�f�q��N���{j�J��.�0�����G���(L�f<_��$��x=�0�d�,�>a�cP�}����ا?L�8$͛A3S;�Ԭ�~�4!F?ь[�[����Q�`�H��p?ş�I�e~K�R��]B�["_�x5c U�oaq="����T�l*3O
�a�5�*�Ȫ�؇?6�=�t�! ��l�-��B�uN^	F�����r��?��U[ξ�{�3vi g�����+��e�}�ĺwO���%L0d�xwV�b�\�t�ʬh���\,a��Ќˏ40^��<���G'MS/���{�a{Vc�6]*�Zձ��XE�L���͟!�@"�H@B�zL_=�Ig4��������Ru~���R��v�?2���*��s����ʬ���]w8��#X��s�I�v	? "�����!�2y~�+k��u��� ј��S݃59���GVޜ��_�M��?�X�mbfJQ�h���f;b=�X&Ɲ5��^�#��f�8h@S�|��6I�¸s�Y�Q;��U��-︸z��ʽU�z�6��/>c�2��a	��bAŃd��	G���{��f��YM`�ߌPS�>�7��`@1U�,�z��V���������3�7W�����do�Q|���.N}Zl�疛��b��>ѥ^ƌE�0��#y8��c�1��P�r0?p�g�!���#E����}�*�/9�7�ڗ�![h`�����H�h~n�</�w�.��N:({.CS�Q��1��Y���"��G�K�je��0(�2��*�R�ؤR�/yk>4&���jv)35(u)GM�@�6���t;�#_(AhH��&:Ή��z��nIp1�J�]תJ��2�um�k��O���z�VԒС	�%Z�l�e�L�m2�8l������5��m�.��I�X�x*����i��pk��⺲��xe-�>\6�N4�_��M��0�lӜȊ�m�)�N�eF�S#K�u� g`��*���}�8ۋd�'{�3�9���U.x\�3K$|��0���}/e�T,��B����Tvx������낭���~W�\N����T".y,D(-9ʱ{��a�o]�z�.��$������r��ΗXC��hVfx0:�*����{��YRF��_�m���5A����d��ש�n_t�=[Z���3ޜNI�1i���$j�с���Uif�(����snaP�by��B��]]y����j�!~c5�@��x�q 1}t�}B��~���Y�f=+@ޘ)���đج��
��0�xZA�׽�~������vQ�ח�^�u�b���yF3/�L�	���q���e�.�}��
��������$+|�J��D�v-O��b���O�qh����,m���o]9�QL��z��*�A�n�v�e��Tу9�Jd�D�e߅�t�~�mg�����ϙ�Ϝ�d���B)8��F��7����
��K|�����5�C���\��o#�ir�4��Ǉ��F��u�8�}��;r���H���i����\��w���(�O��������0��A��t�ȱ���o���s��A,���H���
e�F��w���C��?���X���pnҷ�cz�߽�d�dQ�MKd��Ð�,*L��AZp�!�w����=\T�fk(q:CZ����l� � B�t��rOU���xwu�����,�W�19	fWyz*�i��o�6ʋV�e���O���<jdm9i��'/Rk�A�&¯����h`0����?���z�_�4 .O�M^C���ƠD��\�6څ�E�J<��|>K��8w0�����}Q��˻t�4�����'覱�h6"�&�}�)�B�V�w�3�;�n)����������I+$��������,���S�t[�2��ڐ�����>�i���x�w]q���'��2��HD��g ���&��oFA��������)��l�}�M=��N���m���-E�5�v���hi�PBd�B��A/iJ|�W����?��	B�#�5��P�1Z�c�������]��"9���Qh͆P��� �� e�sc
�I��\���.�{�0�	!Z�Qݎ��_��yמ����I�N�7'��.ږ����b�h�u^���T�{�_ΞFn�0'vB�Q� �72���e�������>
����7]��PA�)t.t��>m�QA Ou�'Q!�����<,x�H�M���7I�,F�8f
�z�1A�`��5��AѶ+/��N��~����,��������:ͩg����cI���YSަ�2>�9 ��d������Ui��?l�&�B%�)]�c��K�H�:�����u��*��L�Y�L��ܿ��f}���Ӎ"��/�^��j�#'8�l��8�޼������:�s��w9H�m��B�d��5�m�:��뭑b���'�)�҃n#rE�4
NZRU���
 %1�:	%.?䁼�x���opO���%ג2�%�<�����ԋi�z���̶;n�1a 졡]Q\s2�����mj��c�䅀rv��d����gQ8K�9�o��
�Qj�ǡ%�O�ڙ�:�t�fj����_Y���c�-��9��K5=�wk^�� �E��Z�P�i�3�w�YwN��b7u�[n���8�b^ܖ�L�/t�>v��m����V	��Y���zw��!?i��n0��ڲp��!����{s���r�ЎF2U�-��]����U5�3�Pl�ai������ݗN=2�;��C +PU��Y��ۛs�_#dU��22͝��ٍ)v�j`�4����;@�tEP�V�����ֺu!Oo0Dm
��}G >KA��1�DK�Zo^Ú 6u ��0�a~r�|o��9�3u ve�䶥a�wB����`'��6}!۱�u�6��\6����2�8�)���ǂ��-���o0�/����+�NI9 J	>Z�HT���3�{)�h���#K�����`�p���H�u����k���!,溽9
�v,�[.�S����Y>A*��!

��z$V�5P�&ie��_<o׭/d�Q	�GY�k�t7��U��nR���#����.�p�>��7���UT������ƾU��:��7t�iv��0�����mr�;�fБ��4<E;��;P�alU�>z�kC�����
l��#$��O���]���+b�C�8��;^Y����/�[W�]H:�C���T� �?<B�3���^mx����US����c����4���[=�RS��t~^@R���7݈Y0o���A�,�[zM3ǒ<_]�m�O�����"��;w�n�+�x�
O��}7�Υ`�JU��i�N�Ȥ(H��)":)�8�U*�%�����?{$U�x�tP�[��&v=��<]������GLO��Xà�G�$�=�h/��pPs`+�47�W�lD�H�"�o���X�I�VDR��"�Z;����9���y+;M��1�1ϳ�s�\�gZ�$�������������uoW�ePb��l�׈��||K����l�豈�?=�UG�渻��c�o���Zr �����ʉߜt�M �O���BP�9��M�b�\A�������&<4��G ��r.��2CT�ź��QeNn�T�a
eI�� ����Z9�p�5T�'�����r���@�7��9�?�U�	�C���������,-'
l�wɕ�It�i\�D>K��V>�I�j��S�[��;�k_i\��uE�u���UX�a$�;��%�{�EP�YHx b>stmdISjk�����L7�Ur�R9���!ON}�wc>�{��F -I1]���Ȏ2�q�!#�7��$�dG���|�?K��[W���4�~�ƽ���9�Q��ාz���lї��Y�ՠ�^���a�Ea��������3� ����cn��;P��qS�'�|�vO|8v�e�&�g
�|�U��ZڶL�8_~��_`��bNc��ن����A�\�\� �O'97+�~3�̏A%�] 3��v����z~���ܹ�;\|ĉ�����0%
�G��8��f�%�
T��wjń���I3t��k�^"����+���Ժof�и4G�M|熉Ã8��U��13P��z�зgK�� D��	HV�̋��c� ��p�+�3�>#)�[Ƀ�o�З�.g&ε�F�W�������Ae�YS�C���!����t	l4�>2�s<�������7���zg�^LC��!�q�C��j?H;א��Řx��9gR�W�K��(�@n.~�!b��ޔ$i�7=Hy`ݙkD|nKs+Qw�ϡ�/o�ښi���g�!�Fz�Gￗ
�_A��壹��`y󆽈^_mj�P�I�)쳵�%R?���>�P}ǎF�i*��R�H"��?�/��/'^��u���"I-�V#�IL]����wwA��ϐI��#��k"Er��4m�͸8��V'Yb--c{�v$٠�ȗ�����$}�ף'���%�+[�͸uo�>�Mܨа����r�T3�V)�>p��~�R�s�by�i!�O�QW[��@{�+b�j�EP���{8\O32	i��tL���
����G��TX�����Dߏ�ý�ה;�f�(�X�`�ÿG�m>^�@�t7�5�� 5������\&��##q���8̐�5���صh{B2��N&��~8idzG��J�G����]���Fg��T�?E�z���������p ?f��z2Y�v����+:�r>	(�G\$~���3�����<�s����ݑ��q3�B)���_��[1��Li��S
L��1%�и��[q�E\,T��=�W�p��M�G�:c:�'� 10���c�5!�r-��#{����5�O{�>�x��C��7�l/�$kM���͏��+m1iR�W��+��I��i$�gK��L��1J@��n`��h�#�]zHW%���k�U��8*�[vD�X��	�HQɁ�������"�Z����p�Sy������ówԽ5���ީg�,�2"[�f}�c��4M �yݟ�sV\]�X?�ґ;	�=����'�O�� ���(@�����n��XpX/��BPa�a	<�����(�LY�ꌈ�u�*�skȁ�gi��s���-�c>Ʈ*چ�V���$�%�/:B!B��
�x$�\^1p۵�ye�żI0%Ė�H2L�ߨ�lк���6�͚J�%g�l���d�O� �26���1�v�l��]�=�x!��x�m���R�N�@��xN���� ࿤C6����J��IF��&w)0�BB�ʡxӓ3l�<H ?�ͅӧ�4tFO:ܲ��y�M�S�G�ǰ$ψ�*�b�魔�|.�)�x�y���)�7=;a��q����D}J����柆Kc<G����F{Q��#��˶�D�a����tLEh4���\��%,��)D*��FK�򓼊p�:����Ăf��g#/�|IIF^�"�IX��-x����>	��\���策��J�Ep�~���A�l�E����߈3��@�>[�̾���t�g�Z�{;7C>��v??�Mt�
 ��8���ض~�ޮ������TLn�r���Q�����}~t6���H�Ե�-�d�_�4�0��;y�̊��"g		�[���'/�bE%��M��.�g]��H2tgR��Y���j�W���i��Lⱚ-��_�+K�2�X�rM^`�i��ӱ�������8b薪�Z��8z��x	�T����P'����q��?���A�.Syf�#:�ԡ~\W��c$��+�:z0�՘����[�	� #7� �ǂ^��.�ߩ)
������je�l�͈�m�����t��vԈ��~;{��ǻ:S�ؿR)�F�����^+C�2&J)/� �yڑ�O�c�
�L���Ԧ��)1��Q�	��{��h�e��[H�^�+(�#�ST��Ip(Dn��Q:�x(@g��l����)�?� �u�Ǡ$Fe��Y���uVD����pnܙ��O����!�﮻�,�J���
X�p�&��e�`��6��r�����q�q����R�nzX�/��a.ⴔr���w)w��6�8�_�?��f��m,r|�H�g���='[�(��1��ڀ�JˍvSL%.�U4kpt�v��l��;��9Zb*���:ѕ��Iw�����ҥM�188���V,�3凮;<H��`��$%�A:唸��[�կ�n:�@7���0�����,�ի�h���N],'��r�`�'�.�����h��c�]����X;E:�����K�ws����b�ulLT+�}�A��Ga3�2��׍�tz�UbK�<K��s+�s�:VY}��Y�<��˃"?,Q��Sg=٭ix۸n:`�eB��v1q!�1��������tV�g��P�ӧ}�s��QH�0�9�����|���]�����̛�hZ��>����v����5/ii��@S�ߵI�h3 8���H�+���!CT�/}�F4�Xƚg��e0[$�U��=��Y�U|
����H�㖏��K��k��De� �`ֽ{*�5G���25k1�D/�	�w\�ӳ�8ټ�K�e�b����A���e�:@�0�
�E��G2�R��<I�9�`�`��AۥX"�0Y��/"��R�4vj�B������w)�<����Q��D���m�n��"��
��llQoh���8���DJn�Cj�R`:(/�Ź�01R���A��'̖)���a�ܱ��ƛ�����&�;^���di>���:ϔ'cA�+.lZ����8EwZ���U�ݜ} ��bq.�b]�k��	gG������� �?F�
q�1wğ�J�=����i@o�n��dбJ�e���TBgw�D��֭��#�����!�|�C���x5��K<��L���-~v+�ái'�Yd�����q����m7��w2(�ɀo�֎m�ag�-uiEH�> Ĵ��'��u����Ҋ@p΁��|����������NV��H�=�;@��o����bt;��c��ZL�E��
0P� �ݱ���Eo���f`�^:6T��剈ukI�����w���q��By�y��$\��]Ξfa�ms3�~~��3���C|:�u^6 D<��5C9�-V7D�0R܄W�YZ��ӎcN�&����!4袞�	�9R��6h�(��ԯ��b,��O$e/K���+�ک�5pJ�5�g�,(7>��-�h�;��uҪv�.�?T�����O�*�R�2d?\!�m"�P4�~?칁��M�YW���˺��^�p�Z��kp�ZZj�&�R���"|��:���-t{x�+y����..�T&=� ��NQ\�	@%�"*��w���7m(��n�,`c�rr���w��=��+0����#EI��Q��|�����վ�tY0���Y��Ô��i/�e f�4��p��������SL`s�����MmmJ��6;j���>IG��B)%���$r��C�_|T]�*����],��m���ȓ��*AߏA�Գ�3w�q�7�zj��woփN�J��^~{��ϩ� �r<g��&���>E��������
���Aއ��Y0�۸>�:lP �_-$�*zH�:Yw���Go�&���/�"�W�V	�,����z��<�&<����6�Z����A��)�tx+�>qԋ���N(�5jYU����^?7V�ƹD�³�bCh�G��Ԇ���z�GF���¥�B��4Z�@��l~�A?�4Rq�8��K&0���1��:��4y�L
a{*s��jE}Yd`��^oOkY{�Kߓ����Ĉ��{�����%�>%�T�Q���g�R�E7M"}��KJAw�C�f@��ǅ#oP��}V�k��k�y&rsv��Z��DwoqO�e$�:�k���)e���gV����>M	ȠR��E�Z�G?�6F]࿑��'޺ņe�j"��h?�}:�1�I82l<�Xe@���"�ƪVDE���s�	֞p~(�@vPE�}M��|��.P���c�z �Bi��ڠi�p�+~�:V?�M���(�-!�t��!�:`��L���u|x�p���s:n=��,u������)JR��憎�q��=(�x�H3���/n0�S}w�{j,�}��-u]���T�r�t�d� �
����o���׀1��8�R�{�)�"V��@����4m���E�m�hֽ%+DՕ�v�R,�}����Z���^>�%���Ub�:>R���{����B��-�p��[%��
q,�=@�Wש�|zA����Su?�B+�pw9����<��I2��gP`"#\yQ���`��������yb�,\�&�z���J��]4���� ;�0�v&M�Ƞ��`�c��i�� N[����}D@���}^42j�*N���<���b^�E!м�&@<2�Y�l>��LY�����;d!�l	܄�n�V��)I=�q�qPKxZdZQ�uԐ!r��v�Z�DW#X'2t�ڂ��=V�^�n��A�{xo�-�e�(k�I�?>)2]�<b��|��xbV�nNέ1�o���J��H7�X�%���.�AE S���Z���Zy�t)��|�D��`��n-R%*SP-�����%�RC�(��Y@�~��tZ~����!�Q1J�z���M@��5��Q��=�����%;3�E/�`P�����K�L�Ȁ�T	,��^P#�Z��(�n拀p�bZ35v���?�y�8�[��8���]�?fF�_k.o�x<����KՆr��7���� JGco�ƛ�%z��\�C:	'I�A[�T"L�?y⟌J��
��nNT��%�4�Z��z�/��|��f -K!����������M#�*�$Co��|��M����	;�;�1e�]�aPw
؂�i������Ũ.��,�rV�D�:_Bx�l��:�����r0+�@<d�Yu G�]��$#����/MK
5X�):g�M�"h�9)7��G�rS\DM[�/���.(r�gn$l���
���_\?�O���H�� 	�`�wް۬;`���Tۏ�5*����Pc��7�����J��jol��=�9yH a��3��V6k>ƴ���DU ��ŧ�b(X��Y1P�C�߅m�)KT��b!p�QP�B��J��0z��%�iD���2MJ���o����wm��c���aO��sx�/�2���|(�2i��J��DW>Tk�;W"
yd���u-~[��?�����i:kS��,3��ʘ�%�z�u����T�k5��3�-��C K���1i�ēQ�-���ZhlN�T0 �y�����i1N-�;� �	��]dܭ�:���.��|���k��������C�}[�f�?����eb�P �����|�������8=�%�M����Z�ե��X�7�@$�N�o@�,�P�k��f��XN!8D:lH�<���H9�+���!��NH�uD�X=����:|:�0n�ݙc��GWr�DJ���bc�(x�8��E�U�N3�g��~:�@��ϵ݄�*Q'����ڗ�9C����{�����@^�H��p�@��;����s�(z�ϯ��Q��®�ƃsN��4�q�ZFm��Y0(��E{��䩓�;0mӎ�O�w��E|U���8#�ce�tm���v�`�P Q��K>�6PiKJ�/_��sּ�����
�V���]J��k�x�6;$	�0�����Pv�v���M���V��N��Q�QQ�]uV�v?S0�M�1��>�;;��"+6��� ��ŉ�xS`d�0�AFԴ>�)��nW�F�8���:8/U��۰�^��W��g�8��F��>/Rͯ����H�V;��\;�|�G�B"v�'カ���|)��w�5ü�Ӝ&O"�.]�V�"쩜�B��)���28*n���?�_����ʻ��$�Qy�w��qR즰q�0�����S��@��G������?�V뵶��:������K+�X~�
�y�KF[F��|!��'��0�P���.�k5�50I�Kv��� _��l��k�^)<Eh�4�/5LV������>����*ӰE �ɞ�B�T0#cob#���VӸ�(<7
�[�������AA.B��Kח˨[,%Ӳ�2�Ѯ��uk���1�`�c!l��0��;T6T���X!i��c�d[P!q "�=����$��‰p��/�<ߢU�]�Ԛ��S�J�W2��zm�ߑ�5���̙ǂG��5T��c�R2|�OU�}�ҚٹD����F�]mN���k��<}�b�i���ƙ��Vv�T;��4�J%�㍵�<(��*٬�tܮ��h���Ϳ�(ؐl��~�\�Xx�͛3���4����'ɟ?�� ���3�L�J"J�b�~H�
�\�0����,�z�$�b�P�]x�QRկ[�8��}��}��^ת�M���	��y��#deK�s�%GAb;����)��
(q��\w�p��v�!yl�vK��<9�R=�+��؋k4�0,Y���5�g�z�Ԏ�nG�Ў���>K����&�SQ�GP�ד��P��ȳb"����9l޷l�㘃2	BVx�Ɯ,��B�S?�-Srjfc��B$�Q~� ��J��}e��;�Mt��:Y`+(7�R ���c$%(��,�ZG���xE��1;Q)k��0wE��1����%M�Ƶ����_�p��
�0Gm��<*-���4��#��H����BĬ©�X �]$���[c�"��2}%E�|��k˘�l8�5E.'�k��oM�+)�a I�ȡ����T�
�s��:K㽇���/)�[�$�-�f���@��n��3��d@!��`���#��.�G;d�P/��B|2��&�3��h8yE/E��'�?�ӬC��Hcd:}t�����tf�0>Qu8`O ��P�/ p�'nN��:3�:3�9��v��3?��zU�x:g����a�9�C�k����g�z�*�;�=�(x��E�oQ"W�ӊ��*��v�p[�㝉÷H��aӳ��%�6)/07�6� W�����?�B��̻ ��ޔE{C;.+�	|�!��?:�KSij$�cϜI��kE��0)����nb�lS��rWt��	q`>����Dũ��eq@�J��{d�&H2c>�����E��_�){KFO��ޕ6�j�dª�9��}ևoU�\��CuOsc�D̛+ ã�iN̛>��pA�CK�'s�OAR����	,����+�jŒ?H�嫝��Qؖ.��;̻����z���	=�V���'X�����{R����{A�rAz��uU��������J/_��,�Y��a���//f��6)Ş����ë�7N:����}5z;�s��y���9��n�
��Xe��Bֈ��E�
�v�Cb�WN�ƽ�#��hU��仕�a�]�NN���U�	l�ng�ë,��S�&�'���ɮn���աd޻��RS^�|�!l�c�Q���j���b4�ԙ6
�����U��r)Z����lX
6�E�1�M��M��bF���0�?�l�����[R��S ]��׹����A6]��Op9��e@Ϭ!Y� ��T�*�@���9���r3����h�i:��he#���6�$M�k46� �ڣ���}h�c�`�R�������:ˍ,���Ч���9�[�����o�<:#�&k���{^V߫JByr4��mj}����G��:�N]�iv6�;�.L��6|2��z��c�6b��/l����޹��kj�K����R���v���ʫ��y�V�ȋ��F��i�T�ڛ~�i�7f���.�pr���S���&t{p�,����_������y\���(W�<�("�/�1H	�P�8FD������	�Ԡ�Q�O�9��d�k��]sh�4�Q�*iXlR�H{R�d�ElFD7Ȃ�1�  \h�A��X�h�*,�,��`��z}5�3���i@����yw���"sF�i,V3~PN�l�IFN�Z@A+�����C�En|����
�$]1O�55nL���� ��L����x�%��|kR-�j؏��|��$F��(p�5���f)��z�y��6��1d�z_�+BO9Dkں�6d���/��
�fK���Uw�~T�~V�S��q��m�]yBO;�I5����;*$a�����_��ɵ�jY�<3��:�YA���dVIV������{9�Wb�Y֦��XB���}�4=Gi���?������(��BW�x�g	��&DLE���@fjb����:7��;��߽����v���6
~Ro��D��5Wc���&($.<V��Ude�.�U���H��I3�Rx����w�F�
F]�R�-*��E� HCn�*G�����K�C��yߥ��G���.S�S�U��@�����S(ŠQjK�L�`H���A7���$7y)�͹y��
��y�6X�"�2	&��י��{���/T3ՄW!dp��l�a_���N����Z}J��5���{_�Q��M�"��as,���f<U�]�S��i�1��Ly+*x�ae3'/&c�r���/�d,K���������h�z��ư��ݶ�J��o��bdH2zQ��u�S��U�����$�ؑ�s�'^(u\ܱ�㕈p�F���4�SY,���K��k.ּ㭧��"\�yNaPO�Crp��+ ��:i����J�i��vr��\�9-h,�����)Y�C�G^��]����.�əJG��Z+9��C�g�1�_��&��_ᄚy�y%��lѧsSY �֡	�9r�'e�k.E�:���Q�!���+��M��:�<<�L��<*��c����_$bz�`_�LKFLo݄X�l �>��v�)�W	�3�q�V��}���p��T���Z�C�"�?��3��V�I�D�,�;F�������/M�v,����>�t���
Xhu/\G>〴m@�Z������T�[���+Uё�Ju �n(�8t_���>���VnK6Y�Us��9M��)�;�"T�� �/	�Nn<9	N��\����*�,�Q�Z��:/����X�T-�Ě爫)���0����;_��+}R���n�a�SZ��"2���0�s�QG	k*��(:��X|�Keך�[h�'5��:�;_(���K;WA�D�^��VМ�r�C[����F�|u����.Qb!�]9�/�?�~:�+���1��i;sO�B1��8��*�Ͳ�Z�j��dX���,>N��(܀�)I�v��?�t�<�8�_S@����{�]q���Xo��-)�F���6ڱ�D��W�u^�N&�[����kCk�ˣ�5�4���f�IitJt�#��8������7*�(�aj�J�G����C��Vӽ.P��[sFxZO�*t 	&�(W�����n*W{d0��G�[�-�Nֱa��TK��
]���՜`����(S�lL�'�)Ga%1�4���ߗsc��Q˥��H+2���!�Bװ���Ю����H5 /�oˁ���QOW�Й�YW� j��_��Fo[N)2M/�����H�~xh�[�}tc�t�w�t��a��M�iµ�j�_ݿ��k�͖^���?���� __/_AI��8��8C"�E���d�i� A{O���vσ~��~� ]b�Y�T�k�).�zP�<�K@>����\��X���d���A���;0�}o����M�X�̻�O1�-M-�N���t�-h��밚�}�<(I.��L9TG��R��z��3y?���=)U�������ŏ5��dNJyl�Ė�~`N0�)F��u������3%��y���ډ��;��X���a�k�g���I:�F��\g��A�,ؾx��_�t��t�tt��n�@��%�mE�����zA�	:$�֔T���z�����~k: m<�`O������ 4NA5��J�T������k�F����~�v��+̀q��/1M:x�>W��Y���p[���B��<�/�{ē*�n-0�����s$��9�2��a>+q���!����G�#�IM��!�.�J��W��+�p�H�u���I
	��)�4�W�q��1�n9�꠰�e�={,��H�-�A�*cW���~o�W�+9��qNsK�����J���1�L���>���0�bp����ڷ;C��"q��0��-1eJ�u��]���O��$dw�U��^m��_j� ������t�a��^�^ޘ�����ȩ'Y��$L!�z�����5(B4�`��m;N�»1ʜnN��*����ayf��I�B�弌�A�	�~|�(��q��{�6��T�$��]50*�|by�%m-B�~DvՑ�-��<�ob��Yl��e��Ҋ�7�%�^q�s��U%%�w$��Q7H5rxmr@z&.уy�����7���%���AB/��ڢ_%���� �c��rc!6@@]:wOcp��z=#A�=���4���5C�Y?dN���=��"jg�.�,�հ�n�g�$��Q�t�4cq<��^��N�}I��Y�r1�G�Wƶ���P1��pѽ$�x3^6�-/���L<	�=���vSN
`:�P�n.;K$	5�l8ři�ccV9��ׂ����L�����%�<��\�ߎ:�&*IhX��{������T^
���Vk��gNؙH�2;dV�J�B�s�O&��/&�J���������!䤬���F茑z���䌘)��yr`	6�]"�l7j�c�Q���U�ƼĨ���ԺR�#���	�('R�#���_!Θ�Ncc,H��m��4 �='�e������ƞ�����7�K~#j��a���^߄����Blm�;��f�v���x?�}��H�K�8�c�]�����%�v[ś'�i�f�6�����3�Tq�Eݹ[1�}���F�.�g�,Ք(d�` �J0�w����v��c���Q ^���t�)���ѩ�i�����`"
�20�*|(�V��8��U��[�Ҵ���f����$�����s��݅��1��u1�Xx�A��*�0��x�4B�V�6���T��Uo��x����>9�sUW.��e4�A�7�/Q���A[�!�׮�⪎�M����S��[s�G2w�B$�	1P���	��"��(_�V6m�f:�Y�f!���z�l���ᖞ�ez���?F����t�,�}�_���Mz���@�8P��M��6h�����N'�w�	{m�z����{۸�p�J�tB˧�q<�|�b�cr
��o�g<��:��kr8�;���(�s��Ue��S�-���h������B>��s��pKc3v$\��~��D8���Z�j��nQ�Ƅ~��]]�R������ˉ���
��[����T���.I��z9|Y���e�* ���t�O����{�s�ɷ%r�m���;��e�~SA>��*E0�������Z���u�ָ�ԹI��.���"qff�1�=�3�V���q��#��"^?#7�B){^��,,��NZ�n�g4�U=��2��l����vb"|.ъ�EE�+s�	,��Z�&��:4������8V�=>IQT���CZ�j��8`z�77��x�H9��"�f6t>f�}F�C7�OZx���V�v]l�_0�&v�	�tz��/ٴݴ���pf���'����ik� ����4F�/E�qbr�~�T!�C{E���4�Y��o���1��mKa�~�����1�d�y�(�S2�σ7�UWH�q�����p2	 6#��]z�վ�&���>�b�|���`��d�����Y��*�Q���մ��3�M�<�Xf�p��'�g���j|�;��[�ֿ����i��kN(Yʾu��e��"Ѫ2;T�F(S��> �
�(��aܧ]��-eն�%�ů���<C�G�ۢ��@HuI��t���֎Zd�	�҃E�H�-�o�{cu-X�~�Î�Zރ�UO�P��
��s���������r�}	V���L�9����Sn�rl➮��;�ė*ފ���V1�FC���>au���Q�7�W	���0mr�ü	��*_ln�s~��݋��Q���H��t<%V��垟�-q!��G�a�M�k(��Q�R�aR��P�����o$�O@�?I�)�6*=��pL�T�
�$A}3k�ѻ�K�rse�L�6y����%��[�w4�I/b�^\z�Hj�X%����@p�|L�ć�)�-�d�N\��$�2�{(Q^�G9=c ��m�EOY>[~y�i���-|�0�v�W����,����Sn@#�� �ׄ�A3�7>(&��Lq�rT��f4,����z"1.��o����-��mO#��B��D�h�>��5u��{55��5�t>�ۘ�K�����<��we���:Lנ���E�p������	����s� �;��饠��\�{�����b�o㠑l�I/	5rY�\���RY����qc	t�S���:����h�¶�t�h>���u��d�� �L��btc(feӓ���@>t��]�ӪJ+�8fш�T���7������g��e��	��������a�Y��)^��g������m�˯���b���ͳ����T�z���m�%O�HF1�E���b����r�_PϚ���4{E	�6�n/a*5]F�11y��v����ۮMp�Py�t��zO����U�^�JL�r [B��2���/�[����
 �1k1
�K��m�C_1�`V�6���!�k;[q��4��NPA�Νvhr'����"%O�� �f�B��� I?:�K�	�f0�:�ZTa�im�,l4���ˬ!Rm�a��Ͱ�KHx	�$^	����F��7`攒%N��>8�	۴X�&���o���kbNy��g�b&@�0|�ҀV�+���Bl]?�"��/gQ��� �E%�jZ�x��߅��B�F�0����P�?$�i]J�l!����id)�=2�Sᱫ�y��'��F'WقQ�_�}�8��?߶�ʙC�y�F섃'5� ���+�*���$?��b{0q3Q�S���e�c�f�"�/�j��'3�����8��%x���%sW�E�E�Ғa���b-�y6�c�PI�� <^i�+�Y{-��d��1D�4�\tD��W����ؾ�胮�0��|�-$Z�J��w��\��T�Vz�t�e6�r�va����	�y�L*�̵s4ޣ��C�c�4�O?�l),�I>�Y�X�{�L=��X͑��[��`ÿ�S$���{���A�`�������!�
>��e��	|�ZN���M����ק�S��	�ġ�;�l��fҼ�L`���x9P���s�����7+?���Jg�N�W���A�:*�Z��*��esP[E����O�S���^M��7�������ŉRO��< w������`�gF]lz>� a�66+�Yv�������U��t���[��+�6s}4n�EJ�FK��N}]6���A&��BK�B3���i�si�1MaKU��N1
2�@J�$W�UR
3�����0R�T��<N����utf�;��]�~��娆�{��ӼSV00ի�u�A�kcF��tJ1?������n|�N��s�u���!�؃Ɓ��N��j��*Li���GHҾV�{@�؞�>��I�Y���#����"��!%l%�.cqU���X���;��������p%�z�~����$ޚnYE'r�Oy���?��H]��Ქ���
�>
��f����U��<߯��M� ������@�p�l� ��!�_eT�� p�~�ǴjΕ���$5_��s�s[ ~�C�Ґ8�]����g��C#��7���\�N�c�lk�G�i�5o_��6��$l���7����i�$�K��p�ECAC��p-�pg�R��I�-��]�J+,ی:����e-2�R�Ed��|jdR2���Q��O�Գh���B��l?{C!���L��!86��"�?R�n3���պ�k���t��Jۮ����pe�|:?�?nA��[�b��3��*��_��=�a�y۴�oD���w��zǆ�-�p�	�� ު��.�%�|q���������y�e�ME�O�� ��ٛ<���z�/C<d��գ=!rb�Lc�$�m�[��F��3֧�{���q�h�1Ӡ��+-���.�PgP��O���3�+�m��Ю�U��F�=j����R&�i��&xeB�$��u^�I`"�g����{�$[>���4�2ξ-������$�	�����r�%ܶ�u�t���,o����f^4���E�f����O$pNp`a���D�������\��5��F�������+�9�N0��$��w��
a&�F��H)!\5�y[D�]#��)�6qB��i4TC~�+��1i�ĸj��kW��n�'`A���&`���U��������w���6}b�:��{sh�e-ۛ�F�VV��~ �@�wT��~7����
�
��Dbx�_�F&��g�u-�v���r<][��FTr
�jh�!*IE3V��˪��S��1�8�o����S��S�j����}��r�l��9��`bm���:=����zE'�Щ4��8<�yJf&+/�4v��H+کs�z�
�x�+�����%V�M���>�a+�]v�v��2�{���ۤ[�2�đ�5�cb������5S��m=x��s�p��-�e��ϥ�cp���Ы�9-(��8��=��S���}�{f�vS*��4��s�}�X�)/�oi��c��j�$���u�3����a)�>��D����8�bۛm3
o�㵡�)D����� $'�#,	XE$���_>4� �2~*�y�[��Prq)n�M�{Ɲ�B �bT�e���>�+N�kc_��dڕ�LS{^��GY���`�!_��M��x}*���ދ,Z�1�c���8��]��5��_�J���v��!��pȣ��Ë��^�Q��,@ �%/��o�FU)�c������vi"�<(�BĭK�uo� �r������B�A��1��X������ɞ>ҋ�E�ਮS�j(`�ȌP�(hn ��?ma1iK��$��M�nbe�����\! 
�u�1oƦvu�u�˨;�ktP҉d
	���L�Zl
|;x5�{�,uFU��PF�t�:b�K�z*Nu�t�Q�rY�D\"X���W%�xo������8_�!�Ű��O)��8!$��|3�s?a�8}I#G�.f^�F�!Yi�4򫊼gG����>]�bf�������/F��,<UxO~uWГ��b���$����,�68}�M�}@1p���e
�7%����#�]��\�����T���] ��.Op`�SA��nԮ�������o�]$��6H\b`r�cI�5�:u�����c�;��H�&n�u��[euN�jd����
,�E�PAk!���.uo���ٰU^���I��33?��)	�����Ս3�ɟ��0��<Dz6����zC��𺥽�{8&^ou?"��w�����0�ښy�8b�����	��[F�w�,�&�����sh��>�'�슑Z��0@�Ve��a h X��?��N�;\�$=O�İf��T�Ø1�_s�ٛ��y�w!��En�Hћ����2�c����CԈ燉��vO�h(����3oV{PT�2����qAl���/?9�i���3�q�tB500S���y��D!o<��C9d��7����(����F�䠺�I����xK�s޴�g�נ�U��rO~ ̰h�O6�תJn�l���}q�����)�k=�p}�o��'�(�-���H��wŁY�=z�r�p�1���EA?�n����#1�H�ݼW�-Yⷘr�x�爵�I!�A?|oS��P���,U�#-!���_Y�=��""�%3F��W�Ȧ�#I���T`i�r[����'s�~_� b2
[��d�]�B�v��GC^fUt��i�Y�k���3���O�W$����o�ސ���T��o�����\�!2��c����"�Ȃ�9z��U���w�-��x�fy{R��#W�����|����X�M\ca���n�>ߍ�~r3�f���ʘysF�wG�V>�c.��!8�.��3X΂g ��|n`Z8�j��qqy����&����������*7�!��~~�$k^��P��6SZ9�hͤ;�=�$�4B�B�.��VJ��h��7*���φ"��a��s�R��8�%�I���ď����k���)tYF�K�T Ł��E��ᵊl�G,��i�Sv�p :�-v�d�@�m�H7)�8A�[S��?�`  όH{Q����'�	�.��żS�QP��z�:��W��s4a�K^��C����ܩ7v�^�p�3��J̊�r$z�o���oK&�`9�G�ap69��r��!(�Y�����(���Ko�t�Q&0�.ܜ嶶�.T���3�#�훰�Aץ]���r1�j�&켖�� �S��Y�w��|��=h�dV~[m��ۧ�}2����hc>�~����Ȕ"��}��pS!Hю�7b?�6�/hU}9�"g���TZ���E-HI@�o�E�4�VSP�?����vf��Q�_���uhQ�-Ry��ŭs��DY��#+�J��E���f{���!8�f^*�G�u��L/*|)ӹ:))|��*@�&?hΟ]����+�S�j�s�F�g�&�FQҝ�%�Ý�����pC��D�*1��I��Nܒ�U�F9U�ߢ�� �W���:� YG6�	���#�S}g,�~NZ8@ IZB�ly9�dD�E\`7��F��Lˈ�*䵔�)� ��W�����)�t/1�>4��Py���s׸�n,�0m��蒪�Q�X�p�� ��XSE�7[)��`x���e�:���' ����q��{����ҹ��c�ޒ�y�'N�� 4�D���D�2I���!|2�䴩1­p\ZLt�l��]�t��Z:!
MS�uu�b��I?����z���Ǳ��˶��DO�KY�9��>k�`,��pV�y��W�+��@_%�XWVUqOX���Y(�~�y��Kx��-�&nB��L�A壮'��J\c!<�帿�\�}ԭi��>B� �YN�7l0���Ӱ��`�_+OY�2�N�#*f�H�#V�BK�*�4��tr�ʻʎ���3��6�^��*U�@
[5�n���N��	����s�?y2����p����Ta���"Ի���饑�����t2�����ѳ���7z���g:XR�Q��Yh��<�J�a��Fɫ�+��qǢ��;�eհU�2�wt�2�e�����ėajv������7�z3���rM
C�;t���C�X���4�Wm�G@�$���~������m[83������S��_}�A��<
��l�[����?[pV$����X*J�c�0�5i�m,������C���5i�
�=�oet��pqt�(u�ۄ��|���|�H�A������߀4�?y��z4�^���-jFd�}��<@7�;��&3�
�U��ҍ��(4���Z=�~�<C,7̹1��<����h�W��N�	[�/Z���Y�����&�7�؆�S��qI�]�}�x�q��u�(n=p}��~#믅\kuTN0���w�%۵C1r�DhOp��Mz��|0�8��j��� ���lr}�����+����V ��l��%��ܒ1L=�(��;���J�����|;��0�n^�]�:��GrQ0T��sƓm�F�x��������m��i)�a˥`��3��_��w2$���\FfH���m�¬"�;��Te�3���),#ӌ��d�gx�m�8������6�B	�{u%!���σ�D�2I�:�`%H�z�TvpE���`}�:���bR�J�{�x��V����o;���pr����Ҳ��C��8]���|�p�ݳ@ )YsW���_8����� �c�M���aGn�� 8.{ȵ}�Ӑ��m?60��g�%���#B(�kM�	�w`���+bF��+���|� �z��%���S���ͷ��{���Nlr��D���9��z�=}��Kz:�V��tA���SW����h,��ƿz}4�+�G�y<9�����3EKN�ѧv1-'ݮچ8��a}m�~�����Ɋ�7�c��t=bz��kS�T��%c�y;"�h�{0�W���e��F~[+�B}��E�|�������?��P�[��$e��8[�
u���YmZ]� z�j�F�������$Z��q L����y���'��J�,/��RU_�U�
<ȶW	G��=O-�M�$Qk'į��<PAޯ,���3G�;���]�t�'���O[�0�����m�{e�W���������+�[B�i�	H\���ҵ�
O> Y˭�M| ��>���T[sU�_8�y�_�XG���C��|v#/E/L�P6�e����M�4ݔ<�7O�|�,�cR�,�
07E����]�K��5�V���l#ݎ��p���,Vő[ ���l�:>Q���>鋕H��_��`��C�/�KN���ԋ��H��w�'��άshtۭ�� ����DH&:��e�:�j��pE�
e��Y�B������X�{I��;7J�4��DוR լ@�z��*'��
�16Sj:�#X�G������ӷ�n�"��U���&ԛ��ngj=7����2����$��β��(_�$G�0��ܟ�l-�mG�@�D[���������ƫV� � 9km?ef:�?��������L�?b�t���m����(~�|�����t�����"����Htsk�l��4��̢ ��9�e~�ڕ���I7�[��V1�6ӯR.B�Xd�ę��0+Y�!yY0�
m�+�.�Ȗ�a����dt���X����.}��&c�-;��$ҝ�s��MduDM�?O%	��H��� 9���c P�l������p~�S�"vy	���rϪG�V��>�|j$!D|5<#�'q��Р�I�X���n?����~M)�:���V�V�ه��I���C_��4@i�A�+@���0��'�w^�L�P}��@y�x�y�໭�wfoL��6�?����Il�J%�Y��]�: _c��i��]�i�!�Q��)�"0�0�����9V����́���z��X��5�I ��
 �tvc1�Φ֡���g�a��̧���2�"��
�K�[��o��/�T� Љ�g�����*�-�J$9t�R�m��&5P�R�~����B���Q�M(�>��ӑ�l�Ć~�B6F�x�(,/r(cz��cO�HK
�,��5{w����q5���ᅹ#]��}'��8}2_</��F���{��%�ƴZe��u��C7��<��\s�n.i���[��,�Vy�����,0�}�o�`�6�ԇӽ}R�h���L��n����~�T���8�۱��I�1C�H ]�@$T��5��x��!��T��~�	�R�)-�3�Ӣz�ɸ�'��A��AK5�\�x<6�AD5�e�'q����x|`I^z�}�Ϲ�1{�lU��fg4�cr?���O_Cn2���Lus�g����;���#2�_Y�=���o|��6�p���A�cn-�����J-��X+�B����B��~�8Ɛ&�5�q� #[����Ya�ѯZ�ۇ��M�%����n�b�ڄQ^���KU�[/(#�	��Ad�!(�~��/a�1��0��Ei����s�
N�]����4wӬ��h7�y�BXo���?N�-�J��<+Iڥ��ŵ,���ʘ�� ��$����P��O�.W�CK�i�B�X�$F<[�M+5.0�H,}�}yj[9������|z�vЊy����r~�&\�Z���~`(^��6kce+_��-j%ء�]���$�b�U�j��v�x�p�7m7 �BA���2���tG���1ꅺ��kD�Թě��z}OM:+=B=#�Ф��	�,��o��@E��wr���gPPG�F��;�X���]6PӲi��_Q� /�!��(��?+O�8$�[Q���p�6�� �(+T|_&�
������Z4�� ��h��:���Q�����������T�yĨ��U�`Ys�D����3���#��"���,H�C���q�*
	Rp<�C��E���� �V�g�pT�b���Q�o6�!X����o#�j�k���(��l�`~|���!��&)}��ۚ��Z�(׌w��|3���D�v��f�� ��TJ&X�)ɘ��ؑ�?[��$(iM��)�Kv�M�5D4Լ��x}P#x�b��M#��dY�1�|P�t�\����%���'/3n9�������b��Bz֧�iEaT�=w����Y�BS�E���O�1��}�@)٭1WαXEH}����ٸ�d(�Fn~�`�.��t;�)���.u�Cl�)�YK� �f�_�<����]�Ӹ�nu�6��<�h���������ٯ.�o���]'�g�1�NJ��8'���''���Ɍp�W$�d�C����x���!}%KX�R@R��W���c�Z��D� �X�u }T�`8O��S�M�٨�w�m�k�=�� ����o�9jѼr�I٭��&c�˪�b�X�^6k�-��A�}y�c=�wn#��E�q�k��u6�I�Ӛ�6Q�ucm��}F��� ��������<��<)�vY�`i�pᮛ�g�d�4�������1ȣ�^+��sXI8+�z�1���)�~���g����8e��f���s]v4�	>�Y6*��c���MpXKo��+y��=���_����p�c�ʾ�SA��D�����en@��G�V%/K
re�!�Mh�^�6 ,�Č+`F�w�N�i
�G�1֙�$��Zu�@!nI�M�'���Aɴ~�^��}!�Vq�3�c_��wE
���D��o����I��:6�zo�`�%QMmf����S��z��g~@���Ng�{��PZ7սûݝD�|W�q��� I�0�;YJ�ƑگT��s<��UI��]��SC�lp����*���W>��ߒ�
R�9b�ݟs��\-���!�-4�K"�)�`@R��	^����#�\��&E+w�y�s��b��77�;���,>����N)�Ird�`n5��%��=���x����[��c�<�Ӗ�ގS��
�pR��#�;�T����ƞK0���Zs�ӟ1>u��Y��gM�(�8�P+������X��!R(6xA�g	
��4�ؑ�W�ڻ��S-[\H�r<HRS�un�N�?�g�)8��h�W��T7�
��_��@S�#'�U��p��.�
ט�����h�ǹ�D����Ϊ\�O~�"9��&~��
c�Ė�q��8Y��f��.3�1&��s���Vp���.�Vb��~��E�Ɩ��fd����N��K���,-i�������q4�;2����:��6nF%Ϡ6s�
L`��1��٢*�ZK��z����8��+�
jE�OG������4c�V�;&�Ȫ �{&WR��VA�oـ�^��-�[�"�Qz��4Y��a	�d�n�A��иa�SnL�S�����R����e��
��W�E��re^��ß_��ː�4��Gck�as�`� ���C� ���+u9��)Wf�l��� zq���j��qΒ��)(��5t	`�H0�N�|�f1m���fǱ�Q�@�0�6�W.
K$#��18&�l+�%�L_�s��~$`����w�I&�c�e�7�g��$g�X��E'� �zU�����d��sRW�*��`�C�ơx�u�%�k9T�N�QB3��.G6�� l{E�Tu�Q��n��Lo���ǶօYԆ�fu7	��*i�K�
w؁�-;����r�v>C�����CH���,�~�ۧ'֎W�q��0�w9x!�n��X���ѯr�Xd\D��8$h������H�1�gѥ�5ע��2m�e�CF\���P��E�'�*X�l�S���j�S��Ʃ�H��KoaN`p���]ۻ�܀F�9��{�E�7
j�(h��J�b�"v�B(��d�b�m.���c�R��F��.뗺��WTY��@�4����e9
��ϻ�F2�u#��J��_�ӝe���<w^�)���s� ��uB�����]�<t�K��*X�q"ŉlj���,�3��j�����>�)�<���5
Ҩ>	*ߩ�ޑ%�d�iWo�_:36��#����Z��xuɆ�G��^(�V?���z!Pj)Q�p�ZD��[�g)r1���l���+'�g����6�`�oW�V��G&��q�ڊA�n�"�O������t����\��B3�V�N��ޫ8h�R������ע�ɦ�M�������.���������\�Փ�C|�T���������|�6����86�1H�I	:tgDI�#��$��b�f����)�_��P�<�o�����9���]��R:�x���U�oV�]EΚ�%1�&�F8������<�R�xa����b�����%�Xx1���x�-wa|�f�-�I�h�<@o��Qg����;/)����HA�%Zk��V�Rը������
� ��s�@��7�MM��a8����Q����Ȣ
e_�|8!8��p�J�Dr��\���s0G_���D�!�n����1VRؐ������� �`b�,(Q�gtǼ]�t~}J6Bȯ�o�Y��V�9�j'XO�S��A���9�(Ye�zc�h�ה @�sv�PG*Y�x�Ɠ,���x���%f|4�qL���ϕ����:)�AJ&'�`%zbiť�q�	�_�+<M��ދ�f���H���=k��o�����D�f��L��-�V,�Q��uϿ>�d!�l�TTRînR�b���c������s��
���A0v��A|��M������A`���Y�̈����"}2��w��=��X�y+���T�g�R� ��V	�X�ʘ	&���%P
'+B��rx�rQ�®� ��v���D7gq�E�B�W�*�&����ӳ�fAK+&�B�8)w��R��$�i��a3Z�s�m�Դ����z�1���r�[x;z���87d�]��"����F��Wp+ŗ`J����u���BqOȟ��:�ZLiT��^*�&�@��wL�"%��dX����5�i�G= �1�ųݰn������7�k,zroi�2�}>G�^��lG%s��&���y)d�ހa�o�neo��rrԭ̑�vT�h�xA�ݩ�*n����!ęL@����rAl]���sU�mA�KP$��a�h��o���H|G`���}������`��Z����'Ձ�����i��umBA~յ��`6�NA�FG���Bx�8�(N[��"7CBXL����<������,`�%|�{��M�y©ӥl��h�
A��S�z�8Kb3;I��0=��HR�%3��z4ֈd�fRn��`B�n3���|�nk��x���]�Jp*6+Hu�cZ.E����Qٗj#���S=�4��'�Mp�	��d={�ŷ�R.��X������8�ޒYm�T�Ҳ"7�A.�%�GϜ�3 �8SWDX轱���)o��P��'��ʏ��I�AYb�n�#p8����ƚU�j��҃�dH+��z��*E��.}Щ~N��t@��*i�(C��ZS� Q�<��o4�C+��u��e�1��CC#���`���.��3���B����d��Z᧮F�v@o7�;�F��g�Sj���ҩ�Q��ƴ&��w[N~(�K{�N*�}�X�	qF�嚒#�L"L�yn(��K�-��u�ӧ*���[%}t��t��g�$6,�f���0�{D�G���vo�씣�~!��N�"��5y�P�b���B-`e�m��K�����oJ�"�I얳��S�^�f��Wܟ�!���Cqe�.I;5A������&�D����;�Mݚ"H:�U+?����VП���԰Enwtkan��E�����凁�k+߸ ���r
��k�	��y��?鷪�������"���x_�sY��r��4�p��kO�F��X{?�Mc�O�3hK��`����0?sdN���ەS�;?t9�����!��ĝ�k�e>y{��\bF�����;��vI���]��p!��6�示\�U��)/��K�_�k{1����J����v:��~���
��oC#^�X�9ED`��XDxs��R*�iٰ!��j?4�LQ����E���š ��|�D�c��)KY릒�IA�;��e2�^���d�Ε��A2���$K��u������r�뵰�&�K��I�s�����ӄ�4�1x���S�}Fl�Մ
����LGF/AŃN9�¸� ����Zq""���O�_����5��"T�\��_��Q�7�'�Rb����pn};n�Kyw��-�[-�c�y�@��3��)S��k�ޮFU�M>�AA,��",��z�3�5���LH�5�n��U���z�]΢$-���������6B���Y_JgFFs��n\�	ϡl%��D2�%�F�;�ʦ����""��eYt�)�y�^�oM�f�Q^$*�Dp���>4��u�Vс���)0�G�����L�����M���1[�D�a��9R����L+��3�'��o�:����(G�[�s���ѫ���Z�	�#=���}�!8����߰���%��>��D�f"�vqd\>/���Ȉ� ��*��6Z��!��C�J]\!�p1CMn$`ŭb��|qLo�6�&��CM\���{4����],Yb,���)1�c�mC��s�K'G� �~y)����ߑOL�H���S�����BBj��a&%��`s6�L�@x�z���-��HNN�ɻ�O�z�lUP�uT�v;6�c���!��7p$�g�TIq�\(~m���e�Ĭ�*0uv��M5@5 5&�����{���-�[\�I��kzv+p�U�C�u�= ].�$սbD=KRu�,F>&$JP\�.��
�: >�$���cu��n�������CU����u�'�tY��LL�""n$�鳫=OG$��Z���z�h����6�g��}��?��@e>53���ޱ�N�KT�1�ў�Y;��C�o}�H�0M�L�w��h���sj�����BqҊ��k�)��z(#��\��ODZ�a�e�1Z���IƟ
�o�hH���i�����	$�����*�P�Z��֗[NqP=�ӔO�<��B3+��3	����U6O�Ej��+�F0q�L[֒�j��W$�K��$����E�(OM�F�-�)?�qǹތ���_|扐1r�q2����r-RY.���^:�\���ۀCG���K���{�tRn6�)�B���;.� �a����cT��bS���m�3Dǟj�²YC>|⸋Qz0��m���u�4p�p���ڭ]���.$�`���Ȱ0����n�[��@Y�
�ov��<R넑M�~2�Yu��N��e|�«-0��A�j� �$�Ty�E�fkS9�pӧ+��V���q���?Cg��E���_��N�����UW��ĹO�Mѡ�x�1T�������|E�y"�#'��2*��d�kg��!8����)���M_#B��1���ή��!z�赑e�F����E�V���[#�L�8�����.E�H�������d��Ս�^-�j:�,��<� N��)�/�o|e�����T쓼��jKRD�W�i�)���E�ˣ����W�nJ.�n���q��wn�Z��h�p����]���0����<}���`V�>�3ޡԱ���T��7=  ���n���%`1O�H����Q��BW5�`�9���&��̸hK��WJ|��ǖϺMw�6G�� �&�pL���̚�k�S���_�����5�BSج��0� .r�X��֣������-� �p�u������a�<�#*A����y�����Wι\�Vbk�V�!��r��_k�ȿҪ�]�ڕ���ȡ��x�i�r�Y[GA�Vf��l��,�A(Ƅ��I����^�����YC�aVRm��}W�;������E_�p�O��oYS������ҼlӦ�EYJIO�3�N�x�"b�����	��=~d�1[��]��nG�3��9Ct�㐝C`�����jj\�3A����g��^��
ДG��&W��{�f��]�^'��d����Έ��߰`�ֆ0uc<�&yeLHg��Q���F���3N���l&�aS�N�m�����N���j͓��i��C�>k=x �2����*kt
�L�5�zY���Ҭ�t�؃�J���y%Fd���]A�}�A�ѳ��,�j�0-t��{�\���./��ʰ��89>���7o�4�1��#]|�՚��-)J���eH�c��O����х���Y��@���Tl���+j;?G^��!�9yB�w�L-�S����=����vV��L�Q��ۗs�����,
��&�i�k�J���y��~��ODK`J�[���#ʭ�w��"j��m�p7h��҇*!���{S �ypsy��Gmn'�� ��LYڿyf7.@��F�rSo�S:#�=~8\֠���h�U�[hn;�`��6�����2]3�ЪJ���R])��V9N����w�D�j�  �MS�f9���Y��F#`� ,^;]G�9�G0�Ѐa!����e�&��%]�������	G����ȍ4�0?�} ,9oT(�K-�b�#�{�[��+{6���"ԧ�v�����+�T���R ǉ���/ ;_��n�`!�}j�%w�lP�8��L���Q�؄o$��(��+d�η|J\M����� ��G�g�@���e�)��F4*أ�����A����"��y���xb��^���]���<�\N[|��j�!i&HZ��-%����j�Z�����)k`������`N|��{�m�{`u����J����R��O>;e���i�T�@&R=�h�-4�0�pH����g�f��
C,i��q��KY¢⫥Bxt�j��L����l'V�?_��,X|o8rn�4Bݶ�'9��7П�A�ڄ8���P/3��@�i�<Zy�˗�8�e� �]3QeW�i�
�Bz��Ǻ����T��y�j��n��ϕ��K$�8y��+ͪ"�rB́r���>�̷w�-دm{�F�s#�%��C����1��, �[��!T*��D���j���v1]"���ӄ����\�
����K���\�S����%2�RV�m��U�{�Y�X��¿p��kƜ��=��=UB5r.���B�L��s��f
�i�Jǐ���a��*���?u.	֭��|�h;'`rG��0�3e �c_l��ax�n
w�.�_����/�FW�%�o�u�мT�ל7������:���`�k�7��Z���V0{{Zs������2lP���H�yoz3�w��������"�a�`_8N��lb_v~F�r͜��N"�_�`��CJ����u~�Z;/����%X%I�r�}1��/���� �Ϯ��*�{���uGk*�)4���}���[N)�ɵ�E]�򄰾R��O��F�~dR �/u���qC�Y���/��"$
����ޝy��k<��^����ndB�:3s��u�&�[N�¹ �f�J�Q
]F�� �u�[��&���E�`b�����<���2�c���/n����^ޝ��Z�c���&���C�_ �b%B���L	�i�SZ�hH,L��Ǡ澩	>��U�XA"CVDNf9����[$z�qO��cu@@��[z*$*��<�$V��_��I�ydH��D/�L?�H�Eԩ\�W���cl�c�QL'L3�/ɮ��8n�|b�v�p-��=�AQ�I*�x����-(�W��;�ޣ��l�
QY�{	�{���\�lIh����7R	D�K�l��o�נm�W�!*�����S�gq�5պ��m-�R�K>՝A�#a&�%�W*�h#��未o�0�Ϻ$�`�(j���V�<����iF��Jӳ��F#��sQ4fӄ�i�,1���.� t��b};aޱe�i�Ic�Z��;��%N�. a-f��`�p)�&�[]&n�������Pٙ�g�Pg��˷Y+k��S�j+�
uCI�.�O&�%�0W$�8��=i�D��a!��f~���e
B�?m�y�(v�{��R�Z8a��������)��6�Xl�tE&?'�r7���;�&hMF)Ԯ܄�Hp�η�|Pͪ��Eط|Yab
���N��xz���7fw?���msOR�~
:�SК?���s��`��O���Q���Y����8�y��ӕv��%�}P������p��-���O8���SS3	W\�i=;~t%�>�$0�¤��DCQSn "l���>����j�t+���a�F��ጽ%�f���|�oz��RIe\S��1U�����<j$���@�x�*8��������|J�\ =zV��A��(�^J*ka��fZh��x�9_"���<N���Y�%�@FB!0�5��:�Bk"(��A��%^��1[��: �NBu�BU*������D� �K��E�ޮ:����Z�0�vF �Ʀ��hk|���v#߷��%���(C�LA^\`'���e��SEr���^�*�w'��0ڡ�d�?��|	wɗ������ܿ�7l�8�+A�`�m+o�z͈QX��Wy�f��%����Z_���3
�Ô����~�tq��E�ޓ>5��]xU��2�0���>}�Ȱ�xr).��h�(�@)�٥�h�� UEd	2/Mx�0����`�[{��������g7�i@�����te�M�7��tX_��X��Y��������+�>k{ѽ��LA%����R�wְ}�_��	�o��۶�ޝV��_/���)���9FR`#���q�`��HL��6)#��O�	�i�y����x����4�'[�����PaiѮ�I��9�Yd`���ͭ�H5���~<�e�h� ���Ã�*n��}0�t��
�,��}�R�!���/rxf�d�㵩�]!�l����ZgŰ���3�jͥ�$Q���Dph��.��U������@���ƌ��OO�9��#�F���H����?��=²�.��e��*��vʉ-9�"�Z�!����-jb���ޔ���Sp`��ݍ���AD��d����4�ƽ�q��+����@U<+Li�����3E_�[��u�c����"�/ߙ԰���l.�)��	c�.!�Y2��o��|Ù|y�x;\娡���-���vA��כ�%��aD!z�<wiw+#	�̓�hT��Fsf���L��ӳ+�7=�%���{�)\��>=�춛H&(;�	Î�O@����-�KN)I&#u5���*i7��ݫh !��t��+�`�Z��C�cO�ú?i7�m����Ģ9������^=O6�Z��h�lJ	vN�C��N�Xm��o?�3��!9D�b�_�������GK�|�վ"�[l0�={�"�X3i"��
u����8U���r��X�N���ޓ���3�|���T�\�i���A.p����<�Y���Ѝh�g8��J'���P�eK�Xw׍��[�h���ђι�b�	�)�9]#���X$��=�Wc���q���F	@��f���|�� ��>�Sw���Z+I,�n���>�	|��d�F�IFٙ7F�3���ZQ	���X�[��/*���2�#��sSQ�|�OY`�v�~��[� �/��r!&�\FW.��E��?�Dh���e��`A��E�H���81�>8��K9z1�$�Oߺ������q�?�������������"�a�z���N��O�N��&1.I��q�_5(bf{��Cׁ�W�S%�Kۈ��Q��J����+ω�>�6=���N��j|�X�-������I0T�
����mZ"/<���"K��C��ePC��
�]�O��9�RO���¡�-�3�1����H��1o���D��e��ҡ�ڍ� ��>n��`��0L�;<�c�Ɨ�<0��j���X�%�n�Lt��Yo=w��k�3駅]�")�	*��t3r���ǜW�Ϧ�~V�TW���[�����(%�b�I�A_��k�gw��xZ��El�Y'�@�!�T�$d�'�Z����|۰��Sm�L��^�ũH150胿ح�Y����`΃�!�E�2t:�|��σ�ӕ���Ȱ��)},�`��Qr��>䜗�A�8����d7��P �[(�O=~�n]���.޾�<��?k���:)�B����@��Qéa����r~��6���W���hWC�F�96�Y�"��E<����*��`l�P6`
5�9u*���e�	
��ԗ���N�d)LcO��a/����%�4��2�{��&�)[q/����ɏ�daR6iU�p�́�z;�o�QyC'����X��S_�D0}�f!g	�m0dwz�џ��В��MF��/,呠D&2������ɦ���g�k�(��[��B�c]U�'X�0��uz��'��� �k g�#D�7�����*�~�@�Sͥ9�>��]h�@@r����>�O~Z��Bb���a9���:,DD:{��ml�&~!:�$�PiysㅮR(=��j3 � x[N9�ܲ/��G�������[iM�����s�Ǥ;�B���.<7����M0�e��f���kߺ`G�s�?�q��;G�"�Y�U�q �"ic�[������0��0�(�i%��9%�����<����%zO_V�,�'�ȁ���F+�m�'V�f�nA�E��T<Hjvg�������#��!�-�7%}��L'i
��H�S��4"��7.�CA}�v���ˢs����ߣmX(�@\+��t~ho�n|#|���cb�q Ø&Y6�I$�����t���B���ʰ7�%H3X�7��!��)D��8K��~?G<t�-�`PvFl�d�,�E�&�n��.����}�zF���=W5Y\~�'V7��XΧ��L�������%�}����E�W�i��QV[���G���f��ڨ-���_/j����t^��E��j���$A83���Ay�M�gIlb�_&I��Q"?ش���g�7Ij7!h�9,�6M��e?��"�O�cX��7FH���������\���̞YѶ�%i��k竉&�U 䉌���pe��ʠ�ډ����G�p�T�٬pIG��5]��z��O�V���1�Hk7f���y��,�X��܉Tv]�)�l,{jm�(�%��f��F�2�=7~�qӼ��3�@����_�[B��W/����x��V�Զ�{��, ǂ�� ኁ��PvE���pY�h��h�=�AA[�Q8�A�Od�'�UNZ`Hk%s�L|x#���*�-B��J�1n'�+C��7i��с���X�Oհ=1#s,��c+/��%1�/�<�&��"���� j^S�&8�p�j1�z��������|zE��G�rYH<�xD�]*�SSs�g�>P�[B�	��I�)����(�<���GۊV����IV��9� ����*Xg�q�b��O�`n.�C@�W�s��x�\��T�l�˳O�3�=����կ���Z*U�)�Ԇ]�Vs��T��?�أ�x86x�IzOS�k���j�c)�?������e��T#K��6�#�ۚT��d�c}�F���e��%���� �q��c(�_4؉�Z�V����ǣ��Х���Eؾ ����Ԣ{��p��x���|���̚�4�fw�� �J
I��6j�?��,2{��3ۤ�M}*$��xG��yߟSy�"��U���F���l��uaT���@r�[֬W��W���$�E������=h�\��ˋ��F�<3SPo �	 K�8��� �F�eu`�eC0�����W��{��r�C�� ]�{�ҷ��'t�WIZQ���fNvZz�B8�z���v�\?�pX�#�$��ƶN�+X<��J��]�r�ܯ �Dd*���4���d�����z��C�F�o��Wg>�Rh���G6S8���z&�CJԤ�v�7LpA�]8��J8�iy�g" NJ���tR��T��~�>�Fi&�;�W��BJՀ�vI���Ń�a L��ɠÙ	��0k�"�f��Id��ע�n2��, D[هE�z����٨��������PDI��mY�é�ّ2/X����#b��ثɺ��t>�f�h�d�6�=��2t�4U���pR-�ذ��\�����|PN���k7�E�$ܤ�an����*Vu��us�:'��|����}�l�
��\�Z�o�7{Qb�ɿ�@��91��Y=����ZI�̰f�\���֔�&Hqf���	j�*<�J�ˬ#���0I'��1�3�*�+%�FYT����ۿ"_��J���Y �,�h�0���1o�aߤS�qש=�2˟}*��yfG�)���i���G�" ���~rR���J�c��0�3Y'��e�/�yk�x�> �:���mM�{�����}q��#&���V�<+,�t���3
�w�ۇ:*�}"h����@��"�",���'�:^�����O�B�y�r�a~G� ~]�*%�U�ֆ4J���0�����D�����w����"D����Z�����RӳS��D���z�� ��ջO3l��ӑL��yD���)#�����!ߦؐ�&_K��gR暺�$���&�!���ॖ
R�L��<4Ѵ��������~`���������cߠ��?��ܠ�\���
,�Q���M]$Y�Ja�ek��,��K�g���1$�K_Y|��.�&I`�I;�^P]��(�p�c\͔��fK6BpW$�X�u�D�
�GiY]3�[�rņɶ|��R��fR{[�.U^4lO�m�9f�"���{�����u%H٦����"34�gWgȪ��z!U��aƟ�L�ݨLƣ%6�\B�����U8F�����F�M��9S��`��J�P�j
��#6-����������E�ކ�f��~���ج���$�f$xy?P��w�Be]&�E%��;�f��)���K�̮
l��5XVH+��f������}�o-֞H��()���.�XiF�FĦ�y�AVSv����Q��_��ڋ�5�;tⲔ7J`TjOnL���z�k�$P"��w��CE�d�R�U vl�l�m��ՀW�Z15Qg(/��3�4?�\�l^
���T���%��G�-zj�*w�¨�Y�1L��+�o ����֭DWa+��˾+v��&�H[].(hώ��i����H�i�MR?օ����>2�dNoC�󹽣?O��1gE�j��� ���4����wPp�f��=Yfi�.�Ui��j����J�4����%�)�������te���y�7�b�cҖSwε�dI�����[_���59CW� ^勳���� ��V��jK�������OM���[W�ޱzu�H/C�l�0�2���E��fXS�i[	��2��I&���?�vdѓ�דi6� �7�Y�7�����U@�Z-�v�1��W:���II�>D�MfW O-A-hQs�@u4$���{7�S�����J#�K]5b���4tK�G�����!�KB!5�x%��R;u��2��&8O��X?�j�u�	������S"-�@�G�NM>�� ��6%V�-E��`$�_���rS]f�x�A��-�x�N� bo��g]8zfL�Jw�����Ɋ*�"�@�]T?u6si}u=]7|��}�?*���)t��}���P�e֡w�G&�PB��X���^~�`���j�p?�S[�)˒�0ɆO�̊cf|��S�f���@킵ͭ� Ybw�u�P���Q'�]���3ab�y�<��ZT�n�:g3R��?����{&��\b*/1V��wK ��GY'7;H�)�q�.Z�Z���c ��MUhz�ܦm�
!(aY�����S�(C���iY_�e�����#g�g�.'Š��3Z����&O�P쾧0�F�9��C^u}H��5�ۨ6�kw���}v��t��eR�c�6�y@�Z�����.��l�]���s�O���aR�MS����3i�Awqrj8��`�Efwst�ԓN�k�L�Ľdd��?w�%tZ
b��(��q"��>qs�ij�<�y��<�O���p�<D~?M���.b����������B5A�l/�x�dX��%K`�}�dA����RmJ%b2�X������-d>`.2P�dv��ʋp�t�y���VNl�������{k���H�(i��rQ_�:�z��M�r�7ُ7�H���c� o����xf���}�q04� :�隕P���`�);�,�^^5O�C���a����2֘�@�� �-]�<
G�b|:V�w�`�'&��������Wl���E��g�r�f��aP�7^UD���#�*��ğܞ�)fI��<ƾA�<�gQ�P���k]w=��+l(�Q��8Y�Y��Q�M.��,���Ւh����vOJ��CT#�m�=̈́U*N��A{9�B�,�\����N���(d���
ܝ�������*�[���ş�`��v����h��qq4B:�Uq�������VD�����z�]q�铏��2Ü����sa��.�H��{�3���x��c�����qY3��N�J��绪���f<��m�L�;;�W�����n'��j�GR�F�6S�"ش�5�'5���	mÙS�z�=���k,{�yu{r�#�;/;�{:JP@Bu�5�iKip���������A��9�~��g�8+�$w�{î�Q�'�����ޞ���Ƹ��|2T��G����H��@6>-�;��&h�!g�'��8��&E����t���D�-Ȳ��nAgn�J`�ӽY�Ż�ڗ׵�|'����M涔��E��6��
�Y��9�@�u^'�S���l��<iJ����Z�8ް��S���4N�퟽�$�8uf�
��M�p��]��imi���H,!3���<m���$����d�o7N7�g�j�?��>���ۊWy��?1訸��8���8��
��d���/��`%�a�ۭ\�u��W1�l����O�����&l|�5�E��¹�՝���Ky�����~d޵��~s�f��l5�-��x�b%�.�D�zlƩ;���:6�I�+q��F�uD������,��G���\�BGU�"HP��J�0�*�oG�M#���"ߔ�X��j�U���`]O��{�=Y���
�9Y��kauE?=������N&���u�����xRAb�Dp� ۥG �L~�^����F�-�4
�B�{�BDم�!�\���͈�s��5"Ȟ��ȝ��>D�����w��.����G���d6��gQ�m�S7A�r�|����!w�rDv��B�����<�abby"��D�t��_�H9�^B_�b�\x�@
e$��Fj?B¨t��o/g��h���?=���d=ƶ���c�'��@*>	��R/������<���)H�0Ŷڙ�.Kg؎�?Jv�w�'m�==�v��3�Ҝ��

����4aa�� ����'Mb�;0��f��,��6����};��?�0�s��,�]G/�>��%l�-=�S����0��;n2���c�:05�I�X%�����j��z��1�ʚ���0j��U�A���v�6��^�͸Λ�����O4-ؠt9�S)���(��q'ꭡd|v/ ������]�ֹ	�(#�Ϩ�w��^0<V	�x���~�(�"���i�k�ז�h��⵽p�� B�)v!��U93�ُ���f�.+�>Q�[D]��8����ar������D�O�)b�����{׷���N���U�9r��"���n�М�[򘢲������qћ�,yT�{^<�O���R�r�Q�m������-c�7�v�.]@�7���f�R�rB�k3,"cp`��:��\ݗ��K�JD��oц\q���SK�X�T�!Aᖉ]��|�.?bq��(��g���&�Я;l ֩�˟�p71�e���s���ۧ�)���|j�ZF��Y�`� �\}"������W�Q�YJ\��Π��h|�Ev��1F��xs[���'3V�F�_�۾|�\�q]��!L�b�Wx,DG���я�R�+����5� Tq�L!�/@A�u���-�������~�(o�"���K��<��X���A�|=�_�C+�ْ?��"����I�"B(R���Qϓ1�NEN
w(춤R��z�4k �#5YߪB��Z��������L�v��!�O�TP ��5-S��d��?6+p�簷���2��j
kߤNm���'�Le��)��Xn+���w=�j��i�w̐i6��L:��@�K�Y,x���3�]���t��i�K��*��χ@&4'�j���|wk5Ry)x��* �_�8��Q���B�w��ږ˿lblw�I�֌�x�aK��<����	�aqFN��#��nV�Zۈ���g�#0���W��W����.s6�;$r�d��|�Md�����F�.��y��T��<Њ�L�����(��
����/��=�
���I��j�F(�_�q1��vú��z?N� $	�u���xqh��E��%ځ���[+���d���z�T5���E�q�G��)���a�I��8���Fo�,�z��'n�P:ҵ�R��,d���H��e��ة����ݝV]�.�n��Ũ��Xtv��i�vD�����v�v8�1+3��l}<K��,y�!� ��Ɛ������]v�vGm1�z&}�NU�Z��m���c���7UM�oY[�ŀ�ʷ����n�`��?�!��ʐ��r��dI-1B����^?�I���D1t@���	f�"g�
�o�=��Tek�5u�Rx�L�?��j�E5n�W@%�j�/�˸?J㓗�2Ub���U�>Qo���i��*G�uշ�c��t�'���5�s�X�f�\��~:Cr�\,�ʦ�v&uu���[�0l_"]y"4;V�Y�a�髼��t[���:�H 62��u)��#��3��8��_Q8�
��N���,@[���� =6r�uos�	[�\Ai��ˁ�q��v��~̻a�YN���'���vE*qঈ�/_$�O�[b���-&X���W��S�|Hɜ��u����g�q�a�|��+����n_���؝��Ƈ�:��j0����PSjQ�`�����!;�e&uŢ�y*8t��֬<z��e��ҽ3{;�j#�3�oGY�����8�$�gѤ8!�
�E���WEI7~#�a��cHʟ~��|W A����W��Bky�Z��)�5�{w|׾����|�Ө���F<�Q=��3ɒ v���R�W���	��0~�F��[�&=�4�$�}�\����;� � �	�?� ���{����9�R�n��H���š6�iZk���*�3�M��΢MyEIa�14�`gR����NlE�I�(r�tu5OϵN@��.�9u����QѬΈ�6������+E�E�Za<�V}����uI��r�sQ)���q�;_��<64��5���6"?��p��i-��Û��e�Ϛ��TL�ˈ<�3��G˷r�v]}w�Tn��c�,b�_
S`��3���ߴ`�_P�8:�P��	����y[;�Q5]�y���ꇠZq5�
8$�P��a��.���B�d�y|�E�5����mׇ��@�'�hf�ˎ�[k@y7~@����59�!bʙ ���������׸��`�lǕ�-	�ݒ_��)3�Ps�B�h�63KT���&�)dhO�*6��b�vU�-;\�؀��D2�����;�x��f���&��UX�)U������#�����ۭ?�ٿ����Uܦ6Y�oh̓���3z)%ה6��D�(�D�fb�%�-C�XҶ���(kۉ�R���=��g'j��^l�:�'���J�>>� �/Y�$�K��]HU��+��3�I�^�+f����3�u-J[��:=�m��3t'��--��h�H`�b0Ls0�[~Yƫ��f?s+;��K�s`���Q��Vp����|�(�nq:P�9~{��5Ǫ�՞@=d�IǘB�z��Y��lU�\�Z746����s������c�rO�(:L ���i*�VZ��I�;�)C��ÿJ�
��z����l�>$�zt�Djw��8fd�}�:�6���� x.���P	 b�|�jD��EТ��P�/�Ҝ6���vu��,^A�PR�����\�3c����|��y{rO3귃1�#��ۑ�	����'
�@~_��H�i�GkJZAXG�M���x���\�"< �m���d��**::�%�B��s���3�
hlSvBZ7
��2G%NL����o���ZI���3E\=��U߽<�������Q��>�,ۜ4yN��at�U�K�Q�)�K�;�O���Z��Z�v6YD����22f����ia��3�?���	��;WgP�~�9`�0jޅZL�h�OV�X�q}��12��b���L,��yl��߽�be(WRL���[H�kC�4�%R��o�4���=���_�i���?)g��s�4�����ǩZ�dGtMf�x��\�����J{����k�^6j$�q�8<��Z}��O+h<8�����C��h�L�����A���F�k:�\YeX3�rl�(���|5��9g�Ak��c�T{q\O���<��Yp��R�����n�˞�76Bܼ���+s�6�Imk!�E̻���%��D�|Z�M7�Z�]ڌ~IAW��g�5�~����"O&��m*`����*�nx����*y���?�w�Q�%�c��g���8H�w^��6L��nh�U
�Xx�c��F�X��9�ېEt�4N�1`��,�'��)6�a���e_�j���lx�s%�2�f��Ő?�O�Z1$VB�As?w�e�u/���f�4%�z������/8���)^�����^6�ݦ�8�	ǪlN�w�h���4d9ʿ��k$�q!�����N�؄��	�G:�\t�Z�z[o�'��Y�^���5a��"*�ٻP�{��>gH
f8?�G���ᜎ��-!*4H�|��~n�6*�&�/��nH�Q�~,�-� 齼��\`1��������\�U"~E��������{[W�(��K�M��d����K�ڍnk�l��$E�*��Uf�����~K����z�M�OF�"�ݯT�>z��9 �2���}L�Մ�n���S��#��b�����x��1}�k��t�����f���/\��;�$�?!462��,%Q���4U���G'b�,���e,�_#�����(�2Ⲝ�������l��_�8���Л`k�0��6ASV���p��v�@�|�X�Q��	��!�Q���1]��n���f�[��F�Ұqe��\+��4|/ѹF�A(c4��2�h�V�r�Z�'	��f�X�|N��vi�ֹj�a�W���������Gv5��g��X"m!��5����Ԝt����L�i���w�lFީ]im�Q5�I��߄��������F��*x�6�e�Д/�2�����jp�7b(?�|B��p��d�����I"u(1� 5���O:�:��uߍ�u�	�Ѩd΢s~E�<%���v
�a���I���mfog�aw��M6>-�p$���`�s,;��,`�ԃ~���Rh�h�#����B���r;>��ߝv�5�*��8P�����L��E���6H_Mͩ{�ОZ��b[H��xHvN̳ф��mV�-���td�>&����>ƣ��nܓ�ض��=���9�g��@�8��V
�XO(��� ���`��mF����gD!t�k"c�w�ጒJ���,f�$��d1�z�q���o����*�N JAWZ�;��� �����eO�����8%�\G'F�܋��v&������=l���0^�w@�*e�(�W���H9�I�����U9�g�d�`�>�͆�*�)^��2 _%��9�e5g.Dz$J�+����_S���"�b�׏cU�U�a9�~�t���F�l��|�#q��4L��M����9���+
�i6����̴S��$�H�����.:��nƖ�0|:g�է� ���/��I�i�{�83�o��I9m}�Z��s`7U�6!���Hh��eÌ�%,���0�{}a�2\�p�*��I�����S_��!�	5�B4]���PZ��JX����,S��Y��-Z\]>/���uI����J\���?�n�3"8Ć�=��ٽrѨ���i�XocKT�i�"�!����y���չ��ZC��ͨ��:˕�m�֚F.[N�$Q��9��2s�!�=p�$��P��%v����i�Х���p�PB�ͭ��tl?��n)tÙƂ��@��2��.���|"���pcu�s�=��R���s�+IpŹ�%�q�c�t����8=�Hp�1>2w��h;t�� �� $!~���sg���;�,���;��G��g�դ}�<hrh񖰊�{\��08P�<�!���3Iˬ���8�2�0�e�q��.�K�Yz�S�kzb0�6N����N�P#��^�P�C�t��P@��Q��l��JVNj�|I����>75]e�as�("nȕq�-D7�P6�7��%
^�b<� ]Ǣ�Or��~%�ԍ���RѬU"�(]����?��B	5=��
�]��i#N]"�1��d'7��^�װ�\,����/6fò�Ku�% �u�pod'e��+��=�Az/���=K�4�7Ѫh���֛	�[��ʉ�㑇Y��(�s`<�����Z@�����l��T��'�����w�N0��#E_+QE��,���<QC�8���+N�����]��M\8V�j+��I�K�FhUX�i��Vu$����I�X�sB\���0�܉7c�S��V��R��j��>� �¾�������w�7���O��N����Wu)��S��zF�#A��	0m�v�C�)W��ᘪm���&�p�/z06��u����������(��d���a�e�Y��q�Z)����CR'�I��@<�p�U��`\�{�!>__�~ջ=|.�y�]l��Y��[�7�)��!`�f��G�OŎп��ҞV���,ʱ�쯄�C՜����T�w�� &]��[G55/*�9���ʪ:㡺�X^�u��� -�ӴԚ^x±4��	-3[�t��3P�yı@��:*�ΰO���鳲&J������5W�N�+�ժ��|Y����\���z�f�,��1�"D����{5lEp��6㐬h�q�DN.=��9l')_~���]�NB[�P��WfꋖUs�ٝFt�3��B�����TEe�<鰼z���5P��b�,�x��D�'� ����Z���8�~�]��wa)?T�?/����Cָ�C��ͳ���&HQr�����Ȁ�16����9$K�Ři�ب���uQ��V09lج_ç<��Մ)�,)D��x���w���"�VA�S��9�_�����i��G%�ޥ�H%[:)�!G���,`k ��t&(�6<�k�)!�j4-e�;�<�� qA�����0J����� �j��+��r���=d��F7��0�_��ۗ���#��in���`�T��O��5W[.{�(P	DO�j��>ˡ���8���t�Xyy028��U���#̨5*�e�q
4�X�� ��TY��T��Vq��O�t�o�ӋJR�Ȝ(���Y��<ޔJ 3 �K򡙢ҢK�ӍL������b�$uVB��i4�$Tmvs�$���M�F��y(����Yy�q��W��'f�Ћ)�~q��va�҂4�!�@��O���/8���_�~c��(I��׭E}@^�t#k�Qn�p�:���cH��4r<��ͭxT�d��D�2'o$��:���,��+���72y�W/�M\]�}Jj��'�,����E)��'2O�9��6�!b�셩�>H�e0��p^�.P��%�m�
�)��K�i7��)�GiL $	vju������2	�2Fc	��#��!�@c�r��K_Ύ��,
����1���̵���6�7/l�o��ylH�����f��kO:�[$�3���.��r����^T��Jl@��,C�'�~�B�5u[=�=���_r��oa���!��;��ࢱSqMΞ��в�Հ�2v�D��6�"�����t�h�p�� �cMnX3�r1ud�v�ִH<�.��.ɶW���p��j�E���k�onh]>a��{����UM��m#��ka���_��{2��qL�͵PV�dQ5#ݜvm�|�ЂH��QB/��S�J�Q@�ŐhWvp�H�(��}�Ik!��(��ajS�g)8{�.�]>Jі�Ú���ծ��B��:Bn�Z$�|�����.(g�v_!#��9��h#���b�1������$�o(,[��^-�!N�l��i��X�����lA�R� c�����itA3�ZAO����Ο�����=���g���ʗx�������(s&nb��l�(ٚ%�$�v^�}db�~�'�o2<F[��*���7����}G�vE�
�(ĭyfص�o�����n�� �����Ӫ;s�O���Vb���E���|�� �Ǌ|I	��T�T��m[� ,�V*�S�t4�̢�E�KN�[`*lɵ�ts�ϖ�O�l���wF0p����3¦ �?U�ceI9)��
 �W`v��`�̴������f����'���KlF�G�w;>��r�L6Ui�k�[�:R�R�)D�7��'��|E8��R]�yݤ�Cۖ�]l���O�\<�O��ǟ�g��(��	p�k�/���V-�)�Ў #Ak�/��r&? O���6mzp���N�I�,��0y�p�-9�6��$�a� �t6��@q�H=�c��-PtiR�e���B��;.�qk�N�6E�/��
e�č��P�kb�����>��!����g߁[�s�njO �F���JIކ�^^rO(��NAB�^���*:�_Y!x&M|�0��� �ŀ����5%�����Gkuj��X�e�� �	C;X��<��?ܛ˴�́��N���H�sǡ��b��O�`��&�q���`'�-��+�i���R��I��`�{z���=��cm&�l�4��!j�=������ȱ�i��V���k�l�}��g\��[_|�I�USl�/>JY唣��˕��׉[��.��� ���ހy��I�d���0�6Q˘��� �_t��lu��L~���;hθ�f�0��[d¾
���`k�e�,Z��1׹�,��9t9�/<P���b3��og؉w��y��tIS�|�J�q:}�E��ľ �6�ܪ���b%���RhJ�-�K�cE��h�?��LΉ��������W�(\���;�r=��!bN�D�w�`
 ���
#Y�L$^5X=5��We���	F��S�0P� �2�EpW��<>�s��*��M�:�l�W�=wW�*�Ǘ	+K#��{��)�6�2��Nf7�� ')�ɚ�����������G
ִTc>>�P�Y��gJ��h�h(��Δ�g�7�j�8׫�r"�a�\D�[�d�'��gEL��9��4l��#�0
lD��T�ڨe5��ѯ��-鏨P��`�9M~��ى�~Xu`���}1[��L8��-�y�WP���n��-(��tK��b��SJ�����"�f����l�K}$������ōn�;��j���p�A��ʀ��}8���>��,q�B�X���!�$c�jQ�G؆$����o^���WX��?W�^Z�T���ϵ���"7B1��	#�!㲖hRڪB����'a��,HL��YL_��D�5�l���?�#H8K"���^�1CRdVJu^+�mSM*�$��9X|ܸm�߯5��#�T���ns��`�X�mӒO$���*�$7�jM�J�80Z"��]�G	N��#Wr`���B�,.���ڭ�Д�D��Bou�t��;�[��=��8oT�{m/"�;�X������6��Vf]�Mi��,����!r�����z��W��>s������,�G�����g�3��=K<���2����c`)�J��Sx��KV6��._��z���o*L��B�����3	�	�Ӌ�.S�����y��{��Q4�Y��[ڌ����KM�ŵv&J�&���K�S)Z���dw �"��u$l�K�$�P�4~J(�Om;�����:Ъ/�S�o��u��W$,�}\1e�f����3�)�C�d���Ah�9!*>̫��n�T~q�����[������B���,�AC[���ƫo�$v����MM����N�#6�=k�Ƙ]�MR�F|����&ha����⨙6oT��R�Vi*��w�H�����'/���dMrm7�߮�� ��@����Fb�A�$�8!�u"۲%��B�OM{ GԄ���WJaC�v�?��ʐW��[R�G����P��@&�̄k�N��x�w���!Ҡ�&w���+��o7�_���~8��z��vI��0a���i!l;���G'{S]1�k=X�O�\lVi����1oM�>��QHl��64F�\���5�a�ֹD4&O�B2u�uب[i@n��U~,���c\!�	�g���5�ǋ9��Z'RH"��K�ZQ����IU`.��P��n���'���͎ȝ�n@���<�%�ZXp����o��"&�[�<���G��i��u��A׎c�t|���Q �%ޭ�^�|� _��ć���y�<���]*����/n�_� �����qd�ap�%�K�:�j����&���V��72{7��S�1����bb����("�pJ�����̇2�¦O�	���_���~��0&���Ɩֱ�@$���ұZ�Ma�^=�+�4��4��hdˊ���;�6�N��q<��q9.!���'1f����\�(���c�npb�RE�Mg�~y���{o����oUM�u�\ɦ������Š�6&S�0����e�9��9$љ�UP"�����wI_��6q�#���=��_1��rB���<��p��ף���C'���9��P��t"plﱇ�B� �g�=0-¦��V
i�(�d�}�R�Oh�������;���O�����B���&�|��+N�b-��C5�DtI������=��vX�-v{�(x̌܉�a%�0w9@��-��J�=7�*EӾrAg!=�ZKV\��c��0
:1��9ę�j��Ԟ7j��p�6l�G)��װXؑt�Vwz�E�ԙ��8IO�8���s����+����2��hLJ�?�H��V�ġ��c���H�^��jV��L_j���\�J���)� |㌹��U�!��"|��	�4��6�1�����������p� ���3�C�v�3�>�g�N^Ú�赓P�������2���n~6���~f�^�?��M�Μ�p����'s�~�,��W����	f3C�"��o���7�G���V$����P$�ș���o�W+�WA���
Ǎ�����|y��t������x��Н��϶DwS��1Y�|T7��'�y9/��9��\�y"I�Ww��Ph�	ˌ]�樲�l8拗-� ��m�~�z���c�z-�bΤ��k�q�q��5)�T�q�ɘ�D������*�Ü���E�hik�??�|��V��'k�gJ"�L��C��-���%F*|�Ćܾn�85�!���LW��m���]b��w���s%��P6aۢ�P�k�-�Uk�}�ʇm����gZ�;(\�3� (8�&$`��r����pA�>@���Z\"3�6��2��j1c�|��R�e�u	=� ZHu]�֠���<���炯���P�И'ʤ��Ա����u��R�����Zn̋h�Twt^�L�l�l�X�� ����"���!$h~�!eR�=�`<����Ut3Q=�u��}T�?��~w�5�?��˘��Q�t%R�w<��	k���
k��}���.�.!̗4����6��')yz��-U�y����u׉�i��"��nb�V6l��GUW�hT�K�h�>&��R��s(�Q֙#��� R�t�M`��x�g����~�f�y����H��t�!�-�LE���
�L��/`�@\an��������9m]0l�a���4�@.�d�¨F,7u�73�����7���EbX��ϓ��[m���೻aT���p+rA�2-�%��@�BF��F�/%��z>�#�) M���)78�䁗����
�d�_i��-=�g�]�YOs�r%
w�s3�,?k�B�+�f�1��
��?����>�Vy�X0�=�������B5'*��n!�Ѕ��C��!4����������}2R�Q��Zc� �{�����i���_�	+�VW˻tv���a�o	ÿgvn�!b���5��J�Js>ӄ����o�L�|_(!J�pa�_���r�:�9�g��������1�ѷ�4eRƠYh�04���Y_�<m6ћ�7�-��GW�~����=���K��������\t�$Y�E�`��10��ves�}J��sL��L�!��;����};���K�e�o��J��75��ő*e�_�>�ia�$mq�I�=�~PW
:���T���q��$�Dx�҇+�B��}�Iݑ+-����I�j�%������h�ID�'��x�5��
�Tu{\�t�^y���~AE<�n5��@al�>��0,bw�NKD'c��������r�,B�nl��r�Q)�D6��(�vK ��!����Y����!jO�L�UJ��*�<���P�FG�Ʈ���ٕp��-ok�=P���U	ɵ0�~	y�>(��b{N������}�:)APIj��Mg�*#[�q��n�\��#���Y*�a[��eh�H����S 4�����\:ѷ'���u*�B���@7C{���{��|��߄���g]�i��@h���#.�W��e���KX�>@lX��@�����^��Xu�N���`�Ѩ�B�7PR���Wl����g�7h>Lr`��������.ڔ��k0�64C��Z�����m~9�~�1�F��u��L`��H�Ry���,��9]WT�l_�F���wH�ʯ�Pu�[�쫄v �"�{���F�R�xYay��^��ٰ��)�C�V����<1�w��/���¢��/��������0��������A�6���q=(�Ʊє���ϻ�`�p�0ó���5AC����&ɳ�v-N �wҺ�M^�D�����a���;q�c�JW+jӋ�R5�e� X�U�]�hZ%&�
*Jms~���I���?α�er��m��D�Q��_e�J��������0����R�4��𐎳�����RFݬ@�����'H^��qj�����נ67�ɫ��at�P�o�ߌ���z�=��rÒ]�>�M{�*�H/�xu�2d	=v���_�ߍ��i�x���\�]���I0���8�I��6��t}F��-�V�*�8$裾۔�`����	bO;���^�)��0K�W�B�M�b�G,�G�A���B+5���d����ĲA�#p��/�����:Bn����	�� L��[�A,|>�Tԓ��bj�1wX0B"���ڐ��~HQl���@fL���h�Y��~����!�PofxI'=��3������X��y�n�N�帑D�������.� ԣn�3+G��EGҎ�ʠ��^O}�P�k!�	�<ūj5d\����m)|kH��.J����e�%��,b%?)���E��p_e�Ѵ������qs�	luH�X�}�v�F��C�%��ؖ=Ϧ��t�-l����P���6&@:=ԙ�l�A.Yk�J1���u�B��g�{����iR5���y5\�,L���ƛ<�p��?<���Fx@��gZÞ��
������`�M�s�R�{���
c]��=�'���e�D���_8?dl�-�f��}��b�����%����_���mRhk%'�HO�A���ij�dw4���9ϼEG>boW�G$��;� Z�S�{xώ��'<Fi�r�b��[
δ������[�Uq R������T#�{�C�Q�y�xi���D�����$öֈ��UZ8���ř���1{�O�쨾�T�[�������:H�cޚ2�lg����j4�x�03W7l w��5C��1�yAQε���|�X]Z�s��3��Ef�<"���3i)"�jƏ�2��6:a�0ω|<�('�/~;�1�PJP��f��o�VH}�7��Z�l���K>MI8����䑯!7��?yH��4⋀�CGo��B���7������Ԍ�S�q�g!�Nl.  ��E��_Kx�!��l������gB�P\��Q�ETGֆ�r.]ꏯ�'Z^�{��"$�9�%k�h�����=D�P�"0���6���0��#�T1� ѥ{��i}+&�����m�&���<J����S���W	C)4�H��*��s�_'2D ���\�?,\Z=�I�"|��ptx��݁Qi���0�rtZ�9����qMJ�BR���s~�&|�c�:�0@�R疁F@��{��$�������۫U�6���%z��Z �6.N!H�T��|%�n��9�e�=�\��ښ��D0�r���-i�\/�+H�}���l�7�x���t�{G@�ҶJ��e2EK�&�jgI���_#dcD1:�(3E0[�ܺ́
��3����ގ{�~�P+��Q��x5�N?*T��:KޞBY{x-9�?�pD��e��tz��L�rcȺ��<���}��lG(M$HO�ƣLQ�گ)��d�-5��{����S2�E�{�%d�뻃=�,���;v�.�4/P8�n��sX~�;2'����W��N����zw��N�[������3�5f� ��`R5&D"b�P��tdv��a��a���'��׬˕���[! ��<���:~h'�|�w꽪�h������{�:�� �m��Z��D0�	0q(N%/��Tڀ�%�?��I�,E~fb%�pA]�����Zج~���{8*����"��7躒���ϕ�ϮsX��b� �A���0�y2���R��y�㍬�O/H����R�tʂ�l��2�A�������
��{]3���@�=�(5g��A8H�5�;��O/��u�`��PUӊUh��!=��VݴM>�b7h������k BZ����4�3�`6ƅ)c���.��1������y��蠊���J�I���av�NZc7k��i9��(��:�Q�	��P��N��EYZ�T5m�ٰ:�z 
Ђ���������tP�;��_#����l��F	SU��R����dK%����N�3{�Yp�����f���j���;Q�=!7񳩵��f��#
I�s�����!S���Z`�f�H�����ܛF���R�����e�'<k(j	�+�k����������F������`�UrH�4�G�-�B�zK�	<.�&J5�5E�$½YMd�Q���)��\��E�/ �=Ѭ*௿�e��$�	�#ב��Ā���MI�L�����"�t��:�a0,@fg.����e&�E,A8)Cd���U�ٜE�c$��� c�-$�=������';jK87�l�,Ɵd�gt��j��iO}x���2m�����aaQ��͝�9 ��.�$�֑WL�ҁ�o�r�i�w�.�����ݕQP��T�y���� �/���r��e����!X��0����b�ȍ�)�Q��}	��Y�p��Ye�r��!3iަ4�=���{�F�n	�r�N�#�����u�ȕ[_�Nj�o�YFl�q�b��iT�;�jr�6��S���N��@�٪/��@p�Y���m�]�e���V����1M�B`]q�Γk��tMa��GњwM�s�% }Ѽ2j��C^d��t�b�?CS�X5�w��G�F�3���RG	���|%|��ehΝ`M�`��`���Nzi"�����&�_R��+-�t$����e�d�>]��˝5���7D��7��M�O����yp"*-�S�g��.,��n[s�Җ���9���Dc�~"
��g2EwB�8�('p�G������0��!��p/��G�-��[ڧ�W���Waȏk�r�ӳ���	�ڹ��#qQ��m�.�|��i�J�,?E5J�5�^Mm���ά]c����j��T^K����h{��agE��Ģe�6����8,���nS�7/����.Y:��L��.+�Iu��� 5���B��"�#e���'���t�zq��| ���KÈg���1�M�
y^1/
0&����JV U��ג�q!�����T��l�s&�:d)[Zd�Yh�R�,���=BdPq&BA�vM�q��kAk�3��{B�I��(	n=� �SJG�t���<$ rM}�~O��h�T��QK�8�&%�F����i�S�"�)�t��f����`��J����۵Ľuh�E�uز����Ut*ʭ�YHeI
��ͼ�� ��X<ǻ)�*�>X�F�Ƙ(��/s~�IT0�7��|���Z�Q�8:#t=m��
jLa��$�&����ڢ�/��E@-�r\�e����*Dm2�7��u��L���1��ܔɺ5 ��i�b3.�� �g�,G�|'�R��xV�<�����q�x��yQ�����Yr�����p�9E�Y���\����Z�A�`�&�Z�k0<I-p�����no/����F�~�]�j<[��F�)���w�r�z�.�#_L�&��W�$\�mۅ^Q	��q�y�L�g
�:�XW�I=�)�T��	V�����[n�j?����A&з�]W�X�;��������-4�e�ő����6HX�H���5��� F��z]4��˧-�ګv?>�a٨�oS��ʭt02;����"
ߴ5���+"bT��.�b����"#-�4�n���V*�QF#0aZr��;�)�o�k��3o�J��Q�{R&�i�:�:�%�<!}b �	l�`��ȅ�x-mL��b�B��	1�h8�R�--:m�u�R� o�*�:��g�Q�$o-[F����s֜����o\3ؘ.��*�y����I��LK�a�?1���"ă��=VPH�{�y�#đ�e
+#�sp����7c�����T
'�Ψ5=�����wp)��y�m�����n���C�K�[��� \r�>��Y	�y������0ʇ�3�IQ[3y�K�X���,�#�+4���l����TT:w{����%����s���<ZN�r|�=Ѡ�VlPe��W­����M�9߲N0=е��.hֻ��TѦ�ɺH�f������5���g��\�GYՠ�F	e�q4g�L	�=DS����T��)�����a��� �^����N��*�_{!�&���B�cdV�Ν��*e��Wd�)��:��jt?�|���Y�>Ӛ��C�c(�!�Ԅ6A1�M���zCH��[P�v����E��ת2��^N��mj�b.J`�<�O���W���֠g{D�Z�e���l]�v�.�ZH����J �V�.1hR[����H	���9e2��%������^&�ZZ~�өl?�'��Kf=t�,�t������v���M�[���?��쮆/س����;%g��K�*���˽wLu��#UӇ� ��ј�Fl&2LXhA�k|U��oX�0�o� �ݪ�o�-�������HG� ]�z�q�E74�QnU(Y�z��D�Y�|B�lѰ�n�I�@����<��Ј��Vv�v�2ׇ��ʳ��������h��v����ф�}Zi���0��1�@ Z�{Z��B{׬�8�m�A�j[gIH���lT���s������,[�`��RR�I=]�����������w�_���k�ē'��b��ك�D����f�JȴB���&�2��E~Bh���R�·`�W�J,q�[N£0�"(�U��1eka_��^q�9�C��yo�Mq��aR�+��-�Y*��&�7��ݤ��C�	d�6�,�d><�cG��m�Q�$|��4��;[���HI���VS�$�����l���]����?�ƔX�*X��5khafS�{0��wQ���0ײ���d�����ї�A0�/`J?da�> `���/ ��"�{O��p�8��9*��� � .���1���͓hb�1t��L�mj�S�b���ɚ���M*F�;\�C�:��������ψ�'��2�����9'�_f�o/S�Ki9�k,{��l�W[WW
&K����g�\k$��.oBf'�;����&����_�����$~�mD���*E9��񸮖��R���#�N������o�\<��Ѵ���)?��/�{��-8O�����~��|���<^db4�1T�S(�1��P����I!�Ls����`6�c���� �L�;!��Жnȧo���� �$�zA��x��3�n�Ǩ��i�N��"ʽ��|�no��o~�D�u�	��O:�e,�/�t1����Ɵm3>�i�ɋJ��8ॳѿ�@q�p�K�ra�'YD�R�����UWe�ѓ���C4tp��sA��cl�H+��ҵ�Ui}�9�N��31����eR�bj+��i�.��z����	���lNe��"�r�6ۇ�XZ�qh��o���Non�����c�Bd����:N�#4�.h�QޑSΞ���4o6A���L꠬�?�_Z tp�v�x����ک�!eWk��z����B�:p3����-�\c�����ȹ+jJ��v�q�ܲq��X�`e]>C����(�e��9�xh�	�&!��� Yc��x�	 u����Xf��=�� su���i٬���Z�c�+�E�F�K�m�뎶^Tw2�(�G
�6�/�uۣ���%�1���Xh��8K{��j�=�%��J�1�s(_]dx|�;�)�H��j4A����.Y�;NO�I�����V!��F��3%dU-��;���K���0�p����_���
L��l:�u_5���[�D����U��{";�~�A|�/vz#��_�!����n�E��k���eT�A������� �d9��K-C��y݉��k��b�z�%�Q�GU���Tm��<���b��o.��f1ֈ��w�s����u���q�Ť�_�Q�	�/$�����C3�]%�貜�-_-��O2"%�.
����z-��X��I�D[^���b��7� ���g�\i<a��"$%ފ�p=�3��G�Y���:���Մg)�wk�i@r?��g+i8��=�,"͞ڿ䞕��۝���mG Q���/=��0��y�0�+�/z}=�5���ħ
ϳJ�7���+��7)�'D�!��-��%�{��Qqv��$g���\ӥl)H���PUQt��rU %���W?�_��^��\4fX�p����mXb��H(bP���c�����2�I� ���΄�wƯ�Dfq+���P�M���e�����'�I��X�H�)*v����f����]�0�7�_(N�t�P�V���R�B�;KH��=�Պ>$�u�<\V���x�q���w��K�Z�Q�C%���c�D{�
P��ch��Ɓ8k�v~J�(4���u��!d�A��/	��P�!���c<�Oi��?^�E��\3P��� ��'��6���n>��gk�]H�GK��GG0�Lh�ssԀf�wP�c�Dkfg����l��X�Z��({x���fJ�BrfM�agx8- -G;���[mI�`������(��.��L!��s��� �'(�5q(��G�Zx�H�G�ڐ�pm�f2�K�7��in���S�G�'z��ۦ�?�}�}"�;c�*����,ao��^E�r�&�5��|�2�����En���) ]
���0�.�k��aF\BN��E8F@s��~#a��m��sӏ�n�v<��1zD�֖�����|^ �W��-��V�Ӽi�ɫ�M]-^-�j�ht�aA�'~��v���8�zd���K@z�5�.������b��F�V�E�#[x��$c^ayt�s��^����M�_�Y(�¤�P��{�5�S?*����Ɗ���?��E{�<?6��G%
���l�ԩ��l�\X�b��JjA��P�iɀ!�J	�C��[��&��[�T�8�ăF{K8����F)����z�Np��JRb���|^��xG}i&�U6�I,�����w�/Dە��.�l�)5V{��J��@Z8(��?�L�)�,/�J3}g���{�;itޣr���}�v�,c۽SɊ�J�,��xZ':ҺY	q�0��U��P"��ٚ^Q.sW�Yf(�w�]�R8`a�29�S2����Rۧ�6b�D�D�H����m�s����!?z�~�bG%��Qb։U.I��ps�rg'
*�4.IM���y������yB�F1�f s/IO��¤���v�;����4@�|�(Z\ɬQ�l�?K���S=}(�yն�D�����o�@���t��vM�O�?���d*Z`�U�[X��9ܹ�f��k�%ER��R����َ%���]������NL�_̷�� �G�';70	#2����J%���V[Q�Y��l���� ���е�d���5�>xҦ�MW��A�/���m�����Ƈ�xd�kg�du�V�[MioTǋY��L��Lg�㷵��f�R���_θ0�j�P0�-��o��#�@�c��d���Q�2�1�B �D�ӕ��Jq�1��,�� S
%�a �KF/qEqƣ�����×���R[F�Y v��4�XB1U֥� #QY��B (�*��%d���ht0/�˷{��"��e]_�7�d��t���	w<���_H��<�@r̮�U�?���a�:�@���>J�x�Z�$��*�I�~:���!���� �(��tI5VK�o�ϦT��V���$�==��UG�������?;��I��m�V�〈�%,808��]t��Gs,~5_����� z_�n֓O5���3`�)6_�K��0��wn|�T�T���~�9+q��,�ѭ���OC+�Ԯ��pyې�2��<��3�^ �;�e}qr�~ؤ��ܔc�{�Q*�2�y��@7�Y�OHԕDd����g���Qz�s���Oa��}[�T�C���3��~LO@)�2W�'a�pU�T�b��\ ��x!'v�ƀ�@�`���0m-0����u��1� ��p�E��z9Z��$����|�B�)�<��SPʮt��B��gG:N:�ug��#Py�D���_�סDW\_Rlga���9�5���2Ic��L�\����.�a�'q킁d���<R	5鳀���hd/�5�x�=z�,��{-,�NI�.�OW���x�c#ȸzՍ�?��@ި�5]���` *��GO�<�~��=�1`��ێ#����a�\'칺j3F�A�K%��љ��֑@1�b�j:�Qc��T~�\mqe�:���yC\�>Ŭ�'>t S���4?�*�(�T�����Z-��A��g�mX,Hݾ��p�9�+���~���E;y�񧎍��X�V'Q�/�n*ۥͫ�T*�\�G(Q�L0�s�����_���U_�Oy�Xfu֤��'x.znp����be����;�����g�	y���=��te�ى|���7���:~�2�x~�l�ڈ(�Bgv�6�I���f��MZ�#o�h����S�k�7�䒻c��U�lr[���?�����?����>R�D�At��eWʶ�X�Le�IEh�3����r��X�W[�?���Kƽ�:�w�ǃ�&'��{�m��i�Q�@�!q�bSު���e;#�
"���xμv=�k�]�U#�ŕ�_NJ�agy��,ʙ�o7%�!�Ù�8��Z`� +V��q�)�S��k<2%*��'���ݾ�[�S���+Uˏ��wnN�A��^��g�
��]��W�Y�z�^��� %��$N��+�-ڻ.'����"�0�([W���?��5��?��׮��^�k	��Z���>�H�-�۲3�9M��#�x���dpvG���2��P��@&��69'�h��Ѱ}��Y��EW�h���4;�g:M��>��"��N��;��F<r`��6��}�*�E���jT�R�0��%iy�LY�W>ҿR%mOPH��㰄���!�����Z^��XŔA.a�V���"j{��ə�E��!5���ɔx��x�V�o��Qx�x���VL:����1v�sm���᪇<���0�-��m���a���)�����}�J��<~�rI��Ic��l��%����i����x$�CW�n��D�a^����|�A�M�E����II��d��X˂��qYsp�9N	K
�b�5x�=ս�+��l~Y��S�Y�}�8��R%�
z�����ٓ2��&t�+5�&���Z#侂�܂fֺ���.�nQ� �ۺ�-<)] x;�' 2)�,���:�m0�����,]��"@���0K�7jn(^������:E�yaV�7\r\�A�����A�5�FO� ���	������ͱ�^ԸTDP�����ΐ�!b��F�F��ޑ-Ɂ���,��}��Є��,������?Ac��g���,$ţ�ob�j�M;3�A�Dd݀l�������F��Ƀ&�A zg�I�bf�Å(��+Z4�ΞO-�[mo.��IY�*`�)�������N�L$�	�����vEJ�Ffa�s�z*h��U>Y�2�d���~dˢQ֤��a�9��)���n����rzy�����|�k{�YY�hm��-.��?8�RJ��f��BE߿��b�v���J��Y~=��}A���X|� Ru��ѦqJ�fe0����9�=���y������*�56��|m�5���u/G��.a���vQ%,TK�Z�!�k4���,n7ÿ��L$�*�hDf��m�
�.�-��Rr��?:>����-PR���tf�i���t�B��=ux��Q�OB�YkҰm�VS�ApS��ie��h5]T���� ��?������������>��-{�;]ϙ˧�1"�{�%97����S;�6��g��&�qH�Q��Hf�-O�X�t�{�:$����/��ƀ �n\'��S&L��
�q�A��ѫ������ۺ�>�>��5�nblkb`h �D�K��*�Ϲ;�͒b�q�0�i%zgzB���C�9/K\���!�Uh�t?��P���eI_`F`F�[�6љ� ��#6^n07~����"�#�����,!XM;�_��������q���~���0�B¢�@��6�"	UD.#'Q�UAp�R<��PJ��W�|Dz�w�ٮ�Vo#Ш�7g[�Y|�y ��3,�L��a�A�ن2��w&e�9%�:h���$�C��	Ұ3q�۝m�M���,f�vl�tf]�d/56�*��O�#ke��(t����V�i�Eqkb��Q6/��/�>��wT��o�y���8O�44C��,7��K�@���q�B�H��`Vݛ��9�P�����e�E}A�ba�n�[y���>�&ȸc?e.�:$S�����O5��'-�;������(�¤��j��i�;B|�>��I�� ]��7�*L�B�ư1�����`"g�m��̂eĴ��Li�A����F��C���A�	7N(�Z�h6Ɓ��<2��n��R��BU��0�]2�^@E���'��F��� ��?���d�8�E�2n���&%>Fr�#���}Ԫ�А�-���籅i_��Ë!�h2dl�J4��|��TBS��;��qT�u�=��D8U	D��=���f��j {�ٰ��3bG�e�
�}�㘤�W�줚K�8�n���\�x��˔���Ӣ0nh!�4�?ZBu��D|[ft���%l���H]�&*�%l�#�'�b7S;�뒄	�H�������z�ڸ��Z`u`���"�ԀN½t72�I�Rk 8������c�iv��n�>�9����U��G��T�S�=1?�}HIc�f�B2/�l"b�Wf�1aqd�l}������-��*n(���^T�7	�"����T��s�_�o����p���-3t��8_�����UB�{ ��.~��.�e�3���O�ŖHA���@��9�ա0�Jt���O�*pm@�i0���N��Y胬"xj������3����^���#����Ş	fX�k8K�e�tc�T����KH=�e� �	PӐ$=�R�Ֆ�]k"�'$^0��"�L쪣^Ź�R�E�ǫ��4P���(4(���Ko%�B�e�`���%�)}f�#>�`J��Y׬@���۠�.lf骄v<v����ص5�p���!�g�Efo���%nQS��Z�{&#$Tq�evً,wҫ��v&o _�&��q���:s�Ii���:Fv`P�ؓB���n��35�>��<�]��:V�@��
����S��E�/�p�U�����]��2��ҪM�:g�Ov,���{��������d��D��y�ŕ��6N�j��y�S���`�3h*�H�'����'�Z��%�h���n��i8$�������P�3f�\)BYF��+H��oǢ��OǷUI�����_����Ց�7���S2���`i)��轲ۇ��fIx��z��/�Y�uJ���eFU7ˢ~+.�	�}H��xO�
|f�Dh��K��Kɢ��}|C��-߰YJ,�l��ӆ� X|���;
�R���^���D�����8 /3|�jn�mI��Q��/��u�r�s\�>q�Pa�2
���zJ��K�ߊ@H��d�-���O��?�0�0S���������o���L�,��`|�q,�@}�?� ?LN����@����ve�����X�nA�i���d�Q�	;+i|M�Ҭ�g[�ʸN�aE~���9�����-�����r�
�r�$�)�p��8(6#�<n��0�QղJ7dK��<u]e^I3�ќpOlၥ��{� (�S�7�����5�̣žx�{;FX �g��Ah��,��dY�\���lV���HL";%a�v~ު�_b�!�/O�� 7�{�B����b�Z�j��	r^;���a(
W�_�jE�#7�`������e(Q����:{��`S�3 r�H�DO� ��@�s]�(��6Y��P�02�w庹���]"�ҏ�����5�x8��h��u��uMr�3`U���1�����B�3����#F��`�>�7+pq8ܧ� ��~�'\�_Q���^�s�� C��ͩB��A���� D���^����ْ J�b��՝��FK�i���,�N窱�;c�{n����.ExCT��+��:9X�5���������T��_rB�T�/X�Q��/�_V*7��D��nZ�Wd�6ޓd�Į E�բ�;����IHZ���B�SQ���}Z��ABN�)m�U~�C'���Rh�e�B׋]�;�Y�/��h�;Ex�Cʀ���HѦ��:�}A⣵l�<�f���PY��8=�Y�n�ZT"��z�D��~4�^Ib��X��_j(���YX��$��5�q�9��O;Gs�c�x���A͔&]|����;�8l���@v�
�~��#��VBi��
�U�e�4d�h/���&��W
��ĜԊ�n�Ď4p���ʹ�px-2/�	 S�^�9���<���V=�.d��2WL��$���N�e�]�T��:��&��ǟ� c6K��߉�Ȟ�ؿ�?]����hOǾ�F�LIǑEס��z����Ą��ڸ:+˹�J�t������i5��a�/�aVx�,@�Nz5�J�_�#�ܷ�/%�!��:���|�G_`C�u������M����G@����~;.��=^4<AW�g��4��<%XT��xJV'��X3���Ec�%�l4,���U����5��@�D9
�}m�+�Z@��7^�x�3�޾CU�b���}���k)���>�"�T����q�WAmC`<����G���H=������q_��g�X"�^����"N��颚��?ZK�l�qm�yQ<G�����B�h���0�O����f��D�J������/h��f��B�q zŋ8�l��;�oEMFa�9��n�_S�Ռ?qF��ԭ�8�%{Ԉ�����
4I�z��향-A����wo�?&WQ���Ŝ"7CVR�v��Q}�Y*S��ZK��O��(g� �O�ठ��֘��{��V�g@�G��M����@%�+���AN�	'��g��N�l@~ԝ�y֠�#�*��٦*��C��HO�}<Ed�\�Rw���w�8~d�ߵo�|`NM#W��u���V�R��d5+��U�(\� �޺M+F��1z�3j�v8B�Ĳ&c`j�i���#��N�MQ�"Ì#	�����l��;����y�-�h��ǐ�c]3���'�1���zA�
����?l0=��*$Z:���m� �Եo4�N���*YI-�Nɂ\�ڳqTa�_�L���̞))��
�J��R�h��2�R�3yA��z�0&��F�
q��%o"��	�
��V���������Y_m��IsS�A$�R�]l���C?���m�������؇�̾kA��"�=!*)�W��zSNkc��68PFo�=���#�W9ke[	�&���J��ZE�/z�`�\ {sc�g-H�[�D׾YW]�D�y_��mP��
L�	g�E
�Ҵ5c�U*��dvG�Mlh�7W��i��K�p�'Y�Q�v�ek.��5\��u��,�KM0��-_Uj�/B3�$kN��/��w�!x���T��J��9Z�X��$D%�}��	P�TvSkGҕl�����wW��pF
6��ۘ(�����m�rOp)*��7I��	\���g��#U�0�7gl�d����ǡ����G�U-�19k�I�MƲ^�䴄�����}v8��W>"�x�X�W�8��%?�����n��)hx�Cs/�k.*��1:��=z2�������@1h_�E��S���oy�
f�
���dߛ	ُ��[#�(a�Ax� B+j���.�q�r25�T�pc���b+�h� "c�nbG�����#�-s��!=푡�(����~�z�]�I�Z��|�4�A}v���������e	�� x��&R����""������P���q`�}��8���3������%wł?�j��CH�C�Jq]G�g�',«�-O4��JV.���Do��r^Q���Va�(�Q���S	?.	x�p�I�{v��Pq���������xw�>٥�� ��Jn�ahў�(���}o;��/V���`��A|w�%\�M��v-.!ˬ�02�M�q�{#z���ʏ�C��oGVʼ��kx@Z@�&`������5�����iR̓��)��O�茦�j�?����XJ�S@���<���6�F�U����b,��wf�Y�0���Yk�E�p^�����l�|��h
���lڿQ�C����mk���9���#�ںBB�"�[H�>�2%�ٲ�?�3^�쩘2�{K	�\�4}X|�9�
�@��a⺞cy�"U�p�w�`cPoPSs�tC��G��@~�%�P.u�x
TN-]si�,=�1u��,��ę7���G��=�{E7�㫢lE�
��DE�}d����]�u�i,[`��	F�yXi(���&k��a�U�@̕��cg#Q?B� ���s���*xl��o�"�Ү<J����J���?���H�N,0s����m0%3��x��B�ý1��U�e7�� ��=��ϼ4�؀�:�\����S��Z���HZ�3��G�J��&�X�*�ƅ(�h%���3v���]�������c|���-&?�fW
#JE6;쩥n�2�#����Ǹ������׶n y�r������|m��c�ubRl��u㶺Nm6s'1R{Bj�vs����4x2$�f���@Q��S���A�8��/��Ω-^��}o|��!_�ڑ�����E�UX�Vr� �.�N�8im�y^[(�CzS�E1nf���R���=:4{+�T�a�k(�Q3���%L�8ij���A�Q0��ǣ:g@*��Fn��J�A5��$�M�l6��e�'*���7�/^�(,Ey)kD���˲6�����@\~e��P?I(�T#
�&	���l�P�ވl�)�m`mG��bgʦ���'Hv��*]*~F��[ ����aQ���׫�$�Bi~�.���[������� ���I�j9t�`������&(�Gde9�J�I9Ó����>�?\��Í��DY$��w��h*\�\I\��l�?�U�Ɏ\��@jT1��H:QmOX�I���'�U�3��{�g㑩W�M�q�&��sk
7i��L����DJ���3N�x�� F�UE�����.Y�n���Z��a��V��j�A��4�;ݗ���A�WA6#��"��f|��u�4sdD���{��m<� :�����r�ř`��kr�K���&�̡yl'��&�.]*Fs5ݔE�@���>�����]�V�5,z۲�՟,�@^���ʆZx�Yk<�p�`bHI�G<2�}�Ds�>�!X62OzF �<a83�V����!�L\$N�t��<8�i}�S�r�"#�*>Ja�P�\��$�0iV5g=+Hѯ�?/EcH����,�S'�B�MOl)�����j��'af�XEW3R+PK:%,ߧ3�%�E1܋3��g|�\Y�Z��$��q�3��e&Kܫ���5�&�f)�M~.��@�4�6j�~��6iyS_?>����,��[���u9r@T#C�҇��N�qA�^A�E�������^w�彍��"�e�"5�o7����Q�hkn	��2��@�s�ū�1zF�o�4.ҡ����R��]>�?+x�6�m*t�$��M8eO��lK秎�״����z0�ضŶKƆ� ^���n''&�MT�G㻫!΃ة���)��E�+�&��+]��H�%wLjmhr���n
���z<2�!B7��'�'Z�S�/���#� ��2 ��M�N
� �vBk�	���N����[����0�ck�FV������V�����1��\I,�6B����V�����쵇Kc�_�\�Z����1v�nZDU�r�m"��6��5�����h�^������%�Ȝ��~w2AрV�ih�֏��ۮ���K�0Rw���lo�{NX|M�H��X�t�߁�R+�C2����:��#���CI���ך�������N2*�G+�3Ɓ�Ƚ+&ղ�ys��h�B�YW�.D��4�������f'/�E,��ʱ��l�c���3�G}P1@�]�<����~4��ۄʰ^�p{b���Y�{���#j�d��p��"�U(E���	�ж���D�ט���)*4���Mq��Fn��%O�рB�<ꃏ�S�����9�yU����^��I�1o���-��9W,��L���Y��6��ܽ�@�n�+
�d�����4eY�u�K��z�Kz��b�$���lo(wP�
Q�ǵ�葦��b3y��zFؤ�X@�K�*�e��s>�~�So�u�
���8����{t~�[���P����L�5;�v:�,�6��ߢ�h~L��QF�j�)�-hhe
EViV\v�E��c����%/"qe�I+�V=���}!.ɑ��|�遬B��������:v�J�ww�i7�dI����V�H���n�t�^;�D�.a���!�@@8���^�-*!�Ni��c���Xk��˫�6Y%�Y��Yi��S%g��i#�Z��>ZsQ��1xۆ��9uF�=�0Z��?A��7AD̀�I�Jc@~%>g �:l=+��[f;|��u�/� m���Po&G�I1��j���gψn���Y��Ȼ�*V�2�~�7@Ӗ��=�k!@J𮼺��_�G��Ŏ��5B��~�x~d�@�8�\*�V%�| ��=6)���̝9դ�N����|GD�Ɗw'C��C��ReEA.���/�t"֙��l���%�Xa;2qmG��5���e��d��4O��4yM`s��"G�������n+B�Y>�Y���/0OpjNK[���$�jJ�ل8�%�� �:n'�D��K��r :�s���y3���4V����NAO>m�̋��i�1^3���l�h�e�q�Y�������>�QD�Xp�Lcx�
#�f�X�BZ ��2i�3��u�쓪�#��J:��{�?vhP>U`h�x��0�⬹�9&�ê�~UB\�;��i���\ܘ�'��R��,ښ�*�ߚw��s�t�J*G_W�́�G�}a��9�_���v:���JxF2�A�G6�q������A�3�s�J�2+�[b�)׳c)�ׁ�p���Z�Ǿ��S��\[*5�K��$G���x����\Y$�f�$9صc�����������Y<��:�|�K>.&�3��꩗��4��|q>�*mdi;!?�T��D�A��{���L(E���:��]�B�ִ"Yk��-9c3����)C"�G(d*Jr�k�}��a��Y�.Zw���DG���7�⏝3*R�]�Y�|��[���O�Ց����oN�r����vJ���FeR�34��4^����YZ�T�������e7{�N�!��r�`b�e`�逸��`<9�g�^ UG0<I(L��	B��Ğ��yL�<J.�A�;\���#s'���N�|Ŝ\���F��}�_� xP/�N��b�2E�IE��47e��ڠo�.D|r��_�n"�7;o����5���Q�"�^KD�&�������2�H6�t,/�?��]S��:�(�<��2mu��d"��a���a��n�I�����SiC>-��K�&����47���Z�1��tY�
@�P;�RO�2��W2:̋���G��LR�i.�$r�V,x�&�'%��B�p�Ծ��>��g�Z_~���	a0��NJ����anܑ}�{��^r�I�K�UO�q�KP�d���H}-����?������1��T{�=��	���pbg�'�U62b\���闱U�,V[-�,�y�����Cu�_��g+�7,�̤|��Jcc�91���N1ֻ��f�`4���P���kq+�et$��4��h�N��%�Ջ�4������*I5R�D�4��Ҕ\���]5ٴ��ݽ����9Z�����qk�)��|��h���a�
�;m^7�>US�%�a�œ�\��[�i�)<j���C�DeO�"��ZMqD@9�zT��DS���BOH'�-�x�:�J
d�3>�2��~d.������SZ���k2�4H�r�.<���������x|\EX��7B �
,�3�v�`��Q��Њ	����*���HP�*��?5���#����2��yX=�#��otV���<���=�u�	���3t�pY�[p�����`�i�&���X�L�G��y�9��Q����Q�`�.t �K�R�Z=Qw)��Z㴿&��0��
pk'^��n8��5�0H����LYE�����-�鑕'�1����:בŒl�W%�����O ��ԃ�n)N�x"\����� �d�2J�K��h�T�L�@�@��r*/g��9[�PT[�D����3��ҙlc�\��`�4n`rkDC�7�#���[3Y��Y����!l͸7ْ��Sb��=�����Xm�Bµ�V�=�)0_9W'�q5'�S�(X4���囈h)�ژNI}$�Ǩ'=p���KGF"���B�#�۪��$	O\�cG#JϏ�t��t�=KgN�I-��S������58����*�u^�5F�b�8�o�/u L�RF�`��%�hT�N�S���謹ژ(�iTE�Bx������!e����N�{/l�QH̽1���J��K�����j��t��(�SJ�����ݿ���c�X�8���RSS]� ��L��D�ϯ�k&�s���L^��V=ٻ|#��f߹��cc�Z9�oRuy��V�Ogo	��Q�����u�攁s��7�È���/�y��PG�d�-����L�5�I��x����Q!������fHeB�~���#�uW9l�H��g\r�#W��^�R�+e@��N��ؚ��/3��0]�����o���`�s��zW�>`3�/e'=;'m-$��cHTEK�ӵDr������ހ����Es��I��H�ס�/��.~�޴�^�����W�W'>�^�^�;����t��D>!���4��;c���YnmG`�q�J/�
 K�!e,����QU����^@�O���Ӡ�s�!U>�����|K�w1��f���A)V{	f-qrᏬ[viB`��$$go�9�m.�]z<��,0��ι�N��`��!=�2��/VG��-��8��Y����{c�������F&�6-�Iʘ��r��-��	��Bo9�kY�{"��/��O����$����S��c��������v�S�E-hc*%�N� ���cp�gi���z5�Xz���_�
s���t�h�nl��1���Q1�m�`"d�D-F� �=���,.��Y/��������[En[8�V�~����L{�*�v�,�N�Q��
F����O{�1��m�UkT���z�X;�nd��6 �b}�������p&8Ճ^&c����`���y�{r�߭G_%[n&�H��؈H��X�4�)_�oH��L���]ƪ�M�[��������
����|�u�8[xv��.���uZ�+�$W��;����9��p��̆B�\�0���M5ӡ��hBu���p1���d:� }��k
�l�qH�:we0�?M��+�AQ>T�e �Oe��^ԛ:2N�N�O��A�e���b�=h��=��P\gF��@��2]��m�98_���D��Ua���~5k�,��s��v���2��1g���]���I�(�}]�w.if��\x�'[��[�7�	����
��R�krB���^;�D֟�gh�ӿOw{7^�sI!�f`4��+>a
���jL��L�A��KGL�+�̛�m�a�J%:����C�1�@��6�l�RVk�NDd����>�]�)gX�s�󍖙ϔR��'�'�cC�O ��1l\��U�DF%!�9w�<c���ԭd�ä��Y�7g�ĔM&mg���{s7�}"������X��PEf3���V�)q�o�����;��sWX����0�`NG����o<������p��]���L;%����I�^TZ��hw��9l��A�{�h�)�dR��,�g]�m]fDv��/���A���~|G}PIw\�2�y�5��)Em{a�@,�nE�d��sP����z
� �ڿlJ��n):���D�5^�(t.=��D�8�(_�����Jz)���C�Xg��]Eϙ�W1�6�<B�f'{&��,}��k'�d�:pU^�ED�b��E:���;��xp ���jL�d1�0�kT������g�m��f���/���0ȑ� / a�B��l���!�?FW�2H矋��)�ͤ��ܷ��8��%M�+����^	��|z{`#q9ߚ9v��{��f�7D�=^�[� ѻ�l3�F���8�>�ԫ/�	
\|I
$r�b���c�?�Ij�0'�Ѝ*�6��Y��oS5�k���"�%���+�8�*����N �c��Bg�C�*7�S��	��~��s�j���ab۱+f��i���@%1+��HmJT�0�DW��Gt���4�9������>���Ey�Wr�ކ�R�&�SJO6ɣ-��*�D�ʀ(�'p�새�K�I:��*�_����H Ҙq)X�2���c��P�#�o�X�����R����x�L:�Ir��n��W2Q͟0��'d��,���dr�g��iG��&��+I&k���2�vX-��p��8Qo�flwfT�\JJl���q����)��*��D}���� vsߥvC;�
c�C��k3��w[sctt!�(����@,�ۧ���q��E⻇j��]ʂ3_��^��]�=w&P֤6����������:r�e5�!@�V~>��Q(�y�p�76�����s��:��bc"p��o��g0z �Ӟ�o�G�q?9�	����D�>؂D�΀bUi4���6�jZ�Z��/[�Df�a1�AQ����q �8���[>
�u����T#]�vgK�y�(���:2-* �/�����V�d���^�N�YF7r��+� C�{��,��@Bf����%�#o�ns��yS��g��/�/��G�ב����&���mN�:KW;zM��Տ;̈9����Pͻ?3���cM�1Wb�Ə�,1���������	�+�S	Qo�Aw�����I���R����s�K���N��e��7T<��`)�x�>��� �泎� g�v�@y[2%������-LݏS<[��rq�����ejBKO���^8b����UlJ+]�>�k����=:���墯e��,�����D�fQ��\.��	^���<�8:E W�#�&r�:T��"�x��BK���nr|2@cXz�A��yO7}_�q�S���e����U�ZXy滆z;O%�R�S��RO��w��:JŸ�5�%W08�&�S�A(Vէ��T��ׁu*��k�k�P�v&���ï�U��m�e&�A��]��J�~�b�Մ�*78r��`�f4�WƵ�6R��Z�����5�#�*=�P?���J�
k�>�����k�KF�rc��q>ד�`��l��W������u�p`҇�b���$)��oN���	�q����Ǉ̌��cp�_U�}`Ї=@r:�3*j׋9�Y��⒨w��?c�
�(���s���
�"�,�C���J�:��;�����4�2li#\��͇��w�)_B<h�X�S�R�y��ղS@?`�3��o'}�m��衻ւ����!�6��q�ڼ޷{�0�A����%�K���JOLu�_ۨ0�B_{���e[4~Lf���Y���aG�E�X�@��S `ل�+��m���hZ�&ۙ���@�Qzas���I;�Mj�"����b�DK��E�g'v_Qw�՛�C'ou�`�^�X=�F�;�����C����j$`�� �R��H�5G4��h��V�}�\_��:Ɉ��ϐ�[�4� *�*7J�,Hj�R��{&��s��?�e�$�}ޚf���c�Y�����`�f���� x�[�:�"ђ9����[)J�H��-��ZI��<�!��̒TV��
:8�!S׭�$�Cz��l>s��1���N�ã��h��X��T��,����I�)�n=�jX�X~�1H��n���N�HWJ4�oҤ�_���E�U���ł9� �A�V��Vr�V��gk�=�� ���p�F�"Q��B5˄��
���$�2Afzcw�|��!#;���w���D����u-�B�������c�X�m���S�U���b��8_�I�mVz Wk,6����۩���l���ͬ�,˖�=�7�BK���z��`��U2ݵ୷�'J�&�)#�oV�d���f%&�W�3K�R�<VH����|%5P Ц�|-���ѷN���	����šN�ƈ𽸹�3)�+�őxVx��Jh��P)�i���\j_�6ͻ��;�m<:�����I��K�e���8ډA#���'��	} ��>��[K$����-r���3���W��&�E�q<���a��o{��\;��ɾ��P_��r �%��W��,��#�a��2�P�y�q��0�#�|�Iɍ�Z���^��0
�QΛy�.Q�ÿY�C1���p�v~G�����^��e��$��;����jK}��$ji�+�T��t?��&�۰���7ży_ˢ��0�
"m��e��d���z��N&1|k訝��B����:��y'ٍL�6���Ї_"1!OL��Iuy���k)
���[�N��䷖����'zDR����I�E������ɪp��wmo,MZd�I'ƥ@�ŏ`<u�]��P��a����L8!D��h��)b?�Y��Gin���mz��h���څ�AΖ��L�gQ]��N�o����qv8��NΤZ!h�n��O��˨�w�d��?�����em-�厁4�{u�F����Eݚ�I�o. ���b�v�`�&e\����"Ƒ�=g{�~<�/X$��ܩ�� �V�����o�t5�_^Y�#?
` ��*���(M�qt���Ԧ��r�}bQ��}?T$����Q3�&�Q���U䌰����S�@�F%)[�����h%�8����?�ނ�U��8�
�hF%v�6�GŬX��^�kPVؼ��0s7��`CO��c}S	��т^;�j�9Dt�npS�~��)S�2ͮ��_�(u�aĹ�6n��ȁ|��:���O_8�.��W�Y�)��1fv���]xٲs��q�0�?>n���fS�7�q���J!O
����_��[��4���*��3���)z����O����Z�1O�������~D˯�0yw�cb�3���Ϩ�����hZ�(�S�����s_�@�z�l;b��&�C@�M��g5>GlPG�٘�B�{�M�!f�'�q�1�)!�<��b�K�b
&4��-��^�*�ͯ�Q�4��<�9aK�s�c��?�^V��]�(�2�hu,��۹ʏ�#<��9�W#0e'%Z��P����M�� �|s�m)%i�l�����m����>;�G�{<}j`Z����kjO�Q֧SI�R�C3� 4,�FY^K�n��`�x���ՌCa�!�(i¼�������X5��l�p��f�Z;�0��%���9��+�>�����
YXhx�R￵�>�W:8:��T�ҧ��d<Ջ�_0�nV���L��C��#������
IR�6-�\��m*�;�̱2���ý�/��֊��Pb�{��98t˕"��2!��;(��9H�kQS���:�%�R�,Q;�"鑤܆�H4p�a��%�1+K�ߩ�b����$b�*҆y|D��كOv���Q��J��zB�1[?�@~5�Р+��C�9Β��	krĮ�:��ɐ(�G
��n�B��w͟(S!��6Opȿ��d��L��U����)�*�zq�+)�iqE��`f�r�����7�R������X�3�΀.��ct/�R��ȥ��k��b4NI��~��JNu[�q ����7!���քOc���l7�6��`�A�e��$���)����V���$��8����a��62-����5"9�~4N�$��\2:��(��rX$�$̼M0�n7�f�I�χ?_N�8cQj�?�yc%��d�yھm���b��O5�G�����b��\��-K-~뿇>6): .$W�� �<�g�~���%mń�
��E	0�>����I���N���&ch�ֺ�-t^��b��y� |+��20]��{�9
���ŵq���3/8��p�[ ��D�G���hc��[�����ٷ�/�&?Hk���OD����^2CaW���x86�`ʵ�{��C�f��"�
|��
�(d�m�j߅>��48�1���椴�$@[��R��&E���ePk+�y��0'��S�������a}t�䝸�w�ǽ����c?�l������Nm=^~Ng�ĺV���
���t�⦩�t
�#�Pk．u���� ��.�d:W7�c7x��DzC�Cw���c��w�C��� ������*CI_.�06�ꈒ�\}�o��C�!�"���7͓cz�Lck������-
�R�u aǋ���+l�u--"m�Y�(�\-��My&mr��uPT<ď6Sd��R�Z�C5C�g�E4�b�@�P�K,؀Nf<䊮�N����d�Mv#���R��բ��?|����7���$'��f�0nv��1�Q�F���>Kl5��e���U�^�y��"FaL����^s�E��^�!	����7��;j�\f�%�����X���{��H��
1��!-V��{x2[��͘m�ꃾ%�Z�*��8����d�H�tl���>�V)H<�B;��S�l��KY��ҳĦP<�
8X7s�|���7%ig�5�é��b�з��է�}Hqh�b�]�3vE�,�����C:�b�y��������+>�S�q��&#��Fb���C�'���*�z*�?��1�moJ������_,��E��ʨ�;��eS�mX�a��ٽ����=��ec�U|$��Y+�����[�;�(��&AD��+�u���"���L3�D���!�]3�wq�F+�a�� vWF��׶a�H��h�Ҿ��WǸkq�$o�y��"���]�� �v���4ؓ�Ϛ���?���x�朕��6:�h�����Sm�J|���T����M�]���	\=����J~V�#�X6S�7"C�l�`�~������ĹH�Sgvn��f?����?�VK��T��^�;��Ϧ�C7�)�;��\z	��z���0��q0Q�
{I��('�Nn��2o��l�Rh��\���^�t|tn����H;>z�$Ӵ�d�� �'��o�iJ�}��h�B�(��#�T��~N:�-jzs�'��pQ� ��7$$	݂�1��sF��1�j��nLؑi7v+���>%*�y���>���xܑ��D]'���MIn؉90�O����*���lRt4���AQ��@�zy&�Лܗm�����,_u\(�{�]KyELL���4����p�����D��Op���b�b\)�8,����)/����x�@��J%��ENf˄���B~�p�@b����w�rڠ����{<��J��l� u�DEY�?E�)�M�E����x2�߳Z�V�k���ayw6������� dP֓�EP�]�<����'o�Da�(�������7:ϐ������D�����q�]��!QT���$����b򽡇!���5�B`��-�"�:_�1U���e��U>�+�j���(;L`[��/���S:��,Fۓ��U���ȋ!� 2��؊fOI�ϙ���'��Θ) �5���|��w�~d�d�q��5 ��є�g>$�*uI7Z�9vH5���5Â;<}��.�%��V��N�p`
i�+��x}�����P��p�������x�����Xa��E�@��.���A�%b��166��S1N�Ѵa36�+8���u�@��c����':�#���Jwa�2W	W�x�����Igѽ��:�x�s7�bBz��Z�s��uf=p��"���>�ۻ��7�\��LO�K���<&5�����|���@�V"�`����^%d��$Fѓ���������>I�����6��z��_ɮ�"��h���MR���;�Ȧ/Y'L}�Q�˓�#+�#+_-�ey�.<<�	K��q��:�|������+ �S(�5	"y�[�(!Eq~��}Ɇ���u�9�ʮgܕ�yZ�	����5��6�톕P���#x������3���qB�)�Z;j 3}i��sO=�״����L*	���L�����L�z]v�ʟx������WjI[%'XG������Ί����ʸ4G���r�QO���F �-��_Ԉ_d��߆N�'m:	i���6<Qu�I�/#�i�{"J�w�W�?�A�8U�%2I�
�t����ָ���y��Z�ڤ�H�FŸ�s1�<Q���\��곞����H=�Pf`���zu?�@�`!g��'K�R�w������}6��
��e�\��1�Yz�D����ͅ�Y��yb���������x6%�;_�����z(�C��j��?�߯�U�P1A�n3��#�Zp���ـ*�%9Wh�����h꼲W�)%\���l�Y�}c&�㽜匩Xj��w8�r�W,�T�gQ�
E�Cx�]B�Ȭb�� l<S0��8DU�WG~��ܾW��X�b@.��D!�����S���`,���Q�b�\�� (מ��*�����&��)��������WMH�DQ������d��"&Ȉv���\����_@+hAJ.�qK��3�"|��Lw��9��I8��_��6c�-5ǝ�n>����zT��^�|�^�Eą��x�T�f1�h�n�U�#{��q)5��&�7��4�9wv�}��թg��ό����7ނ8��等��P�y|��}]��Ҫ��<Xw%�Z�ldZ�3%�\��%o�|�Aq|�<�qI�m���z�A{��2]�J�^�n�EYI��C�L����Ր�bƙk�" A�s������'ޣ�ˇ��؄�5�]�޼��v��m-<�)�H\ :cA�:Z�'�ژ`�yN��t����Z�4�C�Jst<�ك0�k��ߣ�[����;�)��Q�m�E�ɀ�����!�RH��FpL���͖~O��J%�~*����I��>5�#+�cw��Ə����B���&)'�i�Ep� fW�{���@�/e!���?N �C
"�	�X�1��>���S�K��)")̲r��"��q���*ܭ�����&��?�c��?�W��U6Hh�j!Xx���\����d��� Uꂢ
��;�!�����w�+�Ip�T��e+�##�\B{�̆m�qe��P�g9��]�V��t~���	�q�B����}t:�-J�!*�r�#\<�������"�y�h���S�E^WԂR�ŉ	@և�߁բQ]����Z���R�%�<�p�p$ߎ��K����=��fT�HJ�g��Y�~�*H0|:0!-�Ղv��z�־R�J�.`���-yV�
��������~�R���)G���k!�X����8���V[���$R�9xt�WJ�_+�	�d'k$6�WA�U0]:k�s��.3����b;X5��]����AP	h��Sca1q�$�>&H�U����S�7�bЯs��,W�WQ7}�����Qw��qgy��&�cJo�NE��m��^42�����}���
�:.�F��_h
�.�Tt�0oL�ҨbĜ^�g�x]3&���B��	�!��\'g�.�@���NhQO]���h%G%@�e�wbx){���+iW�_к�ԧ`��c*�F"�>}�y�`���RzY!T<a�U�[�8�����YM/��(#逷�O����Q�N��CX��u/�xP��8Y,%�����te܈OZţ�sa�����Z�J ']�+���$�~y�|�2�'��9=��Λ�" Ċ}Cqd���xA�[�!j��!W�+Z5~��)g,,#��q�'Z� �8QC7D�(�y(5B*q�'}��z��к[j+�'6�6�8�H8�0�T�_�N'� �k��H'���Jʜ*��S�f�Ngt�Tus�n������z�MZ�8��N����`)z�Y	W9&Mk��4�u�H��F�#gdՒ	/�\��%��l��^mm�V9حz+���!��t����؝W���(�j9`��MYO�t;[��'9ޫ���a���$��4��~����7�����S$86����V�`z�ik�a��)18˺�h��B!����:|�r��ciS�m�p�ˎPK��)ÿ����j�.�����ũ��l�MZ�o�c
`.x-)l�S|����
�ݍ���c�	��jm�Ϲ��W7���T����,@b���">��D�jd ���1�s[� ,̪�
��M��Ѱ�[�V%X[�"j��H�����} R�0��_��y�}��B��?�a>懸�?���|��;�NB6yz(��M��<?�����Y�	ĺ�ɭCs��!��9'��}@����՜H�A(�J��lF�_��{n#�|g��ϩ��R	'Ex���9J?��a�Y9���ϗ��B���B[�0�ѡ���YmF@��σ����)�rjD��"O�E��ƺ�X;�:>�lY��t�uD�XT�&㿂�7�x��p>��`�0�����Ju"����6�GlO�D�҈�|p^/�E�R���o�GܶjY�}�=k�興��oU�<�b_�DF�L��U���h2t�E�:���tr�]ʭܚ���<�����Ғ�$�m.V��/���Ж ��W�'К��aT7DG�'&��� /�`�-�6���^����n�{IԔ�?^��E�H�B!�=���ߋ�Y5 �p �z�Xڍ��Kwa��3�|���%�io�F����b�"��4!��&�Vo�=j�L��n���ƞ���՚���	6�/tٍa����Z�
Iv��F:�v��[����z�~��9�RԗR���޸��ct_eTu�c���'�`������]ub���b�'�����'M0f�����{���:�.�Y�m�����g0��pQ�Gދ�𩽽����1gZ���mQB$��-1b��v>���D�����#~��Y�Ѻj9�>S#�F�u����@<-���0@y��R���� '=l�0�H�[��D�Ģ��#De�	D�Kk��MdW�C����{C�RmI�n��&�ӑi^B�	��o���8U�T<���Z�:�?&Q%�y|��V�=���o'�O�x@��8�z4^��~�,+�� ����hN|�L��o*�H��M28#S����//���bV�A���c���i�b�D	�6t����U�"�����0R�VY�����h�\7�}Z�C�Y�n���$���R��7��C�!'�b����VgvQ�Pd�� W}���q�é���[�|A�L7�q�(�V�6�m�����V���;�[�ԦJ�
�h�ӵYfr�Ύ���,���H�����1��o�{$��eU_dn��g�'ζ�zA���-�A#iA%	�E�υwD�S��2�l���;cپ�3���u���>_����^�]%u֒waH;B��B��ra]� `|ia�l,9�:.�%�-n&��`��B�"�d�b@w�Δ
�4 �E��ǩU�l4SFbG;����U��7��R��SZ5M�k� '�?c�W!1�U��� RS"z�j���IwMv�����&"��j�����y��)Jn���T�����!�k������-�ulO��|ݥd��V� O&*?�D���˹\ߋ�lp����bQjB�邒k��P�J�����,;g��8���0k~�zq�6z��rr���s;�桊H��� �7�R��X޿��������>Y@d��Pk��2��R�(��7�T�[Cf�vs�^��!%��x�w�����y3ƽ�e�!o��ݱ^)GT�ķ���q�~����9�^�粼at����idGd��n���Ӿ:�y�sX��ʿ�_쑃��=��ʚ-��R�ŠJtIE�A���0��1���{��*�|g��m�9A��&�Y��a�������};�V���]�A(y����К#��V����G�����)L7�^�&.V�wO�!Q]&k놥4�&ֱ���I�L���2�x�����#��������H��>�K��1'OT);�tz�O�9��5R��n:ne�Z�	6������\7*J��P,6�i�����:�[��]1�g���s�ن�l|��bø�����C,�2{�,����;��UN�#�#D������N�/����6�B�.��P�`s���I���� t��{CQmP�{��[�P��6!�y�?�wd?��v���D��R�db���z;i�%���;���!��^d�T�	^"w�^�VS=K>���D�~)��tɏ�ts^��)A���%�
�fR�dz	o;/'��$������T@��!�ط�)~��i�㥳�"fz����<��2p��1{����ۮ����5�bU�`T�8(e�-�b2��*��x��P^BF}�j(�i��x9�"�DO�[ŋWG��A���]k��r����I�|���av�i��)ؽ�-|�T��\K��xyЏ����SJC��>�� h7�%P�U�|Nu�/x�Jӳ6f�(1v�`Rڦ�o�8�ۖ�D�6��6��$���!ɕ�U;�adg�"'$R?<��5�g�2���b�?�ښ�ǌ�|f�	�Ɂf7̋�|-��$uZ����gl)F:�f3�9�u��j�� N���x�8h�ͺsFoz38�W�p�a�+�M+j�t�XRD�PN}H�l��o����V��;h���@�!���r0���+yFp<c���"�@M[v�",�_�\>��1�C�+�^�"�� ��k8����z ]���
DkWE���f	�������I��/�g�-�$��
ӣ�(��xK\�OrfǑ�d�i�o�4�=�p�5�cʷ���Y]�?mqiS��ٙ�T0�e��t?�{7�\��\�]��t!����4D&;;��=�Sx�e���s?�b�Ç���`v����?B���/a�Ŧ��Q� 83}�zR�P�*����Ģ�g������O��+������^��q�����?)����M/[UK#n1hG<c��YS��Q_rAJ�ƕ�v����kN�٤>��;� �;���m,Nh0f�X�P����T�c7+a}�s��&����|LZ�/�t%���#�KÍ���j�o2��1	�Ή{�)��fgR�$�I-���3��1���p�0I�[��.t]J�+?"-aH�(��[�u_W�i�=-Q���\��^�l`����"ʎ���N(Cg��<�W�!"o�)�ۓFd��S�+*��=�|��+!�'�P��-č�~���$"&��5�̏>w�;�%�`A>_�%y/�qoP�,,����:՜Uߞ���#�l����`/�'r��w�/{q9L��7�f�w4���ܒƇ�:�!:V�tu��%��`PE`EEUnN�\��[���! �ܖ�Grr�˚���\ܯ:����� a�w�0/��-$�f�!�BG\�n�+����Fb;��Y9(��ENR,��r����L^���Ƿ��O6�Y�[�uλ%�r󛷍o y�T�AT�*�y��������y�tDZ�<Z �<c��������92"P'���7�������:�*��W�����\� ��K�O�
����,$���M���D�Y�~���_������HFSGO�Qu!��7�P(�Ϝ�P�	��s�A�Y˜rZJ\x��
�=�ͷ�C��V3�;G�q��5| ��=� A��!☙�#Q������ԙ��*�F�>�ed���C[0�}5��i�޷(��F��ʚ�0��۪@]�˥�?c�~c�3��c;wz�ӗ��f�
N#8��),� ��f�K�՟�G��� fY�V'���E�q蟁g`���؁\㬍�yMMd�w�(�8�:8�
����֝������5�t@Rh�TXr4��;k"�'�bNY��RPV�VpJ���o��&`v#-"v�\��A�W������U*��~ +L8ם���>�\�ns"^�W���xN8��G{��W���a���? ���J�ƀ�QDM���
$���P1WNt�LC�a���rl�vyD_��W��H)��*��,h���<i�ms�G�f���\�2�&�K1#2zE/���޲����0�-1����˯I�<1���eŒ�u@���AvNA�xl ����5�U̟��dqy-�^���A��欮:=x�k��S+J�&ϵ-|2�89k�������6���pttz����5������ғ�����o�j[B�^?^e��	�T�Wnf��d;�g�'��8u�3�������]��ʅ^B�
~ �P�>�K�@~L�ۙ��!�Rn4�Hw~p
wΤ�繎w�IkO�R�����L'y,�n�k��~�*��HH���i?
�V�B� t�!I�s`r�a���}
.'�Y��9���q��RB��z�yd�xg��/�� �$ܭ����`��Mۋ�J��b��_�53����(�����t���|Q�W���)�1�?��Ѣ���ʡN�7.�]R��8оRG3���Qcv�+Ogu����i��<�aʱ��}�lnm�Y`���R��c:WʀN����ٜh��kdC�])�ya�H��(p_܂��F�l���X����u�v��4��Ɉ<�aD!EW����S�<-��؍�z�$4��nRm�۳�4�|���������{)5m�e���Z��@��w��\�-g۠';�W-���-R`[+v��>C슖O�����7�=����C��Є��Eu��ۅV�*�V<�U�U�TgҐI�h��1�а����GdF��m�C��r�?F��w�>c��{Q��}�9��V�!w���\���",��M�"$)!V49��ɳ���I-��A�����o��<E����yV=/K��:iR��֟X�&sW��@��ڬ��_�����v�kp����M~g<��}L�>����/h��4]��M��l��ts�qgU��ނ�����K<�>��n��:B����j���.n�-?q��H[A ��q1*�m#�W~�1�x�&�M;�k��&*K�n�E��n����g�~ ��jҵf��
j����7�+,d[;���j����Î��s��%�Ku���.i��5��z���i�6Gx!`�������'b�/����A��Wqƫ�>�7�@Ȓ	������U;�X�މ��5(+pk�N�'� RёՂcaT$�0�JFy���a?��*�֥���t>}s���wE�tx��P	(E�9�lo��o'Ѳ��r֟� ���T���)�t��(��{Nf�E+A'���|�ʟ�}kۦ2.�z��g�,���<:���޻�{qi�XT�W7�su~��B��I�w�{;���Q���B�d��s}�u���}���V,�s�_�2z� �#��F�_�6c�&M?�Ú��D��"�w�a�����g�'Y?4����zΩ�a��u��ܼ��%`㠹��S�vٻN��YL	��ET۷�ƤQ��.�� ���B�=(�Y����wg�7�qL�a�A���8;����C�CL}c�	�y�=)����yt+����UOu����dkñ��׫���W��D�c&�X� �o���Ǐ[��� �Yn����7� ~�f�d�&cD�P!z=��T������D��L�AO�1�Dp�4rX{��*�w��fB�p�|��}z �eP�N���<!nƽ��%�I}1z�9���]�Z�0�=_=�|X��~����T1Hӽ�k�������k��Z^���1�����a��+��]�T�%�6�&���A�i`U
h_@.JE�$P��#���{���]&��кDyvj	�g�Ү���C*I�E8׮�����mW�U(<��腵V؊~>s��Zd�[�$wr�'�eC�bWGU���3yO9oDr$G(AD��Z?q����������r1l��Z�+�I1o7�R�h5-X��s���mi��f��K"26�@Y��zu���	�h'
�C�'���>|�3J�Ȩ�'�]e}���̯��E.�W8�1�e{��$Q���yBT�m(3g.)_�3�w�T__����?
�2��S��~�2��3�q�9�汗qJp��3E�_�R���3�T=���n�K�[��֣E��4m`��f)
�U�@4
1�1}ړ�#�[�4��y��/j��B��z)��	�ۻ�k�+e�팜� ���:��ʈ�
Ħ�ʍZ����5/nW�cZ�Z������
�uѮ_��"**��bPN�6*�Po�F���*�0_���Ż�E!�8q��3�/�ű��n,��2��3M`����;B������;ֻƫ~7v]=:��qΆHS�A��*���vHֱ�Ig|8I��^�E�c޴�18.�0��M��y��Y
'U�Jf"F��dCPڹ����
L��iP�Qt]i�0����F����҈ �/Uؼ�CR3���a���S���_�K�ϛY�.Z|����]��ŋ��m !���� ��G0d��p;�}tm`��9S�:�b�A�M�w֐B�mՔ!(`v�.�j�O���-��xO��糦Ɣ3,��p#���Y|�	�8�pNs�$���_��~TR"g�1Q��݅H[�a�\�<n���
F��X�{$�݉��U���ָ3�#�xp�C��el�m��e�f�����agIz�%E�f./&Q�p�����kگ D0��hb@\7�?2lw��*T9����.+U��|�@�3�9!�"��/�s�*�[�_~�C��'�%uƎ�A�ܯ�<I��[����D�i "��E�Hr3�6(C\lϿ@����f3��0M���ۑĽ�!O��6��n��m;	#A����( �{C	��<��鑡MT��Z{�m�|5 ~�?��t�(4e�i/s�q2�I��#x�<�\���0������G\j~@�%��vΆ�Y��=���V�ƚ�C�Z��OGe�	����:�DO�r0>��� �76��|�H|\�����%Us��7�s�i�|N;YD�D�&Sr�Cy�/a\�7h>nّ�Fk,��M֬���� é֥>����	㊻�f\��M��W+��.�>L��:���:>�0��.ŏ��jj�;��������Y����4qQ�4(�c	ב?4�Kʹ��FG���Y�Z�������p�e4ۂ���gԮ��Ѳ�sD�Wp��L�~>B�ԭ��5�EZ���ZԵ�|g}p���I0��P���PTIOZ�r�Cp�p�r�:���"�Q����,�n}8k7W�O��l_k;F�\|b*f*V�Ǚ�!�*�,���ؑe��*��w~z��,Y��+V���&y���t��(_�18AtX9�ϊίH���-�����Jlʣ�Y�d�3�V�����L� n>{�%+�L�BT�g� m K��f�oeD�r	;sM;|$"�'�8�GPhWN�$I���(��xd�td}�C>Z �=8�ܲX72�m������$�z3;��lY�)"1�tx8��ڀ���i��U�@^�<�!��9�nO6: uy��l��6{�-�t|���`o,��XG#
~U_�WhMw�3���_�Ф�$.p��o��Gl	8�����!�Q�T���o�B����L�+y�"d��;c�'Kw�$@p��94N\���!����J彩7�e4؏�zP���WۇE�'�ԌE^��\W7����N�N���EXn�N�7���c���p��`�P���o�\��Y	�T�D�zD���ЙАuV�#<�$�qB���5I=�}�8�k������:�A%�|�n��1�:A�k���'����ݩZ�f��- ���a`��Ԣ���c(�_�m�t�<�^�� ��]�Q�Xy������r�@�Ȣ�}s6Y"���w��� �Rԫ�Ӊ�S��l�7���غY�k�։i>�u-���uPuk��AN�]�u)i�Uݯ|�@��{%�]�7I�����Z�Mw����]V��Dg�J��yۡw�
?�j�o�"�����Џ�4��&��3˯���Ur�YRG��k���m��8�A�����^�4o�a}�g'E�T���������E�j��}ϟc�~�UY�!Q��k�n��L�d*���ݽ��J�l=���oyG��E^�σ��>!���4tˇuH&�����p�P/��&R$�൸A�E�!�~�=�����]���3���!���t�ٹ-��L�e�Ea��
 ��[��Qx����{rڲu�:F�,�N���?Dh�+�}�pw]K;�O���'df�k�Ы��.�I~2�Bp�����xh*�wުo"��fb�vsM:vɺۅč��8�s�)h�q�!���V�%��bB�\s�!]����XY�@[�ᇫ��q��&��ۧ^�.���@*��}��A�F�<��3྘d=M���o{}�j��n6������)���m���çu_Ǜg��!��A�ʰ��q�)n�n�}(��UO���DH�ſ�/���i~5�<!�ի�^����I�e3�#p��t%��T��b�Ѣ�<Um+����M�@>��n	Tr�r���4��f��Ѓ�����(F-�K��{����8��H@Gm&���Q�9�j�$c�t��i>	�����$�( �#*���ch��s�#N�(~� �Ⱥ����3�q��	�wy<~�i	t�Bb-�ÖV-uo�q4�kz�@Z�dN�~6	Y����޽|"�ؠ�*)f0ꑃ2[�nSA����%����'=���~mA��&(Umi$"Y��-��T3/���NH=�cxZ��J6:���>��l���-�~K��ݎ�B6.2�	��~���g���]Q�W����e�wG�)��	w��E��,��XX�_��(8d��>��sg��l#��UL�)� 8Ą�\�#�uC����Ku�F>CW��;������Ea�'�*�P:�*���p"Au����Bޡ��@�F�X�]�)�zrқ-�ŤY��t}/J���@0�\ʍąch���{�# ������s�%� X�{�b����F�v�}�TR?���:\�:D�������.a��]]|t�ϥ���ժN�Q�e���hd%z�Q8��S�f
����}ؽXq�<�p����A��/�+dǗ���������41L�h�8oO��s�pY�͈�̠LT���'����څ'�|�W��᷽�j��w���i˾�^Rz���i��J?��V����Z˟����KV�ܻ�g|G��
���5mr]���
�L3n���Q ���=���{�ɀ�'��c,�Aid2�H	��!��|�B��Q�s����VF���6U@�Z�����Cc�A���!k��,��،��ޖ�j��|�Pm7��5�-w�%���r���R�?��xv���L]xCo��9؏����A��N�"��z������#qD��ݱ���Ɯ��w
F�a������I��'�nA�+�>\����*����0*���O���l�&�7f�a3�a��k�A)He��Qc=��D����dN���Wo��xs�)�Ir���x�I�w!^ �<]*pq��8B<mQ��Cyei�81 �v+�1N��{%�C���Sj/�sm|�ᕚf�y�6��=?6�!��Zj�郍�@
�H&��Vz�0�	��GM�C��=�f��ˉ���%යF�!��Ϯ����J�}��"���*����0���~TCW�v�'�y�7�G5'�窡�������Dv��,3 ���+��D��sm��H� ��˛Ds�p��b=Akztm�d�-��!�:Qh�Y�;	�W����FZ�p��,�t\����=F2ќ6k�$]��#O�*w,do����\J//lI{��.9�R�߶�g��c�F���. &w��k;��6S��7V�M������3 �_e�u�8�N��g)�G@`~Ǘ%�,�Ȼb�r�#�rm�#=�ү������5�ܛ���9#�6h¸Ӿ���=��r�?/�`�=�(L���X����R����R���ӫ����Q�MP]��<��ԙ��9H�aɨ{@���GzV��W��nٰg�y�ʃ9�nq�4D�_n�Y���c1;����Ô���Z'�R�T�p��\qJ����MM�</{���yIk���4��NJ���у��B��Ϡj�|�&2|�iS��(����0�w��g���<�΂���T�|׊���"�L����Qȫh����e��Ng�E|"����A��eř���f���#?���nXP��&�C�q8m�.l�ܤ=����F��$}���P�Bw�V�1��s� jP���*4� (���R)c� >���y-ǩ���g��X����}|�>�pf�����p�p�>W�,<�>�Gm�/Ao}�,(���½m0k��i���[�xD?
��G��q$I��7i*��=O��`e�]�O�Ӂ �	��Ek/;j �V�^�%t��㻉^�O�������G5s����ł�8$��^��Sg]�%� �	���H�#:�45��f��05o�7�����0�T8�g����t�]z1X,�3Mu����u��Ȝ��p�}��P��Y�����X�-%5�l.��VeU\�JS�-�f|�Tn���	�6pB&2�
e��֯�N�S���+��`C���;�@/�J�DGʡm=Y���r0�|���2�'�]��@s�������W�a�����yҲ}����X�9�L\�V�����y2M	���R�k	9��r��B��є�g��{�N�xaC`��QNgO�궉$7Ӟ--Bp��2�+l�r����d� {t9%^NK/v�5;�u�r��`F�,~�Ĝ���!�@��gU$�f�h�'GY(Vh��kAm79�����p#q�W�xb�8�����;=���n�Ϭ��� JtB�&w|u	����w�m�P�c��C}�Z�\���n^`���;)���<����+�bO��d���f�^o<E��52�j��Ȳ�4�ڍ�u�Ǭ�H���b;���,Ǭ{�|�5Wuz�\��x�c�2~zPj��7IX�'l$E��9|l��U2�Bn�Csm���t����v�~ཙ	 [�� �?�		4D���D|����J�ˮN|p�%VZ��9S\�<��	)��f4������}�I�1[��S_׸��/�� ���.����Q�Ϭ��e�"��p��.У����~���f�|li��g�G�懫�RTzϖ�Hx���f)pǾ�:H|��\���A�c�)0E�?qF@v��Og�w�4J9�]�@xo������
e��&�x>��,ˎ�(��?��^��l^��!�!Z�Cv
фd_�S�c4b����L���$$�Z<m�X����Γ4��A���r�M԰����.u�_�ao/���T�[(�����=��,k��?��1?��G���x��As���q&� ֖� d\-O��r�76Ui��y�����\r�ɸ��%I�{�A��������p2ң�.W�������uR�ӻ{�ַ��D'ù�1��0��3ϳq:~ݐs�ރ��f[��m��1���Kr�<��j U�Ot;.�[ ���c��"�A�xL�e��8����\=)����;O3�PQV����O�����GǶD�����7O���PC�C���O����E��Kq��������2�ϵ]�?�^���W����>@��y[,�D���z5�dp����Ӭ��9#��9��!�Ҟ���s��p��s�ַ��;h�?ЬT�q�P��)94���K�;�W������ؽ�X����Aw]|�F�P����,���?t�u�饣'-��ޤoU1(ɞ�y~O
បJ��~��%x�9�b�%=譂tC��";�rA��>2���rΰi�c���[����Y�Һ�Cu�z7���c]XbZ�Wv��'��[&
�l���4z�DA�!��������
.�>'���V�R
��-�5����bV�3�k������|';���r��u�8���(�f˖QQ�� ��q�X����t�7��W��A8 �)�時`�[�����ª�h�����\L���)X�j����TH&�˯[LIc�������ꦓO��rG5=��P�u�X-�xBiD�� ��[�fqu��Ml��kaNFv�"oϘz�U�����a9^��,��9ߴ\��e�^l@���>Me��VsI�HkJ�-��?mPk�yl�Z��0�\�����\�ٿꉧ�+�v�����{��,i�u�|����%}`!��()��X�wV�]O����M͎�
���v"1.y޺���?�O|�:��"d&y)Ξ̈:���MD�:ƣ�k9D���Ћ��0��0;��f�����T�O�i����p�����s92L����C������ ��l+V-�� ��4!=���@��j���z]Ò$�>���g;\!��@U�@Y�bb$�e���T�O1�����l�c�#��2Ǝ�8{
z���!������U\��
'yb��݉JM�oE��	�8ֱ�/{a�-���ձ%	��5ʅ2Yy��!;�m-6
?���
�<�ܺ�^C,@����e����^��@W�!��l���
��7( ʗ1+��%�U��]�Ǣ�߀�=Alh��#ћ"�����.��%�ڏ>��B�@�՗r�<������М��αO�ӟQދ�E2kriH�Π����58+��a�*tR�vL�ӵ�P4��2�Bf�ә��$4_4�H,�=���)	q!.Ь�XE}��o��îT�B��s��Ԁ������s�A�!9'��c��	�-��+��}���
�K։�^�����-��g���2Pg��6�����Cl�^HE��$�+}�Rfx�T��]����6z��F����(��Ӗ_b��(��+���S/P��Wy��X;sO����+)&��BaƢ��fcw.G6��+� FL�8�o,�h�@3/�6�|���a�; ��Զ\y���Db:��U�����&L�5�����6�1Ƀl����B/0K���6���a��jiN����˰�_�l��[<卣q�z�Ne�Y�8]*������PV�h������E�0BFF4`�ŽA�hR��;�U4�Ut��~�3L_�����#����pVt}Y��R9(�+� p��9��a��;���!������jPA��t8��[<X��'[���d�{��Րfn/�G�&p��b߅�뿽4|x���{�[��B�t��w��P1'1���v��UE�٭�O@<��^���i_in�b�-sr�$�d>�,ʿB�$g�uk9�_�=W��(���6Yɭ�m0���b�����g�U���1Q]@'�c1D�H��N�Z/�P2��wB��]T6�'۲b.�É_�v�;���!`Z#����)�L�g���F�	M�.����$M�a���h���#��D/m��	L/(^Tɺ̿Ah�-�=��Q���I=��J�;�R�|�>������&%��_u��s�U�ظ{Dl��R��eE�����-z,�`�n7�>�F{�N����u�H��ٟm|?1���Jo��K��d���W�/&z�ﺄ�b�|��rsə�
]P���~�*)	���Ї9�f3s�p�zEIȤ�0[ބ&c��� �D���JǪ`��ȵ�)�$yg�)'0B���ɉ[�ԇ���_qh˿P�ׇ�7�i8�N��{ѥ�����Y�s�<\���	[��}�$��X��'�1>�qU�x�2���R �d(@k��J6u�8Fw`xh���jj�RZ9J}��{]._*g��9Z��kJ~��@k|�C,h5��/c���N ��'�P!��/��/�N�+O�wJۡ7I��덃$�1��³L�/@JF�D֧��)�Wo�W��
g�V"1�o�\5	��a�q�+�%�S�7��4'K��+Puv�7E�;x�� �O�x�ˌ��tݖ�cٰ��1IN	mR�#�/�t.c���8��{V�olWX`���Mm����j]X��?8��y�__ب�p�,�)��8�0`��Z�������]Z�[��M�����`2�4Pk<�8�JK�J㼡��6f����1�s
d`P���p|����ymsz�CY�g��[��X���Q�� n@q���U��Âv:�)��s�S\���-�Dx�H'Y^��>���71AuZގ����fn�T$���t���̺���ORRHe+��!#�h���v�-�?a�Q���r�$Ǡ����5�}���*��V��6,�:���nx�a5�ӹ�B���צ��oPs'�L���}�6����.q�
��? v���U�fC�TcV�A�|���k����dS��=�c�x��QV6YF|�#���m6�ZZ��F�yX$��+��8���\Ċ:�/9�,��~FV�o��I��=A���"����Ʋ@�E`J����y��	�z�Q�e��	^�����b�s4����*Q�,����椿���U9'���s�ß�C��.��{���7!�uފ�&��✬t*a+-4�hwk�뀀�v����1�B8�9|@�,������NWP���X��u��Y��T�z���қ̦LOw�K:�P��k�ǌ��w���7�Ol��QmT0/��|P�5[�Z�{ f���k���4��q̚��0���%���`5*��qNO~�1&�x��w)KAqD��I��k@;�V����T�~y8OJ Z�M�����8	]�;�����f	`+�G���'d����� ~E��_r=�* ����c ���}��^校��"�82��,y`�$� ������?ź����Q���D��#'r�<�hJ��
�˒������gJTۮ����.0�`��2Y?��
�'@�V�>v?L��,m�G��T �-���*�ɧ7�v�ԥI���c�Q��[�"�8-���b��A�(ݲ���Pޡ�A8F��߲���0�18�)�������T���/-KZq��eʐǗ'�k�W��O�����Kc��_��,Ì%՞�u��8��8OQ�)v�Hb_��1n�vP��Dt:WV�X8��������Lג� ()�~d@���u��}$|�����zlu�^*�=I�'�(ԍb����T�*WZYU������@Ik��ACg �?���(�K|����蟹��5� �<,6xG��^n9�#$�� B}\��X�F�u�c��Gm���%0�z���tp�Be~�a0h�ȹs[�9Ƴ���2	f���tï���_�/|f& �ڹM��q���O7B�B��vc�+O������4T��Y�׌��������|�Pi0	|8�⒚WfU8���������柛�.�'iQ<�B(�'� .���Z�6J����<y�$hF��7�ץ��c6�D!x�š��?��W��@�V�l�������7J�.������E7W_x��y���fXT�7.��C�HP�؛����F�������OM�W�aE�z:n�S�R'�􁉎l�-��˲��0B�;�0����ax�6��ʾkv� |���6xG�֝��8�
ܽ5C�OBO���-x���\9���L~�n�f�s_Kr���"Ѽ�%��-��-�"ѳх�7��Uw١�%*T_y���kg6��p���  �q��*�W&3��ݠI�ڐf���r�L��`*��"V3C��0�M��v���=�ۥ̣'��j\�ՠ��Um�G����7*0?��[}�r*�x��ų�����W0Sb�Y��&�`/H���^.~̲X���%&�4���ۦFCz�2f;GXM��2T�������m.0,Q_���"��[swW��D�-�����r_Sz��e0��Bӳ�!��za�~���߭��]�P	[�z�0�'���A�wzP~��	�_��y������@��{���:��d�_i���T}�S�"b��,LUc��:T����߂+�s_�0Kv��.4�9���uc}��S���^�5��ۑ����h��z@������o�~u�J����ߛ�	�D��Bd�3��8�c<��g4	%m�6�VOxU~�Z{��������n����f��{��-.v픅�0��U8EA�Ո���?U�K�����'�ʄHј�uO�_1�C^o�����(�k���ۨ��Wp�H>n
v���:e$f4�zE�r���Ir.(�*�^��x@��~6�ņ�ëL��uZK��I���q�LI�Q�Ч�)�Җ��)c����M�]8T�� ���3Fk������M�K�.���*~Ҿ�ȿj�>��= ՘����%�_j�<�t��F>˔3��$j8�t�SBa�����bkYOkm�h�����������_��|�b��	h�LgHΚ��O;ϧ�a���7YA��"�����1�wl{�6!�	���P�^�Q�c�� ���߶��s���k%+7�]m�.`�����\tE�xes#`�����ٝL5[��?�*ڱ|T	'��39Pa�My_^USs�T��8 Z�A�1L�٪tLPm�b�E �զ�M�p+�5���W��jX4LҰC���s��(«�x�{���P��M����tKQ��Σ��a�	�~�e���{�&!�.J��*�D�;1�	ǍoiT���PZ��E�X2-4;��a.d'���⾍���*Մ-$c~S���dY���x���9߆ݼ�3�����<�HJz���_:T��J��f���dͧ���h��Ҹ�N�c�$V84�� ��v���](��#�d �I�E�Q��j4�+԰#m���aCK�]�����������:����-�D�����?}wg_���2T*G���z��s�a7���ݙ�������������(��j��y�8�P�}ȏ�^y�T�Y�"Yk凉ǈ�v�_h�#ǌr�s�c��s�� � �Md�&����l9(����@�0�>�7����D��f�r���h��nq)ቬ-n���`#Lc>�����#8j��HBj��R��j<��$�,Z�C���3��@D����K�D8 ��Ҥ�}ӡ�Q! l򶈥>܇��#Ih��c6���ݎ{<Z{`yPNV�+8�uD&��h��xS��6�M�&�����s������W��Qn嘎e�W��y��Ct�@���a�f��M\Bq�H�NP˒;K�I˔k7 �Fu(d��x]�;Ң%������	=̌���j-�P��r��3�HBX���٧��_Y��>��*�%LDuRqW�j���!�Ʃj��;���d3`0>x�)Co��#��7�� .ɘ��p���"ݙl.��ǉ
Z9F�=l<��'
@w��V��$��?���@Fp����y[���n�g����o|�)�zQ�8�<П%
p�b��%'���)���瓚�t��_�l�ރhw��s���"����Y��S#uռ��+i�۽.�SQ�y��AnKg�v��ԕ"��#ʻ5Ewo"u\��QɎ7TB��םc0;�k�@aYc���Ä��e���sxF��+��m!L�0�;f��\�Gv����[(�V�����&�}O�V
�e�e����1�,�Z�"+A��,�V����t���y6noB��3e���<��F������3Y�2��}$$·L'vv�O���L�K�r����W��W�loC*ZLXJ����
3DP��*BY�a�DF$���v`�}gɵ[��Ej��$j;G���WQ.P+p#����'�J�!��YP����5�U�@Ɏ�K!�� `���}����B�Ц��<��Z�����/@��8���[�b�&��䌱�	0�vv��?���a��d����U�(��;���Vl�b��uOÁ,p����T?ŵT���������TXzwNPi��5� �" ��4�r��U$Yr���8hc$�j/e��֒�r~���M��A�ޣLV�t~�&I�Eտ$�64Ӣ�|+1o�d����UJ{��x�}�m�FA�ů��:��tS-9����*�������9�F�N��㩬k
����v�!�`�P.�Rd �	̩�p��@�{�8��B����'��&�ǩ��!1��ٍ��G���+g�.��<�D<���dK���I����ZC8�p�?M����'}Z��
4�Y�u���hsp&p
J����K�̙�u���9���A�$^�r�Ed��}JMp&
i�6�ԫ�`�u�����Ġ?".[���g�P�ۋX^����c�h�&�z3�}>�7��HI�^<�S	�r��p�'VO�̷�g㔙��B���>��Qr��s�r�m����"Sf��3�����`Mb�Z���O�`�s�C��\�v��R��
?A��8�Uw(汫����>5A�v,� ?X���SB����\���c�2��i��sF�zؓ� ��`:+����Ĭsv���ʈ���[gY��$=^+$vFR�L\���ёh~�^Z63'�X�m��={6/pNBq�`ݦ��(zӏ��yN0���,��*_�����lha��:���L�#y��;�Ik�x��X�A��,���FcB%�-W�OwO�����7#�CS.��}�u판��'56I"�0qŬ�'h�@�,#D!�N#(K��w-�����IW2Q���%�ʖ	 s}[N�@݊�|�M�����z��j�ܑ�eu9�(�Wݪ���&�D�w�S _2��pʺ/�q'hFrPʮ��G��iP�FC=;����=�s��YZ��^+�=oP�M����Ř����n��R@��ޏ����(4ۏ/hS�`��Do��NZn�д��]k>�#�:"�w��S`��c*�?`Z��l�׶�^��~���~�6]��4�h�w�.l��B�,�����o5-�,pMu-����)����mf=����g�t�b���0g���{m�^�{��@vDM�6�>2w�
0��OqFa_���NH��N���.-�T0-���S��cs��[��-'�T�����~pmt��<��scv1���V��tga�`o�>�������o� �b�d�*�3�U�6|`�0��
*����#G3�X��Я@��6�D"Q=��v��Q�İ��2ǽg���� �^��/b����%�W�EXU��߱0�@�tBx�����$����.���z��*�k����|��i��I
C�z���d����1}n`�+ΩKk:��QQ%�cIB�je-��
D)���N���H�@��H�G�t��=s�Պ��C�@:���u_[Hs@dv �CaEe;Ԑx�����D�,�;BU��+��u�G�!��7�A+8aa󋰐H�徧
)"�8�P�a#���@��3��t�ch7�3Q��"�q�b�J)Pd�|yi�`�)�����^#s@�וr(�.�e�>פq�����@�&lӹ��]�. ��\��(�?#,)��������fz;V��s�)���H���D�3��Ҩ�ͣu�p�F�.-i���v[H5��9x^������-����ٚ��l"O8�Cs�w��iCi��?Ds�����A\��<K4�t�Xj�r�q�o�S�_�j�x]:;�80�|9�!9����r-*"�*�n�_Y ���xZ�CY+�5]���������}��?W�=�t�zc	}Jg��惌q8��R�U����sj���'��'���@�� �/��� �d2%�ܚ�����k?�i2T��T;�qWGd��!�WI�>�k�*Ҟ(c:Z�O��*v�.�>��x�s�=J���޽�$U�:.#a��u���:)���ml}��o.-�/�nvI:ٓ����1�����`�/��Q*i�r��m���$�%�nrNqߺ:]q)d7j��lnpZ��� ����G��&FD�a"8�%AIL���u3��%[d 8|�0���:�[�r�v����K{jA�5�g��o����Ҏ�e��m�dG��	;Ɖ�3�)��A[.<e���f�kS���:.����5���<�ˊ�C8�m �А^��K-Md��������'�/J#j	5�p���D�]��:M��p~�t^a4�M�S��Tװ�/CCj|~���%�%(��1�R>W�j+���:~-���g����5D�t�+�x��u2CI�iF5�m_��X�Z���r\�f��G�޳���A�?~e��(��_�ś@�_8E�c���ܹ+]��'�t���<���oC�T��b�e��Y���[QU��d/�Â;[���J��iu7�Q�mV�T��z��"��w �ro���~+@W�����y��H+�.���l�qϳR��گw|.�,�`�$���]ݸ>�pa�yK���|�b%
>��a-�μ�kc��i�~\0�_a�d)h#<71���)BLe6v����Q9���XQ鱒N��@+��5�m�&Qs���(�Zg�न���;($6h-�X��[f��izi�LQGQ\7s��ͭ�RnYN�rç�F���h���!�y�p��Q9�g���ޗ~OO���R��������@��Z���ω3�%�і��pN��$Ǵ������>2�f�~�l�Y_
� ����0S�rR�@����w �����m���<�+�4�p^�%:�BV& K8�c��#�� ����u�~"1RE��Ś��z6�Vw����1>(������͊���G��_]A�O�����ݕ7ռ�� ��)���n�v�{c���G%�v�����<�4�\��Y�@\�V�,�BI�q{n4^Tx�[�w=�/��G�+��+��`%��(�JSχ�#H�b=A�^�Q��U�N���u��f}�F��7&�1y�=�,`L�r��cx�4�m]���;��S�j��r�x�e��f#(y���9�HzB��d�0�3��
&,ǝ��+S��%�hvJ��c�-Q>�"����(<����s8�-�����L�<��y�g�FX�]*�P=�z��qY{C$��wvA�>���HtY�1*=
��O�z�������վ��_�Yw���M����^�a6�t�'gY���z��=�u�� �ib�g��ty��@��ϟ�W�a����r���i�?�z�ψ��=�����'wAt���}�;��3L_��hb��a��ʣ��	����P06���
	��>ħ�;Y�ȯ�C9�� $4'A��6�?*�G"=q�_ڤlc��rPF:�:ǂ��Ψ79��ٓ���܃��.�f�1�>�Y��E��N89� a>���?��Ϳ�a�.ВS�$x�%��ݧ�uĸ�_}\��� ��Ҡ��ҹ�����ո�o�Jع�W�y�e�ޑԙhζ|�v�XE�j8Nl�Qf�f�81�h��:L�:�V�D�#f��R�|ct&�K�",9�
�فM��H�"1������Vmu�����
^4�Z<��=�e��Q��M�$7�3�_����6Cx�
��;���G/�x|�-�Ԕ1j�ݫ�lҍ3��&H�:����(�l� �y���W���%<#}3 �K.��.�����=U�'8cp��Qgi�^1T��z����-�j���a�z8����&1@�a��(T�vt�/�9X�ӛbk9W_���X�x�
\Z��:1SH=K����=Ƈ�~��BE�2l��E>5�X���Ch�&�0�xj��Ĩ�<�-˷�)�-A�<��=�����#��u�ځ}�5�ie�W1'j��vףϚ�	�;	s�-"�
�`ǚWѽ�ɟ<^G���>{��T(߉���cEuE����a6.�XD\�n�a5������@�����n/�$𰚘�����'-�u�㥁2��p�^	�#M�)4ٛ��42�=<��"F�FA��t��X�x��|C4�4� �W�1 ��� O$�}uS��:ٙ�9��7EI6�)vd6k�=6bGI�7n쿣7笸T�(o7�Q��&h=�h/,�"�����;)UʯƼ�`;`���\2��t�&t :�DS���^�'y#�+��O�K)y�|)��ɴKz������'�;���(�)<i�`���1�wr,�B�H�`�T���*��n��{�ݙ<ߦs|���c����^���uI6k�o��y�A9����p���;�<Y�\y.��ҳ��~2Rp��0����6���4 |���Β�Z����+�����R��ɡ6x_d�{?n��Ӧ][�e5��'�8;��T%O ^�Wۛ�E�ao�K��
 ?P��K���-f5����;-p�R��]ܳA��k�ȃ�P��F�0cA9������l�.�Va�Rc��sa�`�w7:x�6v���#����U���>��̂;颇�܀�~�^7�h62�5�Q�
�}-��3^�`�ܸ�a�#�:�>a o;D��.n׎����_;���@�ug��C�`�lnَ�.�]dD���BT���_��{@����Px����c�i�e9���W���J�v���#��]c[-�M�b���>Я[Gh�IO>���k�ኙMō=r�c�{�9���I�Hҡ��RJO X�i�P��P�B7L;���([�����M�
`�j��瘖��'�i�(=�^K<G'���P��CY��G(4��mxO鎵	&���m�E��rz���~NHi�I�]_��$��G�$�x�K�B�s�fjך���d��B������D�\u�U	7���w�'�d:"��1O����~ۊ���⫩R���X�y����y�C�-%t)�'9��o�a�����;�x���K�O`�����5�T���*w|��6�,�P:+3Ny(��/@�A!���J��%���I�`B�_�9�XN�A�smrW�X@�s �\��}m��`j0Hy�=�d/0�.�:/(�/P���m��,XP:�-'���Y��y�8	��a*24����5��V�*�w��х&�m�c��l5#�����td���H�x�	H�;Ñ_���(�%��_)�74D��jW�>�v�g��+R�4L�V�����+�3���l�x�7N1��:;�Ge����������*�m�KCH��G;���4q	�5�5(xh��5E]�
�ׯ�%S5�Qx;�PJ����(��r.�V�r׌!�c-��J,&b�GK0�6v.�� 洦B]ꀃ�x�5��|��{���g��+����Yc���ѓ���:�]%gcz�V����@����>Ff��3o����0��7mC�� &�"9.,pL��NbW`�L ��KVZ��_�С���=M��4�HU�����cOً'$hju��vA�� 6S}�΄Ւ�R(����rFV� �>�5y4�9P���y����hg�b9�O��/_��E����S�6Tj&���$Z��(�VR��,4���Õ�G���~KRt�R�:��vs�Cv+G��b�q����vzX�O�;	-�~h�G�%�����< �Ưқ��"Cu�r��s��x[�2ц��7����֧�c{:0ɨ앀	K�$�,�F0u>'l%PH��Rv0��o ��p���ݒ�C%O�,
�ܢ�j��6!4�К(��eJ�[l��̓�pܙdgWW��P��U �\�(M�M&߁��p�KШ^_���/�������x�t�c�a{~�]n�����d�&v�ڨ����K�.�c�9UJ��++��H�	m���L��]�
@eS��z'��:�'r�Dx�4N)�i4D�G6�F$Zh��.��XL��F(��+e��ʳ¯�^AWi��6�<�o/�����ʹ#������tt�3��kCDwhO&�bG��𷠁���Q���*��U���7!��� @=�m9��\����{�.��"��9sB�T�������K���pL��B��(���S=�X�(�C5�R����e��~�O��!���g_�9�J���)���E:�e�y{�e-�2����;E�~���yҫ���J�:+�G����TNw�Ts����tn,�s��6�t��d�]�����P��0��bZ�hb�Ѳ���0u��A�I �+ ��$�KvC�cЄJ�$��j-R�ZGH�V}�T2�|��a�]�m���b�Ύ.:�m^��\�ݷW L���������l��[sZ��~Y������8���J���R=Z�e�����Mhg����[����[�2NN�]:��!ːnF$��h��͍O�=.+VXq/8���C.�]j�D�@�Q.�,/+���04\%>S�-��'�A��D<*$c�?J�O�]e�:z�Y/��a�;�}(A�R�n,.��7#_ w�/���h8:u
.r�áo|4{��"��Ln �Ib$�?�D&2q��2k���q���:o�$�E�{�J��0����W$�FU���/#����!s��	�cg�HjN-�]�[l�d�m�\�j�Ͽ�Io|�R"�g؉�)����:lp�S�/��>#��qb�ǅB�ъ���w���.�(f@�w/6�j�~-��*�����/���od�~�����:8J!���.����`հ�]��������c�o3��W�f��VI0ҁ��c�f�/�g5�'�+
 �
.��+!ˬ��V\���p:��������U9�{��Gpb윮`T��@�o�/	LJEg��mP�?	f~�/����<�w��w?x~�(A:=���P
���Jr
��]�_�q��l�C��]��ɪ3~��"Xl0P��y�i�-G㨏O�� �"�b5dM�a�⼍����Ħ��f���J��:ց.p�i�����[�>(�Ȉ�ev���p�7v6���3ǔ�H��j�<�|�q����!BC<=����UH�W��9�X��f�f7�൹��PϕM��N��Ys����ֽ�La�O�d�=W���%��ж��1�2�Qsբ����s��@�Z�DR�+ӵ��V��+m�yka�C6�{�-d3�|[�H�?R�,�*�8���?M>0�K3���t�=�=� e�׭7����j���5����r���d���*
靁�|j�\�b����ؽ���n��a�gagQ��)I�S�Mf���
sbM�\������!�i��ؘ��o q80`��k�)�(褯`����TY3r�H]Ϻ�"%)ήߝz�l7p���$� 	Ԗ5*��V#����U	���3���AuY�E�+1�{t�0;����� ��k�2�pY���v�q�:$�hSķN����Y�Dv[:��sΨD\�ͦ)pw3�#mY��ѽm	;><$���2nCm0����M`^�y[�X�����̷������y1�"�Ub�|d�-��CBg��Fvt�v�<��C�T��/����ʈɏ;1�կ��!]m�d�/!fh��]���6j�2Y�|QW�sR����I�u�i��}���s22�}��A�S-�N��s��0���ʞo�L<�e��-X�s�k\t1s05.�>>�e�n!��E�Ir���7��.��7�NۻL�ˢ�\A8� �X��L��AP�b�QJ.rz�{�. ��w�u�-�uc�n[�eG��oey��Y���ﱪ��
��I�G�,��s\��}C�r�ώ'z1�u��eH@�,Bẵ����?�-�O�^�W��+5�Yty���C����m�MNߗA�a4Tu��� ������ �C���e�3��xt�;F��,b9%�O|��g�Ҹ�����el(�������؂�ϲ�U W�xl|>������p��;���t��B�D}�%s���,&i<ZM��I���xY3"��,ǭ�I�,!�I8���:`v��H͈�E�0}�!ՈC�+v@���!�bl�xre| 9��[X)jbk!A��:#0��\��	��xaD^Cu���ЯZ��������2����J|�M+e }�V�l�Eݒ<�f ^F���2���Ot�E��!~j)��'`�����o��>�lv���:��wc&��}�S��hN*�2�	#�j����$U=NqU*}wQ_,#ܯ}$�>������Zq��D�Oڟ�����PY�E,#O@L%���һ��i�9���-���`����G#c��E�Y0�C]��<�C���1�D�`1���||���)��<\ �M�7������Mz�9����q}(�dş9&:�ی6���~���R����9h��@K���(��=�u����$�m<*�P3>'�Gf�Gn���~�����)ˡ
�"�9���������~p���!�%�i��̌ɂ0�d*�^6V4Y�q/��6���H�)z$N�c�m�=4z9+��˧_"P�!D��=e��ol��'��}Q0{�]]d�(W��鵷*�čy�ٿR�H��W��I��AW%���2���$�����U�5*�џ�UA����}&��n!���24,�G�:*�5>'&���B#�;��Rm���9i��& _N�����Ǣ�k#��rz�}ɩ��2��G�Y-�ΐ2ܕQ°��S���W5�^%�>'<G�� עƾ���:#Xٝ���f�Nĕ�n�љ�)�E�|G�����?�M��/e�UiwP���q�z�+xE�i��Dt�� �1�\�n1�{���i|��{< #�r�O*:�����������ۍ��q����޲QX�l�s�l�h�k�N ���(,�L�2�>�x�چe֮�}CH3�c8�C%@]
%8*n%5�u�|��z��K���P�4M��e�moUp+a8�[^���-�
׿���=ۃ��V��W���C�vCJ�G��h���
��G���e�i2[�#ev���l�S��P� �������2�!{7hu�5`��U��W��Zf<�f3¹-�D�Q����7���Id?�&����gl�nB�[�pO�;_�����bFe��{ aǋV=����'�PD�.zu7��2�]���}u|���L�Z�s�uLO��!36��ВC߹3���l3���s��B��sL��8�iE���ze�������)������,���7�j�>��Y|{�We��q��}���+�������)܄lB�+$�аFv�]���gq��F��wx��������B�M�Zߎ�ʮZJo}�d\o�{�s��~�R�|(?��S�&f�����S�};��#sƲn��v�,H5�l=��P�(���a�ݐ]Ɋ�y���K���-X*��Q������a;k�gν-}R���{8K׎������KH�� ��V�rs�� =ͫ�jU����EO�V'������Q������A%9��,���4h}��il��z*L��>ݬ�l��.��1�ЍR�!�n3�r�l�3����꿌(����ܿ�]Qa)��8����|��'�� �"�z���%�"�8P$foѺ�����^�5F�'���g_�J5��+����ƥ[;�i:�P΁�\�zP�+�&��P+|`ٍV���D�ż�q�N7t[-a���p\��ΫB���x�νZ�*Uy5�� �Y���ȫ�Jȓ��t{��m�*��=�8��}W�;]�$�L|��s:��#%�F,�B��Rի뚊N�������#��RY�*vVͬ����A��� �7r�n�b�*�3bL-�E�;d>��h,����	��3XN��YC���a����8�#����ξo��]���Ur�.�i����l�{+�3��v�g�vu�)��V��a�� q�`WY���M��$Wk5*����\,���y��	�:����uj���������l���#��[fWZd���n��V�M�q�k�]�'���A�9k�!��*φ.�S���)ڲ|��č]�UQ"�=
6 ��d�����N��y���d���v]���m�� ��y�w'���.��%g�S�l���^�HJ� �����g畑sv�n5�8��:�v����nFx�2���I?���ۥ�ۗ�\ƥ�����k����#�f2*�KV��x��,N��wk@��6=�WU<1�0�m��'�@ʥ�[N�KBl��V�o<FӋ!A*��N��q��H��:�I=,��'sF�10�[<IDd\q�N)��װ��!�	���;��'	�A�\W��A`Ԡ斌��1�β���ށx�	����t�G{3N|��2���AݩWT��x$��X
Z];& �ӌ�i,���oa������1Ϧ4)8�R��SA@Ҭ��e�"8`�����8) �Q
� m׬%t<��򏶰�؜^��|�f�lO��]�Ά{7���qOf*;����� �&K���Y���ss���J�o��n:��Ĵ��T'���Z�@��
 �kw]��r]�Q���B� s���ʻZ C߭_��P��6�&_�ټz;�e�>�tBG��.�%Py-mP���oH^�~�h��p:��2�f���Z��r��0B��a��j�:Ч�qV�(s��P�c�=	w����p�y~=\��[�p���[]�d�1X*�˲=���F�y��]��,��~& [��_�y����Ml������O,ڠ5r�
�$P u����p6��-��y ��5c|�6��쨯��X\�6P�v��I�_��p�|�	h�g��Mm����QH%,�� :)��D�(~R�p�.��܁��'J�*�3:q00�r�
o���ގ��/��&)�󏫧}6�Q��՟cY�W}y_�r	#>�P��'�|gF�%-U���"dK�oK�4��U�պL[���c��1-Z�r�]����Ȳ4h��6��UU�eO��U���'���#<�L�
!������+�;�F���Z!zx^����[f�he�������ad֚�¯�[~�� ��Sy�k���@�7si+w[�=��ot(�� �L�x�)���}r�i�TvN
�}��'j{OD��ⶏ'^��-��t�:�(�Sc�3h��>خ=I�N���H�(A���=��{��]X�ֈ_��C�=Z!��2�PQ#����A����8�ky�:�N���=!?a�������+�zZ�X'/��2���E����*Gs�֨����/�<*JB����q=,a]����|����i#{�c~Ϝxߜ�D�w7�W*�����v�V	����J��֑T$E�=DA����^�_3�.o˭��vªI<e�o�*HcƘ�����q�<7�AsM��������@I��j&�.[���@�����j�)�4��ɾ�4XO}��� ��}x����J���_�/q��M���G�q�b�ِ��f�,��T�Hג@�R�V��k�@�0Ʒ�5S�>sBJ3�j�D�'��5��3�A�	�E=��WX�>'߃̘�aR�5�Y�
�̷d�7�kZ�K@��|�|��csx�n���������SU]a&��C�0��1��H��-���'
��B����V��4����I�Pk8�a�B��ԅ�^�|2�m��[H��q�Y\�5�y�=Rv��/�%;��
�T�:�Z�n ��,��5�J"���1X&�7w�;�R�̏�1����w�o����
[L�NڤG��i~q<sa��|Н�����/ ��b�Ad(o Q*����Ph*�5:#]uE/-a�B�+p��l�E���o���o^��L�?������":i�h��U�'�?���w֯F7UN[.�{S�R����[�N���U� �!՜��ޱ�H�$f\`)�_�<�B>�h����%���]1��
G`K�v�̭%��!�i��L�^\?aGcּ�ť�uE�,�b7@��U����a�_򭾧���C� �B�kR��J_2��>|����#�����)�Yb��ܻ�MS��&���.7p/U�~|@�+�J;��}��}�7���[���_ 6en5�]��IV�w �S�^D�~�t�g�����6���x~��~���d��r������w����0A7z�1���x'4���ؙ�X|i��{&�/�f498}�Ku�������g�q����i��Y�m�&�
�ң��ؐ��h\�Ų�1BA� �inɐ�D3VqiȜ�D,�3A����M��:Ξv/�*��m.0��*9�ne����\�Udc�%��@2-��(jޜ;�3X�ڟz������X-1x:p��y}I����Mo;Ì=)�9qsm�� P�GT�|�]O��I���_�������n�1??��Ƭ�KN�M�D���z�0�:���+j�����_v܉n�ť����YSaY#CЇw�Kފ�^3��m�b��F0�0�3#U:���]�&(c\_��B��a Ew��{
�RA�����uC3�I\��m�]���_^�XRVx=�`Xw�WΛΘ?-�r��m�c�Xĩ\������CA�V%;>z�-=Ҳ��W{�2��%�f㢫��V�|��	�&��ئ��Û��A��C��*F�@����*��1��CT�sg�<��m]�2�C����A��~��n� cB��G[�-��ʅ����E�a �֌�.#���\�d��ֿ �;������� ���B��j��R�{:J�Z���o�9���v0��W��9U /f� e+����8�P����^��Gi�<��$���z�G55���E�l��O]�
���v�`��9�dYXQ<ko�����SN�RS�zC�,���m�v�5,�~�����kq��A��@�	����g�a�m���#/�/-X'`K֥"�V��Pqqq��.��U�:Z?+>Pw��i6v��rͶ�zd*���W���kr�EISe#tV��X�� q��jzQ��k��˧ӗg�,�d��A0�c��|�c���i+l�W��kf�_@�u��v�R23��]A�*��m�$1	 �e�Sc�ɷTH.�F	�8T�b!��HMҕ����J�,?*۵g� ����#w������f��r��؞h�W�����B��	TGv��Q���R�sث$O.�6�P�;�}��f���u�Q�E�E����L��$՗!�CX���f!��Qs*��}?�XyE#�\��] �H��>p~���+�Wq��aN��>[�F�.:>�>_u֡
l���~���<��:�����3���f�#�ˤ+��D�ޝ��g8���=\ �<��#��RQ�$oX0�	����KBK�I�'�p��<,,��1u�qfZ�x?����J>3;�O��w��^��Xx��Ċ��̽�@Ia�ly@���@G"̈��6����4ߛ�K
�{G��@3b`�$|B�u2z;Ű]�#�� (�#�$�ޒ����5C[�K|OF`��-�>��YiQ�f�W���s�t�3�)�7� �t�k��V�z号HN^S�|nG�&oI4�y�bT��bS���T��LH�3�"��Њ�e�޿���UQ1U Oֱ�w����=�&ňu�D�2E?g}��KӘ��[	����]�Z��d�ӄ�PR-���Z�YJ}2��������3w��0~��SLnpJ��)���� ��Sg��;L�ܢ����#�&��-��7�����y����0$ɡ�r�I���]�0��<I؝L��ʌ᩹���sX���ԏ���M�[`x�獢�:JU�:u��"�H|�d�u�gR��
�V� Jo��ʣ���56yzZ��� ���!��]+�	�o௏�C��G�젢g����e���Ù�'(Ì|�WL�����w��Q�@.�B�9��䶲/3tP�M�,���'���p,WC&'4�S�qw���e�D~6 6��{m=���H���˓Ek�c<��o{��ՎU�j��|�So��
A%� 'CT�_�)�e���1V�';�a�`���@��&=s=*�Ĥz��ߺ1[ �9i�}-�������ȔF�p_��a=(c|��}��ϔ������+Z� ���X\\������������]3� 1�*|�6��=�P���<"bFywՎu߀N<��k�����,�ӫILR���s7m) ^�o9�-��9��Q���]���(B�Y�u�a��5���B3�=�A�Nٚ㚴�C����e�b�<�y���cQ��zR
r��|��C�	�<XC����z5�.��2K��#�`Ţ�V�k{u}�E	���?)��7Wf�4��b��<��8F�.K���a�N���R������ɌP��x��.�~;;�G9+��ͨ˲f�m?���_`��Lh���1�����K9
�N�T��)7���Վk�b�u�SB��)@�d�֦�b`f�PS����xf�F������,
,�4�U��b�F�y1�`�u��1}���juk@#)��-����l^�n3��a<��ߐ�23�hL@!��3o_Z��:��^�D��.�\b�*_+��N����WQæl�<2�n;'��g������"����k>K�mr<�!�yzE�?�vS����:X���˼z(������q��U�{����	�g�15�{���5ѻD�:�l]�ִ�+3���0�Ĝ��5Ѓb�.h�EB�::
��G�ֳ�����.<a2���V~�(��%���<���}+Fvh��V��x��W/�\hg4E-֎$� �*�Z�}f]���6
nħr��pC0��'�����x��b���α����T����������AJ�k�lX��c)(B��C��(��r�ՐJ5������lq�u�yTle�^����0��R�CD�����K9� �1]�������e�|��������%3�[��)�x�d��P��Rֵw�������X\���m�7�o�<|����J/p�����f̎X+4�$���M����3;��{�i?"`B'�G^�:��C"uI+�Y[�h�aț�����?�`?�M�L?��Z�����5��Kֺ�1������Z���bȟ���"�@�Kc�;��AĖ�$�.Vk��	���G�M��u��o����RR�
=�U+�2��t�Ww�_B�F����q�5�Vя<)¢�7��m��AI||�A�A��`�ԯ���Zld��n�ڶ�H�X
�LI�߸&�q��OrUP��x�`��hu�,��o>w�B�[�jp�E��0Ԛ��r�IZ_��%�9�%���h|�����K���̚��˄�3A�D�m��[L����v��*B�e��C�G3т@�K�^���}�l�����x�y�r�-��,��2�*N'����69�a���/�?��f��7����J�l���wFL�`Sv��/n%�X�u��4E������h����d�ɑ�?t�^D֖0C}�g,A3���3����Lpi�p�M��X3��dm��B�4���D���BuS��:��MyvW퓇93��W�6r�V-"�a�S��a���/�\���Sh��e ��l,%��]�����3���? ��ʻsg�]�<Qs&z�bFQp��X��;���(1�����d��by��'�����rTh;s����pʣQctw&:aZ�\g`ǚ2^	/<u�5�Z=_��9Wrc���`��4)�-{�*��f����D�Y!(�|�ܸRA�X0�R�MP�l�ݪ��	_3�I�4
몯WX6t�­wi��<��c�ɦ��E�C��ᆮ�)WW"���,,x^�Л��]:�Y}���}���t�M��s�3��g�F�1�0˂����C�A?���q>�e�6�5������'�m(!_XY$Nׂ�G��Ӈ#�%l`т��MHB��H�$NJ�9k�xYK���ܫ�Ѩ9�L�&5btԉ��9�	��X�ҲB��2�Q�2�u�\�Z�nJU*?���<Ǣ��O�d �@W���|��o*0�6QX�������7��	"�HG��l.`
J�],~��*_C��	1g 7?�U��T��!wv��fm��|�[E�\���h&J�IG�OG����Z옩��F��-���B9FvK�E0���j�v@\�t����ƶ�=Ă��$z�b����q���CG4�j������V��B���aui�4=c����U-TJ�/���Q�Y49?�΂H��8y�����)�����r�`ԅtڬ��iT�^���` �!6����vK�m AI4,��'	�`��� �l��[Rܙ1V�{
f�H��!J�L,ҖU��\�v�o|�72�y���u�|Fv��8&�,&��Y`��4��cAH�
��9]9{c��s36w�q�?���I��~I���,�2M��Ր�����f�V[���ܝ8
��IL�$�W���8�u�[�3tC�b����剞n��O�6�z��p�5�(˳u;ЈF|c-���;|i+l;O�18IQ_o��y�$K!�6�q��>�@�u��=ZF���	��N��X3��/޺98U�~eΆ��5�:
\Ԟ�q��<ں�˵P�H���HTl�'�I=�6��ʟc�T�-dC�~>��3l�f��d�fڔ�-Ѧ�uv�p�wM�w�8�Ѹ�l)GkT�K�ʐ���\f<���d�<��Dd%2��AY�P�'�C\Ζ`
@@4�s��;�����#��f0q�u���n=� ���a��_�(;�cp�9�!g�#�y26�Cߐ ����?��"�'|w�{3S*��3Sz2���}��'�Ψ�%?dМ��Ai�&��~��>PK����s-�{��p���3[@�ɌJ�,�˩���?ܹ.1�b�����L���J7^)E�m�X�?���}Ni\������0�K�� �*&�e|`����
����1�01�{�A��(0��>[W9��ƚS��M���Ф���'Ab8�4���i��OG�)����z��z�d�;[N��z�8l������Z? z6�q�o�k=2Ȟ=��9K)�;%W+P�k�M��)��A�i�}��,����  _.1���ɠ�L ��\ԍ��;�Ԍ��y'��)m�9�^D���a1�����8d�I�laXћ�����i�^�4����Վz��\5..IC�%��D�]ŝ�{��e����
��c�$>k]��4�?�\�������U��w։zc��k���⼐���v�u�����>*��s�F\��[����K>
1�a	�!�Q���c�(/ �y�V�Q�)�wKp���
D�fl(����_(�Sk*y3�lw��2���ִC�v�Lr�y�W0^� ���BYL�|�=K�M:����Dz�u�=�5���
[���WVM��$�"�,�ɿ��Mq���m�}dV�A$��O�/R?��L�t�!��f�4q���h���9m+�̅�HM�l��)��0�@�J4�G.�����{܋W{�\��A2�VFY�M1?��2<�	�ط�,�r�nD��Sd��D�f�^Mo)�Q�2N($���,:;��z�<s�VM9�6 �,��\��0�u�a�x��:�F�&G�
]�t���<�a@;�����^+IC�sx.����a��qN��\�\*�xt� x�IP�^�@7�y���~ӓV%��#
p@�9U������3~��.��i��`	y����~��4c�U`�G(�f@S�u����q1�ۍ��{�n����Z��ϟ�3q�ki����pt#�R/���R��t�4��Q��UdV �ݒ�$��W��ѐ�*y�a#�b��4�v���DpH�6��ȓC�4?(�i�"�c�c�^���:Q�2��s�Ӵ�껃������G�7�@�֥��"�U���8���a�B�vb�S�>�w<�)n��{On]N�J�e� �@�[���'nF��z��
ֶ�#1<�*���fz�#@&Cj�{s\�vv�E�>*Q��?��r���7�,\��\��Y�鄯/4A=�Qۀg����&�ĝ�����p/4���u��+?�Y��C�_$/�K>)��@�&O�:����Cr�x<��HTi�U��b��]�'�Y� B`���5)��3������=�+�بF"��_��{�-��?J*�A��0�e7���1OHL�
���[�V��g�ȭ��x�|�I~��[�&�p��8��C���c��[�ls�Fm(�&΅���{j_&�%�>o���<���̷�FH�O�����M��^���t��&_e��Ƿ�������Z�.y�g��"Ă�xm��uL�S1e��	�"�ִp5�7��R��Y�`�2v�D�c����@*]��L7����
� ���Q��"�҇�z,�;��=9�6�DQp��V�Z��a@k&����c_�Q5�Z�qO�����������߷��5ɕ�]�uP���pb~A����J �[�5ݒ��� �x�A�tR��1n`�I��l\?.K �V4�������v2<�ƍ�T4W������8����r��j�ŉ"%l�j	��#���)az�s穟�%�6�Tn� �!O	K�����}��S�� KQ"`G����W#1KY�aU�Ns|v�kA���'�����}��$���+�"��O�U��D��h�DYtx���W�M�����ׂ״J�7O���N��]@
�uG7�¨#�O����Mpm"��<�U\�,���	eK����3(�R���=���=r�ܤ� Rݲ)�T��޼�\x�����4�R^=f��bYD�|f�|�v���|�V�ژ ��Vx3�hXB�ʠ� �	4�%psoF �o��Q	C���|Qn"G�����[!�1^99�x��1t���`&�C���H����N��_�Z,��o��E �Yۗ=��bN�TB�9�h?	�7ڟ��t��M)��7��/�z���^�r�e��a��\�8
-�"�s�l4�G�A�R"���xM0dV4�´bR5��_����r!�����R�g2��P�
�݌��=��7�5Ag\�5��i� �J��Q0�>���F�T�'����-�� �W��b��o=�:�'�I�ۡBUn��&����yH��y�j9 RF+0^�'���3aA���a��|� �Z��_�.��g�I��E�U,���z�/��/m@����/�"D$�.ϗ8mW$�W�p���-,c0n���+�29��}T�����/�~Vn0��j"�C�J��`�0��r��[�C���E.�㓧�M���y/�d�� ��$�g�Co�q�vï���q�5-(;�W0�(V�TWH�L��K���0�6y�=wu���B�0*�A��_L�=�4kU�P�������Ԣs�0:�jR��OG
��f�ٗ�=d+c�[�x6�(0|���]}�4����4�����A�Օ@Q�+����#�s���aN~]��K���x��H��a�0>�=N�:m�5�S�`��"FT��$��ܱ�����Ą\�긿��G�F��������A�%���G#;0�ݳD�`h�>�腡�<���'ʔ-Ia�HWL�U֚��D�v}Tku���߹�`/k�x��b�I�H6����*�f����LH�v"�߸w�ԴL�Ц�x��/�r.�Z�Do�	��OL��&;�h�0F�o6��4R�! ��Zq����������-�Ɋ*w��~�4?�wv���
CM�Ez�XUl��`lr�V�><�K�_�Z���%-��QN���%u����_9F�Q�4��,����+��"3�i�5��b Joǆ�JE�m �0�pa��{<��E�d}2A�K*y��$]_d���qaL�<��מ�wb����"43`�(��Mt���g.nr���q?(n���y8��xU�
n����,4͒`���o��O��ٰs�xcΪXH����o&5�%^��|��i�;,a6��\�%�)N�)ĞH짧�ź��۳n�u@~Cа�1��' �Y�mſ�F��D�ưC!������hg�ٚ�+w��c�E�Q�[���8�猋��-�{.3��`FS�y�ٻ,\��ٻL~��b�g���*s��ͪ4�u�����K+17��n���zj���QG�F�&7�T��[��j���g��K�=�.�85�j��@}e�P>p�����j
�-�u�_���2�9��0yO/��
�ڧ�X�p`�L�b%�b%Ju��Ȼ��E��A�����?��k��h�Q�+v�{��8�{�N5�I�����ꯒy��k`��T{C���x)����%A���g?�.�O.C���M:O��-�:Q2�Z#~��s�!�s�䶾U�6��S���Ӝۀ� H�!����w����<��8����)b��~��h����*�	m*"���g�f6�Q�AW'��]�DUMB���Ɲ�b{��A���F@&|����i)_VE�C�V�DT�SG�xou���n����rp��1/�E�Ҥ��t)z�{�!F�˅���gK��vm��zuMd�OS('�S4���dv�]�����Б-S��ޡ���ڳ�aL�F�1�/�2���P�c92�� ��Z�o��	{Yu�����I~,�7��f�O����Z�!�|��ҫ|�ي���a<(�cF<}���l�H+!�	���!��J?k����b����K��f��	U#��?%�r�Ȝ��.%EQa����:?,�zz^�w>Ty���9�@J��bB��|.�p��2��2���Y�����3`;�O�8��	�[�*�z=/{��&+	�,}[@�#l��L�[�C���9�����S�i�~��b�{p����A,�Vc��?�~�#��C�,�k �s���I��k�	m�7�)�����{]�z��J�7���m�~O���Xp,e�D�� ��y�,9��/}�;��_rOh#��L$��ŉ,R���]1�cf*��m��ﾾ��ŉW���k\�����0:u����B��ܴ�]ۃ�(���;�42��.C���,P�E�:ʹ���i��-t$��!^�LT�R�w�i��>�=Em �]��+��vR�l�1��'PS��5Z-�V�-�U7h��+�ޠ���v}3Y��pD+���g �՜�'qу������]Oy1��ݤ�8�oc�៟�~|��o�%l�����(�rM��Ӧ8 ��{�΁U�$���(`�0����}��2s5!�Dn]��,W;W3�����4�$3�r��
Nj�q��`�����C�����jJ�wz������F ��h<���vӑ}�l(s���o%��v!R,$ػ̿w���-A�"'�O#��^T��@NIXm��_58	�U���&�����b��Q�N��ߔVAh�It�	�
�]y݆%pd˜UY0����	_��^��d��dp��"cc����D�YI�]�y��+���C�|�g�X�<�`�f��>@�[��HL�h	�y���VF_��_p+�߈~���>ؒÖA���� ���X�Lu�k����gu$m��R���no���k�N+ :�]_s���U=�w�&>i�m.�W�O�s�ds����##L3�J����P:#��|I��j�C
�$ͷs���rA΅�C�I gm�v�-���D�Az
b�d'%�x�+�FPbV\';�{Z}���,~ƻ$��"����=��AX:w~���Ra'�#k:�@��h��5q�.��f���H�n&"�(4�����S�BUf	P���U;b��::�� t"�W{6�;`��̞�G?�����&<�@��VaJ���C>�\�3s
o��tNޝ�&��0�ܕ��K^�Q�p�
=�sc�PFq�H.��7�s��9�|�]{�A�+����'#�=���h�h�S,T|ݿ�.����Dk贛�nOQ���P�<l��afsdIwCi�����_;3eň5;�q2M���� %�w����(���ˁ[�� "�/)&��9|���-!����}P��|:�x�x���[=�{�a7o�k\����zNƆ�\m1-�&��v,s�i�0NJ �ƸNat� ,���K�c��7��6.g;\����?b�FHN`.� �"�L����¤��R�Q����镋󲥈ƪ�9 ��֧��]�G��(N�ӨU�X�FQ��`�4;��A���wt����ϝ������ݣީ� _,�����=��(����Wp95��7���B4J���p��G4&�.�$�1���<`A��vR㈏z)�k���>��K�d���ڛx�t;�P�Uj~k&�9�d��c��A����?�2?x_;=c�qwÌrPH0��c
P��G&�/�3�#�S���{Q0����X��ۼM�m���$�D/���]A�ˊ|q9u�.P�)�(D�g+x��Z
�y���K��'D`��8�һ��6j����?����eĻ�J�3&C&�����M����,LR�ô$F6��I��. w��|H�ރ�� W�C^ٻco��/�](#�{^�&���m)�v@'���A�����H�c��7+�'�☙�Yʷ#�]o>�L-J�'o��
G�ux
�2�����I�DzI��@�V����ς��c�T��|�k�w�s&D��s��l� ��	��?��c���Xs�2�Q7{�8���[&�Mh��4�IP��o� 
Ah���w��"��]��g/¡�Y��E�މ���stI��.�h�`1�X��R/jmK�[?��&��/q����y�y���̖�{�ީ�!�3c��I�7um6H����U�-h����q��i���D�_�A�^���}�!ɀ[�ͨCi�S6iy��;/���$8��\{���̹���ŋ�H��g�`r��n/��0�nqL����B�oH`����K��v�A,;#~�=Q�G�k�b����L0$U�oȂm� @ʌbH�y^%�x^M;�k��!2�5��a�"�S����!��x���K�C��\G0W���8�r��珁�Q��m�#M�X�Z
��B�X�Q���<���dKM��k�v�]ʯ��a�ȼ5��p&l�h�a��}VW�j���_�߻�"�ÐtF��=v����Z���?D�0�i+Ĺ��5g�g����g�c�A'$??*�CJ���Cm����>ܾD ��؃~�T!�NR�*l�%��C'F��ؾzXg��=/i�+�t���OҤ	h��$�����Fmx|�W�o7���lə�q���k*��J�ȴQ(��3��c��Ū�	\���pZh2��q��N���i�� '`�7��+�}��<�_K���Z (U����h���N�pF�x4�̉�gv�SZ�}�h��P�`mA�G�P�ʑ%{ɫ��?��x@��-�ġ6 �މ;B�_��"'����*�y`SS���En���g N*���9�l$!��߃�z�*.��5 $O+��Gǵ@�k�s�������=Ȧ8�x��q]u25iS�^��P��SH�X��]���75����q�&K���pF i�/0Ӄ%�\�h�twD"�mk�T��'S����w��\�f�"��O���
wh�e��dY����P�!�|��(�퍐�B%��� �Rb4l*~Nd���< @�*U����%��aw�k$%*�keM"7�� z.�P��C�>!Q�JHED>����!��z9��7�7˲�V��G `]�N�����L]�$�)��]4�ʉ�^قdi�B{�Gj���4�z�a0�&y4�w��h'M�����b��ӯ�3$��A�cw��������{dX�qC���>��U=?��2�L���K��{I5��#�J�`Tj�[7|�>D�nX�D����6Ljy�=;>�Ne��K�,ه�s����䆗=,�D?p���8L��*�L�7R~}�u�s{���`�|d�Uދ��Т���4�E~aQG�湷�͛7e���;�#�Jg+���jV��bg<���a�v�4*N�)�.U�/X��Ly.D�tP�5M��M($�=?���{����~����2Z�������ǝْ��1e߾PA�.W��=��S���V�J�/!BU?I�8Av��U�w�:�����<q�P�:ӛR�v�OG#NP �\}j6����q>$Hh!^�ZP��[��]���`�_<gE/���ȶǩ�%!�'�5�0PQos��P:Q���O�� �����p���.d��[�$�T��ն���)�4����ҫp����,E�ȿb�ת�)�w�q�:�����#�>�rhG�i���4�m_��&����l��2�M?�FJñ���68�0`E�e�}SK�t�_L�s���΂VR������/���s�L�Y��+Ou;�b!��:U����N�����K�Vص�z��M�⋮+����2����sX����$��l�t;��-,F��^=����tM�=+��C*ǯ�����H�7�F�F���T�)�t�	 CH�_����qj�>ޘ�A��e�kHkOhé�V��\G��N�%�j�]='?Ğ���C��0�-6��	���_�E��/��Սzs ����!ϟl!��<W�ʡ��:��YF�j�dT��(�&l��G��T-���M�5*Ȥ+h}D&�+A�z�ڋ0���l6�6�t�9�<b,�ߚ��;C�������4O��\𘙩N�r�7/��۩�)e��`\�IvF�ԕש�Q�#J>��l�jx�����&)�M�����%q9�H�郤p7����n[��U�Rv��ؙ�s�-{ӭ�����̴;lŜ�="@��.�%���R�_���n����A���U�H�j[B�da�}��X��v@��W�\y�6z�(l:�>�����#`���n=2.KP��)1�U��ݜC��>���F�蒄ӿ8w��OH ���[o�?�ؿ]s�� ���<�����������ߎ:F���6YꗭV���>D1�S�
�E��6#Ւ:<�y�l�7A��p]Zb��Uh���*�I�w�*�~��"��1'��Z��� m<��D�f�fc�O�fn�޸5?w >����Sͱ��<-PJ�TL|�OTޓ 9}<�5_��f���=����������f��?7e�
�g'8�t��]7����jQ��g�	�퐤s���>��9����b�3LD"�6�c���{��	�.�f�#���cu���R�Jh����V�4��d�X�����;�YΤ�[���f�­f:���
L �?�]�v5;2���� "l��G';F;�\������S�	m�RW/Yky��Х����(�k���d���wU�w���"XP���9�A�2�0+� �U�ŕ��c�|ة|~x̉h>$�vՎ�t�����5� @�	�pF�͠�}-u��sX�|,X{��A!ӯ1�d+on�"<N��b��(�������̪y��Z P�v(�3��e�`CoD��@�H���]���v*��~�!�3	r5v?w��/:��6oDP�vn̞��}$k������k�F� J�4�c��r���D�K
y �9�W�C5ٞY�Q���e?韁�OL�JER-|��ݚ�)�����l۟\�Q��'��1BHb��
��'��怴#���a�[���?  8��@���	��U�C�ë�[8�p�ӥFCn�g�+�}�7?��VC�!_V�(lg��M�����X?O���)���'��	����i4�l�浅 ��-1-&T��-�g��y���Ż���ܱ�>�}�b�CU�K,��T&>^~Ŋ���&`Lm{�<m�D�]K����k�校�Q'��Y���$6���O��`�/n�J�Q���խ>��S�s���$��֎َ��vϻT��Xq@��h��?�8z24�b6Y�TQ[y��r-Ｈ���(۪��� �L��H�r���;b���{aZ��1u�!���K�A���$�l�����/��PX��j��ɗ~�Ů�5����B�+����,¾�z Ne��\ǳ��V5"4�@*�����m�$���~#�}��.�{�X�� H?'.����
j��U���2wW���q�:Y_��
\|�4bv-��Q®�ʊx*����z��p+�����]�N�q�#A���q7S�Fe��ĩ��2�[|�E��&�#Cc#��}5����I��~���6=�|ױ�DO�,)�i&�ώ�<�L�����M���.ׂ��1�=�DF�i�ъ��D�NB<xe'�U��:�9h ��c+<[�N)Jߪ�.�����{Plbħb��L2���/@-��k&p�E5rM�F@҈��"��H����B��#$�G飆���������-�/*�X4�V�r?���Ư��O#�8�ҼQQ�u�u�Sq.4�Cv=Iu��E���	�j�R���Iٳ�e�sǫ��/���%����aV?���|5(K����'۫WT�C�AV^9���CEe9��^a��:�jSq��V�
�/�7*��;�3�8��,wX�H�|\�QF����]W���v��� "ʞ D����..����J�Ӯt�|E�/�O�D�Ir��h�$.)8��-9�����j4\F�\���D��#8�J�d�LG�[�N�<�\U�R>�weR�~��tuq)���WX���+uqF��e�CY���h�^p6>ɜ����*u�	�M��.٭����9F{d���n��V�����-R�m�a���}h�HNcb^�ou�����/�]K�R͟�}�hg�v9�g0b��ԉH�US�j�� S �B��#�/vDZbk�a%�Y�Qp�z�\�QA�{��<cʿAસV���H�f6��M�"Z ܕ�e�;�i�Q�Y���σ̗:�.>��^��@�@/k�5� !�ڛ�!u����#�Wj��&��0<Ҍ���C��j�S���wϠ�m���ȌA>��<���d,���ن�'
��pPǮP$i� g:��xI�(���	�|�Gnt�`���Dz��۬h�.��L�B��`�	�����~�����ql;XM"*u()KײL�������-�k���~��}�PY�v�Ӕ�b:W8>w6�L2w��#�Y��ю	�SwN�I�pc��i�����������*(yB����8%װ:���Yz
TX�Y"�w�H��S����X�쐦Y�=x���;=�r�Y��6wE������hf;!�
���=*����P��R�m�x��\^
c�G���H��u�2˴3��`���Ig(Ty��F�}8}���%Jݦ�m�K�Co?�쮍�E�ǓY�J�VnᯈB�(�#w@�d)�X}ֶ�l�?Uv5�T�~��g����"W%��/����4d�mlw:�8�-4��D��h����g�����\bb62긴��y,�7ri��nk��7*�4]d��_������v�\��cW�h����U�n6�BCҁN�5������ٮ-�5�����,.k�Z�����tvP���A`2r��p�:r�.�������B�~�*	�A�O�+�&�|���+��g�D|�F�B�~;gH��=��	XPF&-�6����7>�Sc��[R;�$<��[����<P ��H�s�~�w)���H}g�������O��e�i 9�L��F<ܻ;#M��쐀�q�A���8�F-E�(z���U����q��T�ؾR�L�/�[��E٢��A;+�Q����<ɝ.����{*aOh[�8��b��a�/')WT@����v������<�뵽zI��i?UG�+ �����m��~��ة��H�/��U�H�H���e�<`b��>�}j���񼜬!�%�]o��D4�l}4|k���5�.�b47�~�bO4]��N�F:�V���l$�7R�:�{c��G�rK,�<{{����я�7p�wY+a��� ��^ut��þ󷶪5��&�=S�[�	�ަOTLJ���c�I��>EUR�Z7��З��:��*ą��:\�|c1�	���ɟ5gK�Qf4?;6��� ����q3�ц�����.m�J���^�t��aq�D�	R=C>�D�'�\�{9���B �d�$D�a��:�K�<�|�P���KK�X䊂%hϝ��{Hw�>1���kc��y �G9���rS�f��
V�WCS��k�s�~�ܥ
0��=�.���M� Y���Ef��y^F	=-�pV^�x��f��i��jR]j��$?r����!ut��@�	��<!�䩦+6��5� 6_����|��`�r��U���l���ʰ��+<Jo�_1��LϿQ�������!®1�'U`�d�P�o^�U!9�Kf��	]ѳk��m�P%�ף8֨6'a(6�I�t��}��|6�R��݁�j�c4XSC.$�o�
�)�`\�g�>�|�K�|'��L����i{M3��%�m���(�~�:w���\()17Y	mAV@KغՂ� ���HN%_I�=���Ȇ�*_Z� ��'0ɺ����|I�
a�&������y_�ٞ��|�����⤥9�|�sS����d#!| ���o�~v��x�6nIQ<BW�f 	���	��)�Ғg��䊖5���:h=�JP�pI���;(vPo�L"�$�>`�1����ş���N�RĊ�>
�/s~vWڒC�I��{%ی�Ϧ�R�r�_9f\?�W��=)��$��� �+H"��j�5�������:E���)@^��ٯ�0=_��?�.�v��#/�y�߬ j[�xU����(U�|��0v��)�0-��z�Hkrp@/�'�W´X%wM�P@ce#R'�)����b�J� *��׸F�V�J� T�N���w}q7�s��I�0�u�O7�B�,8�)lf_h��tψ-VD*��/t����.OZ�mlr�9��E������� �w��u=Z*.$�[�~�M0�
��sBxW�f�0��x-���p1�i��N�]�Q&��F�̀e�oz�ǽ�ҏTsU���'���p�g����R��EQ�eJ�ć�0��J�*8�o~��ث:�Xw�0������o�1��֋sT`�!:wat���_}�!枠��=���U��W������t3��h=������QU���{dB��4;�Y$�=&������]�̹���K���%h�N7޲1z1��$���Ԛ/[�]��J�/���N1����=�;�?l;U�xɺ�,�1�+��"'�k��|��֖S!z2�A��Cz�d���:�Y�Dg���:��b�E���T2c6��n�F������q������{��,
Ï5$�hTzڹ"��Y����8l:�f*;�Pu��7�{����<Y�nO=�E
���G��P��i�a�[�a�63�\A��(��u�n���1�����E2��	�e9O��`��F��s-�����q ��T�����"X�us/�-�F1���d(d>r�b��}�~�oqN�*����:l�8�bB���E�B�-����q���-f�큖�j���N�G��زX�e[F:<dj��0�Um#P� �;)��ZxsJ������~g����`���εjE��
<!֘�ʈy�vA�Q�Ny���]���;��v�|�u����Y�ϭۻk��|�w��W&q�3��"T��X\�~G�E��RciH�L<H7��Gm���4eNkI,u%��ӹ�b������lLZ�O�싴�F  k�����V�+�� O� ȸ��4;k�����c/C
��G�	���_�rN�n�u�JZR���I�e�.������w����Jbl��/s�*���7���v(t�i��-;�`�S�_�<�N����y{ҷQ|l��N�\�sp���̊�в'����M�+�����(��s�ܴ�Ҍg�Z5�vR�5��(49��/�Y�M8�>~�L^R��ᔨ���T�.kʪ���0@4���CIV5^���F�졑~���L�u���{��]D�v��V����V�5�2\�ÌUBsb` S�R�2s
�����I@T�Qĥ-y�R���F^�L���b
j��du@�A�Af����Ԫm�;���a�7��?���-?��b*X�]F�w�ah���X���}9�"h}Uj��Sњ{`2Y<v��r�mS���̏Vw7,�tI�~��\��ݗҨ���<��q���%��$H��>�?�ǹ}Z&�����&��Yc�uБ���YH���c`.u���@��	*�����8��
 �_����iYP@)-�:��U#ɮ��j�9!�u)�:0Q��R���蟊�}�U�Pc)���^%R����K�uy �l0�����=E�ofi�<��>\G�B����r�"3͍i����O1��
�'V8��HsX3�HK���W�� !Oo��X���i [ar��<9/b	݆~��������8�,��Ⅼ]A'�H����LQ�s�n��M(s�=���R�YgǏ��m���`�U�˰u�ܡx���sZO�jX�i$J�iAr�~C���!���ª��V�X�%M�t�NHį惼Xp�	w4Ⱥ�_!�fc.]��'��7=�� s�F%@�dzƁ���Z+l�e��Ȳ&���C�����y����0��i�H�8�)X_Udr���.�%8���x���*��ӣ}TEfj�CE�7�C�e��3Kݰ4f0u�+����z�x�I��ъUi��|Q�o�epp�Ȱ9��O6�{���˹yE&��Fx?>a���6*f���{�k����-����q���?C껚�O嘇�	�>Ds�|�Mi�1Q�/�Vi��[.�����`F��s�=Q�Izj�N5������������u9e�ms��J�"Cb�\�N����B�,�^/tN֮����7��g��FK"Ij�=�8G$0>�Q��I�d��!xA��N$�D�!���%�i�J���� Cc��jS���]k�X���Ƶ�ϩ�-O+�t:8���,�C<�=��/�K����_���K���(+�q1�Q��K���[{"T�V3�B�"� T�h�P�>���?�����6�Z�L���3��
��LUX@$JD�>i�����;Q�8?G����T�ϼ�[%͖E���kC*i��`�U����1K+sNr�M�2�َ?��ATf2'5�=!�6P��B!R��n�~��<�`�'6e`%qE�Iy�5�Qv���E%����>�A�sm�6@�*MAExm\h�Z|�)򣨕J`�sT�=�ދ���p���h����9��#��(���J.s!	",m$���2�T�� ��r��} f�a���K���0|ms�\�^���	�[��)ѫ"=F��M=�bwkق��դ.0����XGg��I�W��@�L�E��&�P@{����Y'^A	��2�����	�#���?S�ِ��5�����.]��f5V�l������<��r��:S{�hq��⩧��L�ZO�.�Ziu[&u:��+2��0�Q\�k�<�V��/��|ߓr����`<V��. 
!�f���)G���3n�B�]v ���(��ѿ��l�&H�Ϙ�@�xlJ
*1�<�N���<��5ݹ�JD[�e	��hR�)$��J#R�����-��B�f$a��	OC�RO�[���q���{���d��G�	�S�J%��v3Xމ�[�� �q4~.W-����_EVp�q~��acQ�n�w�(1������y��jD<����u�g^5��lu8=��[���y̫��ǼxU4�������otrб�(8���1��`�����'��;L��w��ש�v�]���׈���S�>�!B7���r��0b��_�����j_�Lnr�OSZ0��J�����>cy�C�_*Ĳ���C�5�b�j^Q����EF���ޢ���iX���E`��2� ��NI�[���zs�`�Z1RN�)������̗�~"��U�=�*�&���NR#�[� �N�Y�H�w�$�WHH�u���T-�a) z�|-6���
���^!*� �|x�T���ԑ�&T[!�Od��2�1�9JØ^��-*����=�Ml<6���BbsG��F?����R���@�<�[�W��V?��ؘ-<6�Ҝ��J��1�Y���]i�J�(����q^bl6��ς^{3e?�n�<����4by�IZ��'ea L�D�9��Ԯ��u�p�ed)}��M�|��N�~3�����������>d�j��%,�/�S������/ꉑ�K^���c!��x��)pe��-�tΒ]���=w�u�Jd���<D>:+0SM�W�\7��(<�&I����@��Q�P���2�pЧ�'�i�5?��z�\��Y�GUUV�-�/|D�r zr�Q�rI��{�q�-#��+��&�fj��բc���GGx�ͮG�i��g%���Q�~��GA��e׷ �>l��T�G�j�V=tH���#�DĶsٔmګ�}}7��o���-ܕd�t'� V���l��`�t�d����9���tA<�&���ցޝV�,�ٍiÈ����t��"?'��d_��߮���sj7�Fҁ4����[(�΁�O^��	�ty�-�z$�(o"n4B7��ҖB��[���f�����΃�c��{�0�������ĥ�6d8�	4�1 j��U}]�4O�s�k�D���qV�$�\�侩�Ǣw�y��ƾ��'��݋(l�*� (&^��U/��Y]�慻�,�>6Xl�OB���
D0rY��-cO��E\L{�+�'��K���N(�^S|=X���vT+������s��_3vM�!ą8����>(^=J�D�e���ZÅ�"uÕ��ϸq������4��wӍ�q�����o� w�g�*_~j����x��J�b�Ţ�7�޳�9џY|
����Y&�J|��N0%�po�,q��z&�x� $I.�_Ì� 1U�@����ǋ4Һ����D�5�ezUwI�ߨɾ/�7����Ͼ�)�L��{z����wy�̌1ʡ%����B���&¿����ɾi�ʇ���#�o��Gp�()D-b��Y�3��n�M��@RU�'�Ju_��<պ�?Û��ebe�bvJ�@����#���S=؄U;ג����* b��Z��w��	1=�h�$���+:�FyM�w�I���Q�	�PܱRwlҌ�5 M�|}*�ɘ
z��K�ͦ2i���7��P�.cls�Y��8��X�"�hf(\QB>��ʭz<?�a����gZ� ��v/�k�;�AԜ!�!�dI�*Mb�=Mn	��p2$ϗ1�	S��\|�H�پq,��%w�U"�F�;��ؼ��鴩
�K���f�4�N��J����s�x���T�W�J�B���?���@q�C
�S�jD���	��&�	II�'u*`P2��i�&��1���E��jMr�|��N��Cgbo~��$��!�&"�Kgj��P��ͳ�����+sWo�{uϿ�(B$�~�*����ũ�M�yՎ��|�T<�\��Q��:�{	���A� ]�B�5k�D��ݕc���&��՘(�� ��6d4·'��h	 1�"�!��p�%Z鮂��rozɓ�;��qo6�U�>	l��>(=����S׎�3�R�ռy/k��sh��|���(��$��{��=J��2`%���_w�S�������v� Vx�(V��&�3�5�U}W��X��*�13�uў��{�''t)4�d4yx>��RY_�f��Z����,]9�L]2�=��$d�'���pu�ŭ�&EbVK��E�'a'����"�WB�4�d�T0~}D;\ћ�Ǣ���n�#�����S.�4ĕԾ����q�{�%y�;��'�ve�Fo��NK��`�,����`�_�LM��='��4�7�%39T�o�f$�RҟT��M�IqMm��4�
P�
y�4������s=�Eb��~����X��0��l9a�P�g %�۫��B���R�
�S�oԺV��T���~�@�����M�,�<��k�g��Y�N�����e|Ƚ�������� ���R]�CJ�*�Ԩ��бA/45Q�}9R%+G��4ޞ\LÓN�ٓ4s�>wۂ^�HDp,�A^�g���7�΋@��:!��)a?B�D�:�FG-b�ӛۛ��0#D* ��1�����屦>>B��m�Mq|�}�ٜ͞��AWw{3�+R�1U�rݙҤ͐-hQf��o����fJ/������t,[��`Y���X�	=[���Mq������RAЄ��B�7Չ��ZR���k����
�xS����OV�U*��o�|�Ueض� UY⣧J�@|����?�+w��I~�U�;e��y8sJH8�P���^4h��@�}7� 4V��^ȴ)��'Xc�Bڠ骖@X`�����(��:�莺N�UHV>r�9cJ�ѶtA4��d930��d艹ʲ���,]���5͕7|Ml�by��-#]G�B���8MV*��v$������C�yo��(���� ��/�Ӎ{oy9<"��XN-��bSb옄�/����U�_��a��V�G���e���4;�|���Z�]�h�QP��!�Y�kv��L Ӵ1�H��R�,B'����;��?�jc˓-��V�Nw���˓���|.��
��l5|�x�,`�E��N��׺�,HKǩu[Qxhsg�5=�y�]@2�y�7�x����S�X����h���<t�
|[ec�1��%�|쇊ר�1��)Iv����%����M��+���z~�B��8S�J^O2 �W߫6J�^Iw��5���H���s�Buth�����ͻW�_�c~T�z�������	h+Mh�â�Z-�W�y��H�Ke��*�W��Dj���C�3q񋅓,5|�HB��[L�j�0?^�X���^c�J��hם|���P2�b��/k���e��[��s >����?G���x�OL$�����=C��1��3Iwzڼ�n���1�Gȁt�ȕ�8S��C*�љ�\/�׾����T�x�U���;�ؚ jX8��I��R��@��ІDo�#\�6���`��I���w>&�9|��N��p�X��ɥe�vR�&B��\�B�ϹnO܈M>�*��U#[�S|.f�*�L���JO:a�����pA"��
n�hߒ�Q��+�tsŕ���6+��a���1�I�X� ��̓�5Oar�V���r�Kb������ɐb�
%�c���4���1U�i.V�ݩ�� K�&F�tδG�����3Ս��1�͛�[P�����e�|�H*�9��W�O�~MA��\"��T��l����[K�O��`�O�&��^#$�X�Oۉ�Z拟=E��'��}'�i�p�21��:C�2�r�H&|+E�X#�, 0�������<���v>6*�����C�Ig��[�:鹍���6� ?vg���I�(W�5ʁ��X	�n�����J"�6[��*>�N�)������f(vJ	9mWQB�������?L��߈��V�w������+��FZڔ�BP�;�aF݋1�D�a$�x3�^��s�,�0��� 
�����Tv����	�v/l3�2��^I��yG�G�Xu�4Ƽp};W݊Pm��gg�D�v�M���i�;Y�$|����_n�Dv��8�g�h�<g��4�C�l�f���F=�W����)�ˌ�
��n�:�2�� ��hd�� P����YL�~,w�;~W��ƪ�#�ѱR���N�릤�#lR�E�,�.|����^
aYa�-U����|��G D�p�@ o|���F������Bg�0]��ް��t�.fP����E�$VS!M�A�(�_r"B�k�����#���I٭
�e�9�f����񌹃�izNS�� !�R8{=7{Tܶ4Յ~��>��Yc�у�9�;r�\h:h�2�G�H{�~�,��@���`T��P��9��w�����5/)��Ff::����*9���g���j`�`�M�'FJӗ��%b�b�'�y���)�|�������OW���m%��臣��,�Ӹ��ȼ�0Q��{࡛��k��1�¬B ��ר.c�ݿER~E!������@��`<�7�� &5���E�4��_炻�ݷR0��O�t�\HJ��~軵��*�=���W3����6����> 0�Z�_Rp�Q�',f���bm��3�H-d|A)�՝x�����k��
��D���:���V��C�֑�E��������?��D��ѣj�~&��*��S���-������ECw5���NO7��&����?m�����E|� x�(Q+o߭pq�o^<ă�x��������S�s�mq��%{�:+6ҾC*�!��5��b��dj�>�� ��t.���Utf�W�Y߂'�2�7p=��@����^`i=�Ubg&/q�K�5G�J�W홍�1�u� �lL�,Y�,U0��*�o{s�#�S����u���8�KM�����iW�^��P��q'1�̻�R��A�/C�s� �.���%m}Lk�a\���=�93�@�G�ޙ��<U�?��XxZ���Lb��0�R};P0%ԫ2i��uo�(?{p#�=!>�+[&O��-g��1��Q��/��+O���b磸H
���B�Z�v�G[�'=;m�k\>��ݍ�*�.q|��csg��� �4�o<��/G.��q�!D�}��$��G^�;�i�֍����*��ZDl�;�c�g�tN�TO��yȳ�v~�/���"Ek�	��&�����.~�	�L���
��ڵ�ڍ�Z;,�N*;L����jr��#!����y��ɜ���/E�ٟ��@8X��k�;>1|6D4=G�E�ѓ�PSR?��MLGD���Ρ.��Kx+s�Hx�5�r�qɌS_h�$�q��&���-��x":�繩�)��-� rɔ ����m&�x�|�I�C�]8�TA�Ģo�8U:��F=E����~.�S�>��=u����?�=��]!y���E�4����`�6��d"]���b\�ݦ�t�����s�l�����|�V��ǟՁ|A~���Aٔ�
Uf��@5<�G�i~S�����̻��4*�&�4[���H
)C��G-`ֆRe��M�5a�;�O_|���Yl�=[e�ce-l����sQ �ٻNM)���_z�8�ة�.5b�h3l���@~u͗X�� Gy�u��b��r2bdm�z����P^ʏ�<ἢ��-y�!6ټ�%åڗ7�.Pg�l�]�zҷ6k)t���m6@���_l��~�A�|"���W� ���8I������T��d�u��?�n�lS�F�}�US%��2b�)- ��D�o�{n�Y���F�Z��sW�
���i}��u���;Y�<���I�-����m���\��:�=q����h�~8����/���żo�`
j}���Z]������Z�,[pg������o�>y�,�z�oA�\I��R�n���s��>���ж�7R��IwꬡtJg���u*J�����Q�7Zݔ��������Z�)��{�MpC�h��\�&%p�W�q��8ޏ�>��x'"%��2�@i�x��4O�w����<0�������"S{o[��Mb~o��p�!�Ќ[��ף��67�$+e�O8��XdzH|�#	J�����4�I�9NDa�\5����@���>�W�"$�-�7�M�#��~�g�(��^H΅ʮHO�Q�j�X�Ò��B�t�ɿM*���4�<��ʕ�o��*��9��pi����]�o� \Ğ�oɤ��e��d�_B� �_㋱����(a�0 39Y�&![=��f�x��c��o ���������?J�pyt��Bs[P卲��Tr̥0��Q䪎B�ܛ�V9�\��ȐA�%���5�!�ݯz{��,E2��&��w�I�����n��D����H� �����8˯#a?$!������8��IX�|D�G���Q�mq�j�G4?���7�%Ir+,9nX2�~vVb/�3�?����H2�@
��/�J�L�w�$����7<�Mtb�7�_�u��&���y�۔ۧ��bѾy���4��H�N�]:{w�d����Tu�J*q�Z��v�B�⑐WP��(
P��Տ�ߴ��a!�uʔ��e-f�责Է�߇��=Rޝ~�*��X
��z��(�Hq�w�7��(�e�C%��E;�A���辋5���p��nv�௧�P�b v㻩�wX��=�z���nu�?XlH��=yZ��J�&E�o��O���e��E�.>�/*4	�Fz���b�(�W���%�U�#�u�!��@5�����)�ˑ!��Jk�<�?1���A�j6+Ŭ���e�:�#�ݓե���st�]���_Bk������b�6���TG�G�8b���������D��%�ZE�І������O�B/�h��Y㶇WDz��N�t>�z�1��QDܕU�+P�����0U7��=�=H |B�|ejo�[��s���0S+��D�����7*��Qv�Y�!4���p14�ݛ�����~�eJho����7j���J$�H�[w��X\I���-A���4G�Tۣ��e4Kʤ�Sp^
��	F����uv�J���Y���I��Ri��.q�� �'��T.��H=f�B~J$w8x�����n/3Oq�v͓6#!�;aU0�q����o�,��[��c��ިy�� )#��Y���N���+�ť�� ��<���9y=Px�Ա��XN����u������Ȩ؇E�S�$ǲ�zw���ue��}(�SN�&�=�\!4X��-;Q�ۅ\��WKD�O��(���"\�I������G�~�8鹸�ވwz�֢V�_ήHޚ�]�xv�ӗ�'{�{���М���͍�XS���K��\�Э�r]�\�Mܮ�Mq^�����
̆�xn\Ee����̊�H�:u�S]\e��\��ta`̳���8��T�����J0*>2p�})�f�
iHskrBY��+l�3R�����|�_1�V�����24[��'t)�SJ���;@Vd���E�&Z�R�M�M[���>�K�Z&����#Ю�d��ebS?�|�M;
ӅX�#�J�=K<3�J+�#��{~�#��B�r���,B� ��
Wy�W��d|ڝ�"����`J���t� >nE�,0��7�p7��f1�>u���h⍋3�����#&!��I�ʁLK��3�X��]ΫvL��ǅu]���z;�w`�o����*���T.w�;B�QG�������r4���V���SP��=�a%�!5�u@ɉ1�ǥ��0m�\�z(�#�J�v9��� ;�uy�[�>�5r���[�S�S������b�I��3w)3jaU������P�@f�U���'�-*R}���%�fA��b�{���~�9yl;�_w�}kb�d7GA[@v���I�$X�T�d�(]�2�M3!�r�W���T�/'�{B��{�G�I_J��0���́~Z.
������1�Z���(	wmLR��q��л��F\cSD�n�s�~����0���}r���߳IáV���Iq/nn�g�؞�$�;հ -��"6�$2�-�)��m� ��F�ys�gS �6^D��4t2��$ef�i��%�Y#�K�/]�D%P��9����' >������r��IK,���3Swrt�;4߾V�9AG�=*��C�7{�5Ҙ�78b�t�9^�r*��}3@�ih�֟����,κ��i��XF�uH�ΠN(n��Wm��ty�k�=;$�����Dcfu5��B:T��,�G�V?�s��u��tx8�I�s?BH�:�xIкT�,h�)A��A�0�wq��)�# "��>�W��W�?1��E~_����
h���eȮ�AԢ(ލ���>b��d�p��Z�k��3��1InBn��h��>�-��#?�/UY"��.��t�}׎{�6��g�;�1�4t��lV	�����P��C7�s`�#%�	��/��3�?j�&}��k�с�Ҝ�6�����*>L4-���$�:u��V��޻�.��.9�_�e�ָ���B��+ח6���h2hU��ԏ��`�B��i�~Qi��[�����K���ð�B
]j,�z-W
��"�'Vh�ʫ��o���+HFVU��I��uKk9l�l�nT�t$\��=`j�.:����Yx(�8���h�ٷ���?;֫?�Jy��w6����[�ɟ�������3r�<����q��Tf�C=@Iy��qqF�VƔs�g���8����*n�G���`�@*k`��q��D��l<���O��,�A� ��Tgv��5g(�uMzV�Y�ICG2Ri�
⚚��D���W\���f�t�n�[/̱�ЄŘd*x��N�3�x�$��I�Ί>|�.u�rc|����r�f�Z���/��X#&5�c�')�="A%$ު���CZ![��C�k���o=w������'c
=�5�e3�����8p��Wt�I�TY8����b�|W�H�!P��������tlD�!�A�Q�{,����wW٤�JK���%U�M��\�{h��]�'��qŤ�!��'�¡C,����#yr� s�e������$B�ړ���N�t����*Tv���%�i�m-�?��"<S�o��w���e!�΋�y�G&$j��q��Fo��M7�u�e���H�~Ֆ��f��y'(Œ���pG3Z���/q%�Es�y�]�3mc44jVJP��FV$ӊ�y��N}�r5������՝5���t� k^{�"W��:��S�,2C2��/����������R��3Mæ��'w�^��Ѿ(P���<,˻\)�}��C�DAw���擵�G�<���g� ��ũ� =��8�߻|'x�����wa@���
�8�P���ACMp�����͜B������8Cs	�l��t䕱C�Y�T�3O��a	��һ���)2�r	�{1�il+z������Y�҈$zD�m���jݕ���3��.w��������s�%X���I"l����ԊM���ܼ/�C�3m����T�.{d2�E�r"��ܞK=����my�&�&��Y���Z��Q��y�����i�\�z�2h4g<�= ��N��kE`|QX�	�pG�>�]�ЅN�O�=R���G�M`D�nx�m#�#�����0w�[���������>
K����A�ܕ�v󱩔�|JY�1;�覟��M,�U+��I�A��_��<�O�$0�nChs�A��Skwt�cJ���;�������0x��gV>�]贈�J���GQA��rY��T��g1]�>���4\su�5�����5�(����"
�T��DPj���}����M��6-󀚖�<�*O��n�L������E�e�b�4��<�/W���}�=gU2"Gt;�NW�Zv��ٰ�a���Ux~�Bz�x#��|���<������ѕTщo�-�a�4\�xC���!��/J�z<y�ޕ�������f+�|:�������H+��iشZ�D���)����lr|�����n�� �[J}�V�ә�R�T�����w�t�8f^�ʻ��I%^�C��Z��^����zs�36D�d���*_�z4�{]�0�0K��nD�0��<_������L�P���٩�>+B�F������3'+	��K�xa�0���V_!��#K�z�ھ2���RJ�;���uV���/h��n��=�!�%G	�gY[Q9����_-�kD1o��s�c�}|�q��w�RP��ܶ���J�q�a�ʵ��Yu,�^�b�_�d9��?��K)���cr���)=>�M6 ��ҋu�W8�@�O��u$j������	|�D�)j�#e?�K��a�t=����w�M <J;���ǲ���sU�=6ΰ����=��AF<B���f�l@S�^��]OgŔ|�������#L������$0���g��y�T�B�q���	7ƈ�tU���dw�$�<dXϘf�M����܈��c>�^��a�s���!b��o��5�v��99E��~�Esf/��8��@�M��fpK��*��]�ZϹ
n1��H�P��<� �Q��)G�e�P�t����H+&���<nX"�K�i�����.�Q�;1��l �qk�����4(`(�����Y�GC��U|4P��h�1���P��\�71r|�ωŧX�)�Z��,[{� /D.�M��Fs�w%��$����֚s�[�Co�0:��UjҲ��J��Ϭ ��k8�X�h�@�
�{��)3]z���'��ƍ���1XN?�m�|ۼ<����M�'e�k�|��i�a�NA��P5ro�H�b"V�6�H�@�_}�Jb���Wn�9�%����[s[�Z�פ���^��#�[�hB5>c�[�E��,:�Ħ����;!��A��V���\W<�CٕvD%/�%��	n۬i�o�4N�ߋ9�2��pʥϸ�i[d�j��7�����F��_�nUV����lK�6uvS���%(�Е�����qp�]7aP�~2Ճ�b__H~J��ԧdf���+�kz`9���Ԥ� �· 9���U��"��8О<�]��,�+GېT��T)���F�^�ꠅ�`l�d�ϵ?�e��?��#G� �کU�k0�u��eT�0Ml��56�y���W��ny�����`)�n(ۜ��V���u�G��HՑ�(DO˄c��O�=���&�T͓M�IV��/��4:���ŕA���Sٮf}��Q����d���ը+Y����$�������^�3�T?n�R\L�ө�⫬��lC�d�5]a [T5�>�{V�I5�	�Cߚ{�!Ϊ��W��畕t
毌Dqgc�O��'��X���;�Q�>�����1�WS�����h���*���.��"���d����'U��=�3����7E+#9?*��ΟR�>(_�i�O���#��k�E���A�ҝ ����p���x8=Y͢g�Z�6�k	������4}�~���x�{
��+�H b�#�������P��w����gEb6pΙ`������ȥ�C����/�]��r1�/l� rE}�p��(p���:*u��ˣǭ��)W]���▝�2�|7u���@8�ٮ� `��=��D9��h��L�,b�&P�F�ׅ�+��+������*��צA@2g��^��C fy�l���Nڌu��:{D�z%ۥb�$����Y�Kݜ����=�(W���J&�N0�g�>D-'�%i��D�*��&�A�*�1V0�ҹ�j�6P_�}��
.�? � s:�z�ˌsQ��n�$�����3��^�|NZ���uu�X����D.d��&ew���c<%��0���f�.�����M����R�jף��i��e�7g<KՀ;�q����_����N���EWd$���bb"�\6��ުY�E�,d�cו�毅Ñ��sl}���z��k1J����Gd�& ��N�}��}^� �w+ׅ.�BA��C�K�!����t����Z���<�eWC&O]
Ƚ9C��x�as Z�
�Oֈ��d{ٰ���h�8&BC�N	�=���boև�PQC{[ȡ{�I�g4�w�fnƂ˾��D��~n��vӻ��y[s�8��H�ғ�F.=,�#��$JKȚ�r�2��@k)�iϴ��%�<�_M��Ա���Z�ٞX�vS��]Ͼ�7� �����L�^��D�v�;��mV���Ͽfj�(�}ݵ�J�����T~����_��&�	��-;{-�cEx���V���#�y���b��SyS��iȮ�%�O���İ7����_��<sG��:I*=R؝��@=̭n�=�h�ǌKʿ�H �3y�8-��-��Z�[T�����������])?>�M��}��*c8�m�:�vʧ'u@R�z� ��Qzߖrz$�}c=>h��f$�"y����Q㹄|rs���>Ԉ1۪l"�+��ފO�6���٩�󽭍[#EФ��x8X�m2U���@U��*U��sJ��0~/}t!��ev@�1~H����	���
�л08��e����Y��o>C����,D���!����#�4�Y��P���o�78�0Z�pe.�&m���������)���<z� UJ�W,~�b��v�#� �8�
�?|��2���`9�-��������H��x��O������R��{���o\)@ޥ�QyG[̀[>E�-�{�L��na9�����W��;X+^�Rih'�U:�Y��Y�ة�W�-`��<���A����+Zlӗl��B:�6����7;V��N�[�([]�]�8[���Q������2҈��W��%��M�O�U䠢������'_�n5'l�`�#X��h�Z����'��9`߸�e9����m����
�xʩ�����E�\fc,A�޺����.Qs�C������nf���r�q�p�a�*��I��/�3���hA���S_$/���^�vT(��m�u�/��L�/���F��AMW-p���Mu��ۙ i�Y����ǬH����v���Ihr#��������4NzHԛw< �4�W�Q�o������*0"C�L껼EC�M�Zcr�����H�/7�v�]�6����@�3]��5q�7��I	Л\zu� ����HMt�&ݦ���`q����	,���D��(�gڇ_��=@��ZL}	!�P������yZI��{�����p'�'��dC�N6)c�C��~�9k)��A�^�_��p~}tfqk��52�h�A���GVR�,s]����	�]N��k%Y`��K�q�����J�T���?,Md�|�^d�+|�#���X�7_�}(\�'�j�HLk�e�+�=������+6�/�௚��p���*��vu���]�#;Oe���a~�ǽKRP�t��Y�1b�e�2)�|3As�5^�Ga������'��V(�ߪ��1���B7�W$�@N1��q5
w�˗I�;p)�!Xf�=ۅa!l�b�r�٫(�(~�F릹����"�ޑ�i��������7�n�&]/��5��q3�5���<�K�#G-0��L��5�SV����ɛ��fƉk䱭�2��'U���͢n7������1�!@<ؤ���*�����e���[���ީ�0-bb���t�1��>/��Oz_Y@~��6�nP��G�i؎B�d��g�7|�Wv�L��6j��ϨB�m:�&���(e��<�=[f�gc)��)3= ~����y�P�=A�Y��"�w���na��r��*�7��a
T�"�쭌�y�����aI�=b��k/�v��#α�eL�M��"�8�>G&>�!�L㵬�eG�[���pRJ�0(*F��c <�J7��N�\�PŠ2�c_����ٚ��¨��}�EI ��I����˃��(�v�l�B����tٳv��ԫ�b�Q��Dx�l�)y�xE�P�y�G���kZ w�_9���C+)���P�J5�A��*�n�Q$�w�����{��MJ:��L�y��fm��������q�������k�2�
�Ӕ��n��3��[�ýx�� q��K�qcA�D��<!��	+�T~�h�����G��青Fs���]l~P�:���~ ?	uf"Ӎ��%�/b7UZK�M��pӂ�|�`E����O����Z�H��&r<<ΘLjAږ���L5��j�<@:����t������  }�OI���*���Jd܂�qa�K���%���f"\8r�'��>+dlc��o���/�֪2��9��1t�܄+ b�,ƛ��JZf<Ӻ	�V��Z�G(w< �d��&�q�a�������c��ޡ��L�g��@������X�uAB�Y|��z�Ɣ�.=�D��"�����6S_L���ڲV�����w"���e��/�R+��L��_�0|kidA^uv� �L��T%g#���D�B��Ə�����_t�2ڗ#5�~:�e-Ge��C�hr��Pn����WcG��]F�����^,��3�n�m?Me7Z���@C$y
)�G	��;)�b�W�`�a��!���-!6;鈆a��x�4.@�)?�sZ�����Z�T&�� t��H���'���a�^����J/�oͻ��1�=s���:���s7J4��]�����C�L�FAXQe��Yyҙ��F�Z`�� ���៶W������s♽���ْ�����RA �E�EҠ}�vז*�������@���0�G�ȋ����vk�g	���q2l���/_]�_���͙ ���!u�Am*G��.�R��v��_]����E}�D��x�]W=|�E�,HRpC
3b�r,��uC�nj�]����\Tc�ɗ9�>5���h���2�0rPC�}�-*�5�Jam�/~(����Q=*Z��%��w�?�Zwn7L����޷�Av��d�Y���z����AY���"����0nŗd��|�#<���UO���g�\c����(���"��5W�x�Q�xnS�,G�Ksd8Q��Ib����l�8=�f���2��j�A�|�ph2��N/#i��q��R�^šG����ތ(���j�H�3�0	��-㑯��"mT_��䄐��7#���Nq��u��m/z��n]ˉDb��h��'�=�E�Mk���sy'�eJ���iP�>��;ȵ��~���P�M8E���AL��ub��ώ[O�m6�F�����S�ѢTԫ	�W��H�BR�k�D�d̘�;�G��:��f�n�f�hJ��=r����x�5���TB]���\YW>!v���_[3���� ,v�F"˦CKC[`���z&�(+#��D�J�[�:�3Լ,.�����FIr����2���+��|'�0�j�ћ�c��NI���[�����Hg���e���N��)�:|S�EC�mhJ�,zzb�?]�����W����=����a8#�1sn�)���W�b���hw
�{�Ϟ沰�;�1��'� 9�������$!G�Ҋ�R����,�[ꀴs���J��j���A�����q.Bٙ�j\n>̤R��� �����T�~1�t����\>@Sk�W�<��p*�/��Y�������Z��\��<!Ӏ)����~�hoĬ�%�bwg�B���}ƻx���슑�'@Vsj�x�̈́ �ʏu^8�2x=0D�6��K�c�0p�7�PH�r�c�>�nK�_�"2t�S�vy_-�E}RMc�L���<�/ڐ�v�Hj��uug.�;�����_��&?��I2��P����]��ƛJ-��� �
cxT����OB���-P�rn�i�!����_�Q�,�&XWU��a==@M���ߐh��2��
c� ��W���P��	�{k ���1c��fT�b�ڄi�����������g�Ǡ�)3����#�0sj�����{���Z0vD�W��-���&���:E}u�_�r��� ��ѫ@��-�����<���=rV������N����drS
�����^�apO�vv�+^��$=���6�kVѢ2x�K�ڋ2�^{����)���ܫ�2�!�w�}Bl�fb>��[���9rP9���ɦ�p��A1İ����ט6A�,�D~���M�ޣ�ԙ[m�_�	S�"�ݲp3T�n��J�q��c�h����;���]�"ʆ�P��C����>�o�}+��0�[�I*{�9��x��jHe��u��q���~ls�E��JR��F�
���F��_z�2�V0,xD�����<a�
���rF�U���-7f�J�iF�!f_�H�k3�HX��k���`����r��k���B���4Z�W/c�V�#�w�Y�e5��v��fl�;n\����Ә�6p�.�����PJm��f#@����^V���tU>j,y g�(�)��um�;�� lc�?���;X4���<�ұa�55��u�Tn��a{��� ��n��)6-�-mؕ/�<
���SRo�Or��n��y`�!g�Y�Y�3�q�>��gG\2�Ĺ�s�n��sc�I*(�&�
��Q$_�Yf�޽ǎ�l�W?�P|�3�@ĕ6�޲ѭ�u$�Bۖ�_���n�@�t5/b~
�׾��aX�Nn��;��� �&e)A��i%O4�a�p�er�ܮ}ή�*�|:<�;��e�g)*P-}��b��BA"+���i���G9R}��K�2��U���"�%n�8�T���C؞p+�1����������O�+~	X|jXxg�,\�q�*��+B��-o;&�O�� ؅��ʬF���Ax�꼞�S\�<�l��o��o��QqG;�õLa��E��e���K��nU�߳'��z�>�5�Y�*�,�V��EF��V�f�y]j6Ѣ�ȸsG��A<��q�ƅ����tV8�2"�s��k��w^��6�ug������ƺa�7�D��fr��	PV�f-��^�� 
�f㿣ĐOR��Ry�W��7����IsN��6�R�Q�y�{Ӂpc��3��ƽ�s�g��k�<�\���C���'MA�.�a �Nx4rm �rݵb��uԮ��uGh[�Ϯ����suԎ#'�S�W��D���m�Hag]o�����-g��b��pv -�s\��d��ƪ-[A���+'�5���5����/����X1Ѣ�)��7:� ʆn�� �-����xQ[3x���^�J��<>z�W7������ԮkK�i�r"�v�gt������.�*�b��YH����au��G�_=�X?�}f�'�8���7#�)y9�K�^��X"�_m/��I�dŀZ�Ͼ��v���}Z�&@�Ơ��������w�)M�%:�-��Β����y��B�>)UB�I.Љ���.ܔZ-���@zB�0n)��U��q��+��'V��G�0б���]�&�d|[>2���Xř.c	�&:v]ȓS��	�����3_�X�mr	"��Q�|���o�#��ܷ~�����LnZg�����ʉq�r�a��Հ������/���E�P�U�ɱ��:Ad|jG�a*���j�u]���c�`���Z�8���ݬR�%�sf���g�to���+|��Zk��ˊ=���`Pꬶ�G-��!�)��o�h�Zm�ϵ冗���R�ܲ�c�S��|y�gW�5x�k��o�奾��2�KV��]cg,COw�`��&?NI`7N��\��>v�����N�P M2�;<��f6=⛃Tx�)7�2OJ�(@�����A�qmj�9Pv�s��/���TL4�!�Hi� D�n��ۘ�/���'���i���<�������ؘ%���D#D�Ω�t��?�a����h� � ,���l)�Ozg��
$(�iH��G�U�h�>�G�HΞ�=����|t�W�bDB0/RN$�6O10�:���x=5��m}��L��������NE���*@���4GR�t��)���=1�@��P)t�����=,�ޤ�;ѱ #�rK�|V�a�$�>�r���l1���=�Z
�zW�����CiO���fd�t���G����74�Ϗ�iyu�qo��^��	����$~U��h|�D-�Y|�))�^Mn��`4$����X�dL��$l��P�b^Ų	����],�H@�υ;#�I�N‴������d��,���ɼ��E$Jݕ?� �s�(�e�)�=	���8���/̗2��Lʫ��Z�Q?�v}�ST8f�f��<0�I�򗴶fE�u	ƙ�X�f�i�{,DB��S�!%}{c"uZR���/�=�O*b�4A��Z��9�۔���0��T�2���q]&1a���N'�K21�6��Ysr3�o�S4��Fb�Zl+�\�������˰���UM��s��J�l`r�j�Oُ��*�8��զ묒���L5�/�U�t�?*d��XL$����%���c)�c�_z�'�y�����ϸ�J����֪o��r�-�2+C^L_�����縧�k4��>�?���v�wm>ՠ��?@0�������6�w�P*����ʼ9��'$��ړ��9���?�Y��=o)�LL҆�����R�!�z��̪X���3�~L�W,���C�E��}\r��\ 	n�&=�4�>�4��� ��Hp���C�l&��pm�}�k��Fx]E���v��:
}�`4�.P�x),#�����˵*�W�i���A�i�{Y�9l�V_$�£"�Mh;!1[�P[��r�x᪱,:�j�\i� D�/��&��y�N�&��G�tJ��T�!3Rv�y�^��u/��)�<p���.���1U�@ͥd��"��M�@������C�G"w�j�2�2ʴXt�j���l9-֪���H.'\��jF�-�p�;˲�Ǒ����_s.p�2l>�>���#&���@%�Ǳȓ"�E�{*)�����RN�&	
:1L�������:��!v�W����6|0<���PĠ�І��r�3�� ��	q��@�Aڊ�+U�]]r���y;]�Ex�� e���/P�Z���	����5HF�I����#��+!=��ʲ��p%G�b�(m�Ƽ����v���ª"�R��ˀ}�
/�v�A�3��ν?���f܈Y��ӽ�Q�����	���*)؏GO�܄�M]�����[�P���,�0�}��x�d��<����"p�D��������ţgP�~�%�F��J��Z_�J�3�ɣ4X����f{�+c*l5y*��}V�UY�������"�Nl��GӜ�I��񄦸��}�g�&�v��o�1))�aA����o�u�o�1�������L�}.H��# ]��h���UYq�ݢ�h��3�)�.u<2��JG��3k�����:p^~�����&�Bo"�`�T��j[�̄5QF�F�!g��7HUr���^8�;j*	u����_����\	�:�*��L��R�q�pst�:��*���(����.M���0��Q��q@w?�c�o`���1��d��&ϓ��<q�ryvL��9mil|#� ����ph���H�C���X�<�ё�4����س[^�h�j��c�w���j��^��:*��WE�!�l0 s����`̵����+�]~	��!���N�P����0Ԡe+���B��'kFO ��!��}�o�f�t��A-(~B�j�\0cǅfD7�p����XKѱ�b&�y?_��m.��<XG|���.WSغ��;";���|q,\�N���8�ouh�2�$�X�I�Pv6M��eH�0�G �/�]T-��YS�hr���Q�q�R�@Qi�������q�	�z�z��G�o]C.��ߜ�����P��#=���:�R���3S�!��=}��8�G��J^D�fR"L�f��*� �}֠I|AV�=���_q�`��J��#N>33hґ�-.ɧ��ˉ�Ω����< ����Oo��ȋǏʙw�7g�.�N��m-��H�g���z���Jb�Y�6����w4��!��ڻW����D׀�UW�Q��Lh��"� 8�/Mȴ2�BqyQ�1��L�:-��Ki���|�������C%& m���M=Xz߫����8�]n�S���v,�h_���%t�%Y�}��l$n�̀��gQ��zv�-��3���p
�#�ﰜ���rxr��Tvs�wQ+��r.O2����Z�UX%iPi
�d.5] D�3������;�ė����&N�y����J�:���z�LR��w.�执�#�r��/x��b��H3�q�������P�U��[�W�&��v�ˣu���s�=$�y�2�,u��������@Iub�XO����?6ĭ��c��P�(S��jk��^8W5���$��)z����r�JL%4�al7M�������&`�,���d����V�Tp������SɼLfW��S#�!(�`]V�\��n�٠p�^��o��O�z� �?��D?�9���'}4��M���
�G����R9]��`��u�1ǽ�꾦ȏ�ߜ4�o
H�,�w��Sh����o�Дsx)l%�����>V�Y.��ŅR�8�.}+����ӚL�� k��K�V��ĳ�(�Ζ0�o��c�$�1��W9_U-t�^^�0�0=��kj��6���#�<Ç2��p�6ei���7�eo���?�g��,�V�ژq��7m�t@�ʲP+.���kurL�G��R�P�u��t���Q5�[/�NތO%�����O{��� �7"�k�a��W�n3P����n7�uf҈��Ju��r�'Љ�#YT�w�5h��ܛu6�#���S��cf��%���c��у�(�}8@��z��ƺ���ؐv(b��mE�����Hh�$R��A+�a�V��(%�mq�_�D$���Ց����G��\��Ԕ|���Y��#\P*c�:���j!"��f�G }+{�z	�������(��J�X�/h��^�c9?�/b��2$���\=d�����%Pgl,"����^����UQ���G�P�΄��6�'����Ȟ:�E����͒zF[ͅ��L��zm�T�H>ӤVC���	�%�R9y%��'�9F��Ez���5��P>Ƿv��2u'���'ۏ�~��4y�����+-&p���9@�w��f�STX��N�X"�M�%tC�'p�?
zN�� k1��'��S���g��4\��u�R\n�Ģ��q=S���h��94�0��6e�=e$GdW;ն���ɇ�U �[Ձt����r��X��;/����<g���m��h.)��{�ʩD�r?���>2Z��:�G��P�
�U���x�hz[?J&��/�J}Ԫ�ýFm�1�8�-��S���N�|��Q}�=H�#�I6�p�ܲ����\�1�f���в$�MteV(HX�_k�(�%�*���/Zi�'S:L	�6c8�_Us�T�ݩ��O�W"yy��U_�r����h'�����)�S���V���4���3�����l�l��7�7CWB���#>�aD�"5fJ��7h�_bgh��P����>��������u):QZ���,'���=�(��4�,"n�-g�= ����er� r�x�.�o]�/�m�� m��A��R�,��Q":��ޅ?0��O�j���v��p�Sw��c�����c��1�Ih ��k�a�Vؽ3��pdGiI���QT&�P�+v�g���*ľ2ެ�7��Og��u���H��E<���]CO򵖇GL=zq�V�z��v�[|����E�M�0R[�� �{�����	;���k#$��xhTra �L�Xjv .!�(x\�*��7��๸*:���!�*�lv����H}n1���Lef���1lQ|%GP6��5�簘�Bxޕ�	�'�B_�n3@o*HK=����p`a�0�5�щ���t�^7����Z���xu	_Dcu��v�)Pz����zH.T:|�$?�kQ<���y�#|mj����'���l�A�:�y�Ц�W��n��Zv�r�㸍�Ƹ���)��|R���j+��vY4��;1c���#���a���6�7�N�8N����Ξ$���`W��$#��N�`��	��ï��"�dV/w�{c	5�2�,���s��u�!�A��$�ya�Ƈ �t�{�H���)��9�O����Z�n{O��������oh�&����b����i6z#����^���y>X���Q�m�q�_�.˗�8 ���Q�va���eǬ��
����S����Y�Y������cF�]+U�T왭ٙw��x�	j��o�r���H��c�V�\"��F�j.ػ�m�*�������՟)��˲��BC�T��M�{T��ϓ)іY(1\�:�Z�>�s�M��r'�0�l�wҮ���i0�K�y[�@zQ-�B�5z0@�&�������D�
�eI��RS�8�f�U\' �1����4yd��>�O�ԉ�b[�͡C'������C�ԗ,�.�R �3 ����Ji?��w�u;t��I{��W�P2�Q�Iv��wf��wBU�Fg�*-���2��F��m9)����\R�`*g��7�x���Z�n��toP�LV�j��1V��Hx���r��Y���,���*.���֋��X�����b�Ǘo<Q��mVUT�m"�]r��\q����z��ּ�s&J� ��	�Sw4^5�\�L��ﯡֿ6��>˃ڛ��Ϳ�T��q݀3oN��$��b��ѥ���`�}Clc6&Ƽ���ʌ2��M�;�c�I��DQ�:��F�����!Mp��)Hi3@i�����𐄶�����[y�+�ݢb���4��]��z�Ҹ�$�9
:p~Cb%��P*�h> V&���i|�Yv����Q_QSpJ�n����3;Ɂ��=fc���tK-}�����.gI��hU�v2�}�t� rQ_�tSvC.��3���2w����ܧ-�??��@��Zd���ޜgY�̠�f�+^~ �A�l��T�������h'�'�O�$�0�OV�����h] ��3A���h&��6��<Wk�*9�p���H<n8��, ���/��.-�����o�Ҍi����	��{��\�B��
�^��C�X̝��J.�����Joɖ��k9�wD��<�
e\"7�9�n(U��U��Q޾�hl�Pآ{�Q��u<��T`u���]�y�-�/�y��� �!�Y�(��H�z+�k-���v��3�4544z�95���Sm0��C6Pu�'�2���B�2���\~)�>껳��ݘ+JvIq.[oޢ0P��v\\:�����qt�Sd�㭽����`+��e|���4�X5 ��J�E��ֽ��T��vG��W8�'�>$�[L�)�9�M!v�I�_\)�-qZ�w2����IW�@��?�����!�Wp�!�ő7<r���f����ck�x��Kfq�JU�dX�ġE<�.���O��0��d�xt0&3�E�@�P��~�&�P���cʜz��5�$�f'N�7~�Mm���#`nCׁ��쿉#g�:|F��\*9����=k/K�g�"��4#�W��JbԻ���=ﭺ��u�g�x���"�	��e.%�Zv�.0�U�'�\�Z1�vG�M�rh5�4,g�L�`+}��p�-��7����5dQ�5qʥd�O#`1l^9Fi���EɨX8�5/2^>s^�(�m�G����Yzecb	<U1��!h��5�[[���mX�2��BEc/k���k�Ь/�a��������f�I#���؊�"{�sr2gk�K4����)Bu|��gg=��rϷ�%���$�����@�$�z��rll	/t�@_f���}l[`!�dS3���S�;��9dJD��Nvu�ۊ��O�$��~�i}�Ɯ��a���x7Stk�.�inMA�l��Ȯ*��+�-\�">I�v"��~E��D�����"&�AI5�ڱ�1�+E��s8���HT��gX9и��1��~��WC<�q��[l��f�Su�RK����[�%j��t���E�ڞS�`�r�f�Ȣdq��w.���ڋ�5�S��Y�~
�A~��4t.�Ԑd�� �e�+�=���G_`���ҍ&���|j�Y���O\6�tv� ���
���cV9Ztڶ�o�Nej�o��ilST��O�� ��Q+B���.QH��'����黚����W^� �����$[<|L
��J�[��=q�3I��@�9����ln~?|{V7�c�X���K7��?�N|�/]��X���
(]�x��\_��Ü`a�0�[U�+���P���S 0�H�j�K���=�n����m�kU���,*X���Ą��;sk3*aއq�����b�%�N@��m�F����5�X12�:��,1'o���CTbWC���=�d� w�i��V|̋�H��K��rS�:z/���f�Og�pO����\�5F���5�D�H*�<�$�v�#��뙖Pʺ�/�����x1nQ<�*C�e����P��(�'��\�H�7��eJO���p����A��p��ɤ�+9�nf�g}��ql&&�ErX����J�&��.�rMg���i�+��S�m�d�D+�ұ[�|รfT�9�S���ϟa�
�9\co�z����zv;Í�hD�j+�],ew�]�MG~B�t8!EzAb>9f��q���k��������e�/��tx����1J'�}��A?w��2j��ן,*�����NI��j(�?�N/��?CAq�]@ )�����i�/&�d�`W�T�x�/M��]չC�I���ӭ£jѸ��0yT(-�ޝ�R�ŨT���N ��ɞ���smt�H��6�.�lm{.�C��R�B�Z��͝�-)L.�x��a���w9�-��.��a@�K�B��1�n�W.��?!C/���1���c��ZxA��25��aI�W�x��QD&�_���ɓ��H ^y�N�:��Y���i���/TM��xɵ�X����>�/PL�z�4�P�o)Ҝ10�K���@$���P`�~����������2�\�ق�#��FD��1��c�W2�o�q'����䧬�B�h<�.��{�����@%;�C�u\��o�[�@�D��bzKA�a��ڍ)[�k6��_}�wVR�V����i�"��q��Nb �n�\�%��"�#�Wlkޱ�~t9O���78=1^��}��1v!x���l{���3�a�#d����bI���ձw�!�Z�P��?A�q>���	=i����喔CU��e�M<!^�Ќ�26�B�CRk�p+�'�Wg�Z��;�gR�.)�*�F�����a��QT�g�wU��,�$�A7ҏ��]�H��\N�����`�#�sⷖ2��@�ě����B��|�+J4��I���Ϟ���|d��;�5Zc�<��ǲ�����H|Z�S,sJ9�s�J�Z��q��IP��yk��r����|_zgx2wO�8����hut��QN�Z=m}P���r�FUr���|��r�Ќ7�-r���5�C"�R� �u��2�|x2�d%�G�Q_�5(��� ��ܘ���l���w�׳U���/��	"�m�0˧{ː[6t���7�X��q��v�y�~z��I����`z)�������/۞�)94>��e��1�)�"�X#���n��sMw�����m$,�k�٢ �$�8�x�0�\!����Fgx��?���K�������]����@<3#�`T�֊���fvJ�����n7p&g���۰_�X8%@ލg�:�v{t�۩�Ǵ����2{#WgHП�����6���[�4@�59�9�=6�oX+�4X�9L�Z���z�Y<��:У�l*������f|:�*S�1���v���c�8�Ԅ*GPPn�9ū9X����V�� ��xc����pg��v[�_i+[��
����oV*�(J����*+���n#�+��p�5�l��k*�P�޺�4R�?�vv�bD�yr��NO!���>��:�\����t4�d��7ϩx���%��O���a�SsVc;���
���~�I��I �C3�9iDm��$����>� gn5�"~��+����g �dU�ΥgĄ O8��6fgF��q���-^mK�k-?�������lX�XT�G�Ż�B*��Ҳ�9@ �z.8�l�#UC��v�q�,�s��kV�9O7Fj���
j$x��M��I�{@m\C_�/�P7�������~��-#��eG9�`�~�v,�^S
J����p`(�o��S 9
\��>�K24/5��3�8�T:.����&ֵY��h�z��)�wĺ,��
�3�kשL�÷�#�㮪�n�p�5��3=�����4*6��L�E���D�Cx� ��v/ {MB��A��,U�EV�d��(2��&���7ORe�Sb?�oy,hر���YM�̢���ߏދN� S��mq�6mn0Fpx\�P>��1S��A��G��{*՛LBT�\�=�^�դ1�nl>�,���
K�1�s�Ù��� �?�%B@��J�0���������fz�t���~�o2����|�����v�UW_�rL�N�� ���n47q��g���U����=�q�:��͡ x\�8Nk���?\������: ��VtrQu�
?��`�m��a�bO���0�ǲ������@�������^�V<�++�t-t�բ��w�H[�1�{{I؊�.��׏,���{T���3m��c)�nC����IN����� �Y�a!E�[��B������4���4?=o�.�8�|��T����*���w�m��
?X�44�F���(�6K���#�'�lv�� |�d']e�E�fR�����q�5bae(G�j��F�TT��"�GR��m-@�S�����'H7J����&�	���ӋFR��!(X�췿-U^H�9$^)�!A�"��TG�.��������t�yi,W��H�)��p���[�L��!\3�4VWG�6I<&���O��@��U[����hA�́���2}��1�kn��Eæ���C:�Z�y�Z��Fb~yt9���B %O�>��H���0r3P2�*�U[�C|D�4��2���P�qe��/���ew�F+��
��8��ꢛ�@>F��q�H�����[�[v��}�)���8j|c���?G�8N�
�:�__���D�9EI�����?��lR��2J֋T�;wn�2?+2��(8}������<ZO����8�	���b_��Trpzc�Z?����2=���8++�
�6�û��ׅbO/4� t~� �2O����rHZ{OA_����u���o��	�h�bf���%����/�|��G�2����_'a���F��Ā��5�IKH8߼*�/�l�� ۍ�M�6��iOY�xʓ�:��������â����z-T��2�e�/z\4Y��}�Yr�`S9%�S�v\Vb��ݾ#���nY1$pl�k����@��y]{�wi��H��U�Xq���A�&��L�íf��51]vo��*���2���SlIf�,6z���	@��J�/(��A�d���q0����i0��;�>P�t�_����1J{��O�E=����������6�|ꔤ�cU�Λ�l �ܟ�O�	� #������Q�,���o"��"��`F3S�6��Y����Č,���B���@��P��J3��_zy�n��Y�K 0�)#&�Չ����8��<+�žM~b4�#��*�u�I���uQ&�Oiᵉ��I�/z���B�z]����n�T�? \�cG�e������Ɩ�N*gKk!��+��
�q8�E�Q=R,��A��*Ƒ�w��Y(_���o��Z������M,Eg� ͅY������<�jW�b��	��3*�C��d˚W����J��T�1������s	� �m�0M����I���'LPc�0*V�޸O��ei/�lN�7�Lj��yL��0tNs,Z�G�  �%p��Na۱	AON�Ӹ&�q+� �iBt��;˝�`���H7�:]�h ���T�,�P�d���zd|Cr�F���=k&ok���$�k�үP���B�{�&Ѡ��}��[٘�|飯���fX)'sa q�2��
a)��������G���2�tja��J�٫}~c��X���F�gaDs�|˧́%��4t�=tLk=�b^�StM����iI���4��"�?��,z�Q�=	Of�o���q�h&@6Z�iġ�����~O	�}�/��R���Z���`P~�L�ҭ�#$�1�\v���skH�
n>�1��48/���E��~�j.����&a�v��{H�\��;��vL���\,�X�[��{Gb��H��ъaM�� ��%����Wy���#2-��X�?�^�	(B4�@�@�7�4��׶��H�V �+¥��;8uc�v#�<:؀�[y�� �)�<��C��I�$q�g_��tM���`HM��G�v]�S�K�o�����:r{�� ����BW����&5?�4�3����7Ero�����H3 \ɺ
@�$�j�X⢐h��
�O�D�/�Ӹ�dS=�b~�utҮ0�=�O�{e�`f���8��TID�H4����x3��]F�k�Irȷ�VeMG���qE���}��o��
�o��)����b"Jpw���)��N�E��l3j}D�,�5nl�/[��XΛ�VDlpo�p,B����4� P���q�����[����ߎF�߳8nF[��l0�d�~��@�������T�`�e�, �!�#t
S���܅ �<Wۆ/��|0��
FFC�v[�h,��-"�����r�Jd�+�}����q�Cր�C��l	��H��!����Ts�X���Wֵʋ���u����y57֖�n�*�h�΍�z��N���r���=l��C�s�G��Y���%�̰k樹GF�������/F �Q&0�5U���Y�T�ʚ�v�?�w}��Yy�/＠�v6�ҍ�)$��e�D!��K\�9X-4�ս�
�M`O�#�b�ǹ�z�ԓ��k���^��z�r�\�Nꞟ���/EdRy�oq���}���[ؑ�SHg�Sr{%Bv��0/&Ԏ�7	�g*�\��������g��(T�@Ќ0"t���,�[�V�7)K��,��q5�@	������܄��1���ٮ;u���۞�Wم���_bZ�Վ�F(��m,����iՉ��G�A��;
�(s}��=h�~�8���e�?�ѧ�`r�硤yé�$�F:i"���'�F�s������BK��Qw��a�4���)�Q�"k��;}-��߷�/I��\b��j���"X�M�7<���E��R��/��**���E��3��%�6\Uz8m]�I��^��ļ7�t�Cp���[$�p�i�H䙌Qyᐭ��
��/%�{0���	��	����������ѳk�*�-C��7֣scM��(l���'������g�sCa�AP�^���B�-�$�|��,� W2z��ڷ��	�z�.��*��M �-A��9��ƈ�`���_
d���88�����rf˔=��?���0�#�����nLӣ�|�<N@��3'�8'Nai���\e�o�+��$;\���.��cr	����#T;��v�<-M)D�Gj�{�^�
\\+���m�Us׆�b�ۇE�\��4ȝ�I��R�w��k����;���W�^nT��wˋ�L�%G����t�OLl��N���9'��i��ZۊӪ��(	��c+�ے��۪D	O9-)�i���b�W����uRq�����av��V��&�e�R����u�,�j�I$;M�Ox'�uHhm}�O�ʯ��Z�\�w!�~3wh~�^ f�&��A��@"�έ����-,�.��*{��g�V�X�`Π��~2O�~���.��o�8�<d[ݿP\�����t5��d��O����Ƽ���S`a�`x�h9O_=��e��G:a4���'�Zw&���)�ݡ-kuߩ����Ӈ�ޕu\��z	��W�y����K��_�eH�B�{���FŻ�/�ƌ�y�M����w���"X��4qZ�j���	d9�8d�X��Eu�z:"j�K���Q����sJ�L]���A���[�Ɛ#ً����-*�D�)�Z@���(}��넧�|ql�뼶�?�w�z|a�g�F��{� ��j. �ضʐoUj� 9M�_�d�b[�ƫ��u�l���j�h�o\-��!�SA����O�&��{�'7i���ή��1#l���D+�lB�,������|[�h!�Žy	[�h"��%���y�{D��>�����8ؚ�?�g�Ԗ���M�*GSh>�Q,}#1�v��	w���'2�U�^���.;0�Yhp�1#j5�o��Ze�U�AO��H��4)���\ψ��N�B�]�O��9L�-��%Ȓ�9\#�k��y�Ǜ�~!��:Sa��6���m�q�l�Ún³��H����$��ۨ���C��J���[�� ×���~ѥ��t ��sF��Ϟ<�K������j��aUU��Iλ.��Eى�H�X��G�v!��VI��C��4>���20w[��F�m���ݖ^����K��Npރ��>�/��MxQ���ѩ/Do<�M`{oG�Z3U����C�|vTu�����l�ɥc.�N�9�U��u{�Cb$�L�mz TWf�+�֗޶���	�/sR�<8�������F�UȲrJ\�k6k'q�~��qhIQX_A�k<�*��[�e��v!�&54pq�]4ȅѦA 	�H��Z1��g=X�1����ep96�������c�1E�l�N]ݞ?)�����պ}O��� �����#�����Xp�@�{0�T8�")����Yߠյ1=0��O�~��Oe��S!��l�ei�⫦�j��w�_-��{=/�fU,�xn3�u�'Щ�g.`��\a�
�m.E̠���L;�a���!��X�-�Oj���Ԇ�ED_ci/V��	A� � �U,�]WE�5��i�D��?N���/4ڏLW����@n����Ed��������PHE���c�����grT'~:��.�����o��_o�[ā�`����O��ڄ�/�
���� ��c�{�d7Vi���k�B��2x඀�um��[F���̐�ۤ��εꌯ��8���Ҍ��K��G���Vs}KX�n�Kou�~�5�b���y&wm#ɉ$V��]x�umՊG�$����� ʩ ������{R Y}�r��dhRU����^�s'�T�ph���y�:L��:.������s������%�����/�|p�f[�������D����1�kX*��?��Wu���n��E��0�!%,Ψ#)��K`^���rMѱk��������
�!�@Hi�#�s�/����.p@�ǣ�ʃ#@�G��`��A�O�p�zR��rfZ���6W�5f �GX�y�G�)�R`�)Id�����7�2Ѩ=��	�i�8��a�r�|a��TSU�D��,ldz��˚-�I���IF�F��ƛ+/=8;u�`�Л���Q{B�Z�H �.���t��g�BL��˻s��.f(
CZԭD;Vo��_\|�n�8X����>R>'1���G��Z3웍k�6i�K�<_5��ڟ��X�����
t�=���װ�Z��a#�v�=f6c�F` ��k���?G��t���j���}L��	J�i�B�@dRf S����O�fl�;��M�Q��SC'��םt1
S����7�hN'b��%�pρ�י�*���A���g(����+mh�|�T���*q�%��!����H-���mV �p�=w�d��4|3��r���u~��&^�*�C��42� aZ]���q�v����,Kk�n|��F��r�A^�>tQ�k�0)�="�nR�����E���i��s+�H DB�j�G��
�2CKKK��gSj��W�}�)��x}�A,��4z<�G�?�T��=��x�`vU��ĐJB��;{��U(_W�i$�Z@˶�G���^��:L�\�.lף<��U�#�*� ��qt��n�w�y�yfwEg�t容�ĉ����t�l��3�UqA9�qM����$�ov�BB���`>EnM5�l�CQ����{-ifE��5����=�r�V�nS):.�&p��/jZPw�kX�����l�zu��� �t���ؕ�Z�ou��4E�-�&�/5�j��up������>ל�LE�&�яvؑk�P��W����=-a�\�̠��t��W����}
[�b�e���Z�|�|��� ���c';�j'v��d����|z�|S���j�u���J�Ҳ��r�.�𐽙�h��I{OǾ�k=��}��u��FLž�׹�n��ſ �&�Y�������A^��Z��j-�-��(nϦ���rg�Petv+�/��i�Ej��s�lY�]��`�εAf[tp{�n�mĊt���!���&�E!��a`��H ̭� `���f8�5��$��2'^ro�����iڈ͑E�2�O�Q ����b�{��ka�43@gzޠ�s��4G4��?i0-�a33�D�!��:����X�.mm�amˑ���,t�wu��b�!��߯(�+B��@�SD������4_��|�p3:����&L�Tgo��"	�l���K��d�R�M�^A��̣[�o��9������C�B����ޚ�颻O���e����>�d�(T�
�=�څ�}e��H<4d�#󉬕7��c��.�Y��2��������<U�[�q�&���:��c���Xo},�HB�JQ��[��4�Z�:1�@@TYVx;�^�2(���1̴� ��~�1nS�f�t�]@��q|חNX�Ŭ���*��'"�L���P}�������Ԧ���y�SbMUU�! �B1�Mr��e�\]�!{2z��-ܛ�7�&��}u-���Yv/ƌ���0��g��77\��s������`@�m�0̳sv���r]S�)�slK;[X
U�NWuzAeel!/�e�p
�m��ao����q���zЁ0(�#����7Oota]��,j�}@h������{��J7����~��BA�OA��? �8IDq�A����8�)`�!f�"��rey5MIx.���hN�~R_�&<%i�O��U^P�-h��8i ��ѫ5��r���z1��p22k�8 �=�#��$��#"I�?V��	�Et���S��%�A{�e�@1�ɵ�&V���$qD��v4��_��˱���-��@x�4/
��.q�N�Ԡ�ۈ'-ݞ��uj�8>�@R���'|�O�b|��Zi�� ���+Q���4O+��>�ү8�������M���q䟽���yk�2Υr���j7����GUNy��ߝz`Qv��t(�*��&�b�����٫�K�2���:xѻ�����bLY�Bp��ġ���m�1#���N�d;X&�����4��fodY��}��/xJT��ڼ�?J}���	k7p{Ԁ���(�.tg9^��Ѷ|���C� ����˷ ۴]�F��6�\���W��I_!����|����/�@������H��i�7�E�X�r�u�- �������|�M��G��}V5�9F'mR��)���P��ˁ|�
lC�Mۅ�'79�M�վ[9Kf����O�M3��t�-R?sMR�D�Τ���I|���	 ��n^r"�H��0w4�%n(�Xli�i\�<A��(��C���i�Q\i�>6Y'��ʎ���P�U�⛙6S,�N�j�57c�/<����k�
XD�ui�Iˏ;�8�~P��r��;�ǂ�{9�w�$�9Sbh�8
l�0$����%�O���^>:����q��}e�S)�;8��v�W�%���
V�ASXT��e�9�[���Ȃf��C4 ���0Dr�ǚ�(nf�Wn+]�E���Gi�9��\:�cY[.�QI����s�}�U�GIK��uz����
�m�]2U}�h�z|��F��|�`�	"�R�E�jn�0����W����<ׯ�rH�:�bv�����٩��fR�f�o;��9��<�n�o��?�214r�W~�L|� �v`���LX��=��*_���ú+������\>�0�y>t�:#U�[X�|*i��L����{���D]�ݵ�-[�@�
I�@��\)��%���g��;ԅ���{g�v#�����T�J�:�_9zƖB��RK�2�Vl@Mj��Ƅ�VD��?�)�2�� g�vY�:�@|P��rD�mGP����|�3�#�+5��w��x�B??����6������S����{%�Gi�lB�.��M&��� !`LT��O��9�2T�!t�?�8v�kŦ=B�m�m����+b ��+F�	���l���Y��a̓KC\i�9h7qڑ���'$w1ԝ���� ���W?w��5Tг��Ғ�rГz�jd�����lRŇ�BS����y�[U��������H-��f ��A��CtX�n��b����I�uZ�0<����@�'����hSLҮ11���æ�/�A��U�'5|$�j�Mn|%�����F	w�, �� �^�y��'�6H��"�����!ʵ(�Z��J�� 5p��������פV�p���o�/0�r[�|6�<�[��e�C1�>��\�u��: I�bK^�n:�[����Ao��$��c���-���W+�G48v�lO�FXT�\#Y^��ȩ����a��Pscɳp\'��jZ�{�L5a�JMʀ����ume�l��{Y\v�mp�kP����n[Ѷ?nG/@�\ێV�?^'�d��_�,��'����E>��ެ4��m�:,u��M�]Tf��tA-�ꭺi��3%+Tz����\_M�F�>����]�\.u��O�#�M�?{��;zNxY4=.��!/��H]���j͎�aU#&�ߐ��W��g��xv��n���e�?f*�N -�k�l"憭���L�Qh������<�	c��5*z_��LL�E<��f}����W�E@��c�FLz}�:���2g�ip����\��J�Z��%:��$y����¤X���j�/�e�;6X����p��^�eN����1�9;�E�l�@p�O�;�]��!���,���~��#%i/�l�^+���@u!J,w�MS�?S'ޘ�?pj�Wlm��_���5C<�͜9�|$a�b�H\l���&8.�?2b�?wE�{��R�u`5�Poe�C�ߦ���<����q���ި��Qg�a����s�P.�*�x�����?��i~����5J���E��nV�h��ϴ��<���X���2�_�l���������ڿ��4nt�x�7#Zk���JjI��8f��V{�x�4R��ې���)[:��(���U{���-k�� ߎ�]��\c��^E����7�&���^��=C�a���cyyĐb�p�(ӧME��"{G� ����K�����_�Y��E�.Q)~��/p��O|�$�N�e)�:k�m�^�R�_.);�Ԧ���$^�����q��A]�Q�����h�k�ˎ�8��obI�^�VA�P�����˾�nX��Ѯ�'z�E��'K6BQ4�ʾ��ƚ����АJ�S�o��pPT$�7xn���}�B-��I��tFPu@��p�ol�S�&S�+�C��GI��W��ŀ���D�)�`��� �#�j�bv��ƶ{��A���`y�X�����3u�Z���J��:|O�( v�k�Xs(ݱ'}�,Q�?6�p�Xh���o��zn����T6�O����o8�P�r���×d�6�C$ɕ��X�e̛m�͌�z~)�� Г	�9���U�/#����##�B�p��0�an��%��Kͱ���v��<�p��}+,ٮvK&]:9Ҫ-Gp	��'�҈�@�^�Th���=�j�r�N*CD�jb�9�,�����]��p��C�ҁN��Ƅ��_
�k�g|�i���H�:f~���ZL+��T�}"�|�Tt�L��5���_}�p�L8$'�S��8�N�K�����r���_��6��Ѿ9��j�lT�&�u@�]R��.yL:�>�}nHNtG4�ۂ��ت9�z��Я>V���s������k-!��E���?c,�|Ug"�KÿXR<��w���it���|�"sa�@y���z�Z�� �gR���4>oS�ݾ�l'���)a�e��i1AV���t�J���.��aN`��JG��Y\R_����!=��K9y^�%<R���R�+t0�~^��w��i��M�'�|}�;3k��7#�(��&���/Zcj�%����d'4�s�y�:�~,���� o�y���a��'Q�:X�2pv`���!*� �9��4�r�M1�J�Q�͂���} {<O��&�Kl@j
/�Cآ�8�pk���[���H�(c��_lK=ʵ��הp��CI[�,��aы�l�p�R�*�\	�G便���%Ͱ�Y$	.z3���WU�0@Ug���~�A1�OK���ILH��40�#�&R��������^:��gK���3Τ�:ͷ"~a.���?��9�6���֏o�rZ�)�tߖ��X�ڦ�鞯�6X� �|j
���k�~=D�9�����ϟ˞ޞ�a���X�{�Ee��>����L��x���q���v�B���Ze0�W��N7��8�V��)��t�&�j�s��T��\ʄY����X�l��l �7�8c�$�0�r{{e6�9+9�r9��-oM�ڰ�q��]Z�k�r�1V�q���
��"}'�9'�=���]��X�c�ԶӃ�'�j�-�$�M��7M��b1�U���/�&4 n/�Q�
�4�k@U
���F{��Uz�p�GI|]�E*1���7D�$�׫D)����F�U��3��0�B�qG*%�C��{�����u�B3T@�(�S���TW�P=����j"�[��=`�����*��-�$
{*�Ԥ=�B���Pg�Д+^�	G�B�쭩z(�W��k�I��*#�'�9�'�Մm�4��|��W�|y]3YF�����-���~!�N�3���W��Z��tȻ3),�P��4�{@���&��y8	��o;�B!O|�[�=�����N4��`բz@E�SBP�Ǻ;Q����+�-c���;j��)Qz֍�`G�b�d����29ATV�_�]2ς&����a�&M��_(�{� ���o���L��Q�K�N�yz\��r��9X�	��V�ʲENh�Hv��j3���>�q��8�=�M��F0��9�5�z�/8%~�$P�W}%�����V��"{*FG�����U��z�r�P7��) �$��2��A��w�-B��NͶ��ք������^�ލ�j1R�� �Fd�G�͢q�Ԓ<6�4���3��p���;5
�I�`x��4X\δW�nϾP����;+�2D��K�}[!�7aE9��X�� %���J���ƉG�I�d��"(����eK�}���#w�Љ̒���И_��f���+L�h��a�H� �b��ϋw����jŷ�`��5p�C����BI"�� ��o�o�r��_�^�e�mPOą���� �-FJl7o�0�殆�;w��j�LU�%󼘶� x��l��se򐿱R((Ϸ��|E��:��V���؊��ٱ⧈G���=-_j���-x�)�2iD1��~����N���6[���|Eg�3�p��/�!Y�"C��M���k ����J���uCY���*?���_䩃�8Vf������hV����2�&��A�|p%���&<�A�9��'[���]3�4 ���J���Q&)��
Ϭ�d)���S���1���I�)A���ℂ~U�J�)Z���e*����Ofo�bG���W�
`}�!]����L�UH�将y�<.�*BkJ\���i����Ta�n�K<�O��Ǭ���d�xg�B!�dm�Ǻ���ϙs}��I�s�戜�M��k�X��[r�o��;n �y"������=���I&R�=8x�tۏ/��W4���"���z��nd�u�z�H��_���@����gH���7���̓P���T�A�`d�>mb�Do��1���-�MZ��X$�<N��a���o{�����U�����"P;��2rf[a/�_���ce�@vB�N�\"a���nK+T_�1�h��h5����M��v`�J��	S-t�Dll��� �ܹ�p�F9�	,.HNfF�ޞ�t�Y��@�wj��{e:}dd9!d4�`c�p�ؗ�AH���3�X�P�R���q�R��D�/}n:x�YQ��4�I�	�Sa�mi'�1:�Q}2�HV��v�u��O�%�l��7\��-��կrmk�Ƃ<
��*�6���g�1�I+m�:<ȵ�a8c�ZƠ'Bn�	�p��!��h[2����G3��M�t�`����e��E�)�PS�,7T��5W�~����g�}���{A3%u��?�(z�0Œ�i'חM��L���	"=0���ZT+�A��2���[�KF��i�0 ��b�<�A��m�<]3�Ced�t]E�Fu����\Ȍ���	��;u��;�E�g.� ���(�KkW�k�;�+57CFu"b2#%{���HN�����&���jɅ~�oZ'ٌ���S��/9=�Ի%0�
9�oo�T�ۇ{�.��TbH4%w�^�,�h��I��[��7��3 ׁٰf0O�n�a�G���2��R����Fix\�UmR�jA{5R8ضio#2�n����,�@�[��Z����ᙅQ���yظ#gI�sW�ư��詳����$�Pz��C�Oz�67ǏO�'D�~�=�?̶cm/i1��rJ�܀�vR��~���N��B �M�l��C:� ����̓��n��cC�jM�?3�W
�?m������U��H�?���p��O��22�m�i����e3JEw㤾7�����zy�A�|�U�.����+K��G�9��c�5���z�n���E��0��4��^('	�ɮM����kTF�36u�R����=�.A������g�W���\ə@�N�h���'��1�t]�mnc�1j�H���9n{4�Է��x�CR������R�Nӳ�ulA�+DO*\E:R�
wv*p�����2�ظ�9��t�i������<�U`J*o�Chb���]۱׍�*�t���e5{-��x���#�nO�)J�|ˈ��Zԭ�L��.(�p���f�҈��_���9�D�Qw�@$�Y��h��|{�7I摨fտ8.7%�w�Q&Hq%(" 2NZ�ĎU��";���4�Y�1�lK�le�fq��ٵ"�wt+����tȨ*+�Û�% Ci���,��;�J-,"rFnor�KCf�������Z1��3u��������xo@�g�X��Ƒ�D$�Tn����6'��A$f�2�a�D�\g��μ.vOkm4�r��ٯ��&ց�3��Jk`eu{�|�9n��g����7����Ե��B��-$j
�s,���y/����~�+��	Tv;5%#-jz&b�( N�+p��k�'��0[��w� #899YR��<NoI~�$�v�	�@����
G��Od��9��}��Z�O�v&�3c�� rA�Z��բ���T]�LY|e-鯞�b�nȃ�Y�=Kx󢖂H<�n<b����?c�&�R(��%ܤVټ���ځm Ղ�[�3�J`�N��Q�LS�N�.�,����P����?~Qk�/K�ptP.E;$��2,������N�Ȩ�"�b�}�ܩ�8>�ߛ�c@�;���-�s%���,߯���E�U�^{�q!�$���Ֆu�R����*�91���/p��R}©xq���w^a&*��ZR�r" ��~'}~Fv������?��7Z¥���F͇;ŉ�P�b3[Y�����)1x�Y�g�N�0íF(F�z8���p�l�&�s�P�O�1s��	����8��r$1�����b|R��1K�`��'�ذ֫6�?�0�����V�ˣp������T ��0����V��S.�*d#��I:#��;��̈́��h��sz�jdX-=J�o�fzܭk6���S�+�������@k�x��P��P�1[�`�m��A~�J,_����u廴i5�ӕ���Y_ '*w0�����U�����A���D	�������U�fe��I�b��焩���p����
	��4��`���Z:����M���0
S����3X)�����o���$�6*~7�v}�NG�S&WpZj�L
��ɹ�sV��$mT�QE�P3��j��+K|�hV��a-��P�_��</Y��I)1}ʺ��^V	���guF�.�s�h�����3�[�&'.���j�5m�/=8Y�}.�On�����|7�\Q���IgdE�w�w89�x�\#vi�a�H��"�}hG��G��0���#�|��k B��ӟ��ȐT��V�� �]t�z�LG�B�aI���-Y;-�N���j(�Z�CϨ���K�Q�����=V��Rq[��������=2�B��`:�+�=
�\A=���ʡ\@n���~�Ȭ�"u��&<P��[�ܘ(�"*��gH����qr�hH�0³�>�p)$�Q�����˚�N{����qr4��$~-ۍ��.�(�ur�^%�6�ɠl�L^r]�y�����X��B>�\�E���|>2��?�3d�VV�	|��-E;�*�FIYY �{�O}�
�� %E�M�ʘq�����&��c �H�mzg~;�;�	DH�u��/)��NNG�Q�
� Zr�Q8��ꚇ�A(���{�=v�t׿�.?B��1�~��a�#���Xw�1���͂ǚ8�~�c����k������Mh��k����۫��*3���-0'�jZesWt��[�@��N����g8��y���gQ5���	oN��FiLZ�����P��p:'e�����L!K�]�9È>�R�mD�$�:��GsD���|�U_7��U^�@�@���z�F�l��j��"
O�T�nZm�\�W04��(��o��XWbgZ� ������M�}������P��D�j��/ΰ�G���x�ϺN杯`e��*7��J�<A�������e��߆�M�J(��8�j|a� �M�F;;�$����w�u��XTY��^еlm�n�9��׵��L>�~\�Ğ��4�e��3�X�t��OM3�j�Sc�xʴ��y�vv�/Kq}q������U��"%�5u�A	R�	,��s�u.��4m���G����**8�-�4t9g{�.0%?.~h��:ʧ�S	��0/��%�1=��f��P��U}��gye�㖕_��BJ�v_�T��2໑�@�&�h�=x���̉�<!d.�`U-:�ʒ��1�[�����
M{bZ貵�f�@<���8[6�S-i��Ir�p��kZix~w�nqe��:]��׀�ʝI��
�, v�C1�&*=��#���Kv���%�#h�g�'���E֊���n
>�����6#U��xH�+%:ZB]gk	���d��)
�0�<�yG�N�|�'�7)TI �
�0�n;�h`4'��%}�U��<��nb�'ekOkUwS�ڝu�(�R6�ڂ��K�׳@W��K�0�qdU��W,׶f�d�d����[�?LW��>�����fҎE�f�\u�h��ָ��`��v��f<�٘NC�a�wA�<��1�J��π��;	8�<����&�c��E��V�eW��v������3��w-_��nO���ȁ�)=���m�&�އ1V-��yha~-[ݚ`�8��*�̞�.��1�o�KR�R�@]&���i _Q�F%.�"�	����g� ��eN�@i�1X�m�~�����=��@+
�@��N��;柯��&�_p)w�)AMz�FWQ+�I�P�b+/I7���q���D����e�3r�yS$�Q͙�_�#�.�6{`F����%6�y�uA˅���QʓC#��H��#h`L6j���0*W�����K��>0ST��/�#��~��PiT������
��#�1B���0§�z�o��h:JC��ѱ=[���#đ�M���9ٳV�%�ex�֚�飗���UO���eڔ�i��<��q'|Lg�zCW����j����PT3��4����<1�-~&�9�ӳJ��ޠKiS�6�
!t�"����6���7a�� �O�e%#��i��4O��S��fy��d�a�?k�q�V�\��)i��[�t��w�L��!��	�{�u/���]��%�(�Ɲ���$�Zf���K���@ϫe OqsJ���}��C�)��q_���G�;�����,9��6�^��U���ޜ�K[����o��s8t^t�j����-�r1��Jͺ~���g�h@�*��]��� �PW��
uB��fr�K�;�JxA�JHu�T���g��4@��r�H��T�� @���Bڔ�%�Ւ�Òۮ�|�*!Hwg��l���Қ�9]��<��-�8F�3)nay H8�X/C�s2��]V�
x�R�J-	�����#Xٻ��מ�R���U�y�엀�z��_�F$ s@<3шlAa��
�%(T�o��Y@z�4f�D��$j)���FW�3�a4� k$��;(5XE6���cn��9f��f�.(�nI�ZH�d�-��*�u��9俓����*�3�	��ܬ}Xv6�q\J+�h��Y̴W!m0���y�4YV���kB/U�f��LP!��*�9�恂N(/d�`V�_Ii	!��q�K�W#��*���� ������\����Y٢;��7=耨Z�X�YcB�E��Dd�8�����Jr�8�^cYp%�3gi��0d�ל�����g��L�9�[��
������p�J���I4�$ҙO�yOT��8,:��_|��7M�L�*���\!��:i�È�rQ����o�OHL"� ���`����1�i�G���=":�q7%H2iGC�4m�����ug�[v�^�6&a|̎��� J�)+�P���F|	c�}��`΂/����׶�Y�	)δ�����m��2��%���С��I�}`mJ�t��11�c8`���T�_G�A��-S�T21�{�����0�ڳ�}h��l���s�u�z�TJ�$I׈����Zw~���X��`m�����+�E�Fx ��D�(�\׊�w�ؑ�M�����-.��U����J�-�hj� ��)9|�THC�ulͰ�MzxG��O���-���2rכ��
h��A��^iJ��<E�Z��el=P���?���A�/X����~�"�(�H�~ۘ]
8�%�gcgC��HT���.f����	V��Bm���P?�i����Q��fS���]���R�C`�%U�ʥ��>�������e�͙�'����|�Β,�?-�>�%������廦��C�KN��A�.��`bo[����{�7�h� �Q$j����QJ	�l��a�4��0+R\��DC Bw���?[�����ō�?���%PgJ��h5Ln����b���HK_K`)<o�$�>����*hѷଛ� u`��S_�'�����oY���{��4�e�"5�w|�V*z!�yJ��}P�F���1|��s���a ��$!(���("�6�-Z�u�|0�?7[�V:,�&1A�Wz��0�Á����:���hD�����J�n ͇���>Zֿ9�J�n�������3ef"÷���Z�G��Y�/:�d�4��Ր2ԏy6.\3������7�
ET,�3͙�3Cw���~&פ������p���~%��o��A� �V�W�Q)�'G���U2�<#����e��2�Y��'�,+��>����ϐL�'&��_���;. ta�AF2DNһ��EE;��H�ηTa�
�7�7����D�7}c�RD���!Ʌe�Ho�%��"R�����@�hV��ؔDXY��>\PL�$	���ƈ�HQ�������ZK�b���/�S��U*ŉ����F�F�+�:����fUqlO�&`4�y"�}1�
�J��S��3�wHed̅���Z'���#�IR%������!�Ph۩
��B�_-�#�`�[ ���6���I�5rz�(��>����$1��	㷇VFo�Kњ
����2>�.-���@:�Q����d��w��M�I}�>,g�`���o��t���}ඍl������	�DWS��]�&�����(ʇ�g=`9F����˄�i<�
Do2�3tb�W�_�R�h�-��>�S�9��vl^X��s|k%%�2_)�fu6��'��e���u�Y���K�?b`�ԕV<�pբ�@�K�6�w������n�M�
����-�1άr��5ԋA���%b�&����z������C���T�p . i(��K7�&�vg9� e9���H��3Y/�����:J,!�t��s��b�>���0t%Je�զ?a��L��OY�A�"ԓ�����"^�(W����l��}VL,���H�f��7�w�(�kkΊ�
��OM��+�ͷ,x�̩���C�UK��)���;K����Y�{���Jj^u���
�^>F�-��4�ճ��5��nP�P� G�S��"�������}Kn��K�k����7� �5]�	�P�$��#X�D��-��KQ�Ƕh�V^F���zq��M��ה��\�>���qЯ}� :/���(!�o�H���9���g�.7�«?�����-���:w��Z�};��d��\}&s۸�=�o�N������w��CU8���	��Σw�?ǂm��`�tjJ��:�i/�]�w@C����F$R�4A�
b�#����d#��̲��웁�a��� K圃��<t�\g*��ׄ�BϿ��"^s**7j͚6)���?�G� ���L�Z�e��2N�w���\j�,͑^��k-��*�j�Q6$�(�$�	x�@t	����P�Q����bBc%���ٰ������jI���Ŏ'�����7���v���gAb��	c1�]�|�t'���pڵ�h�
Z��S��ǖ���ӛ>��?Y�hf�*E��M��M���s�(=L%T�{i~ a�����K$i���XӴ>�iݬ�z'x9��͍�!�[A�[��d���k{���EQ�9�5������"Җi�y�)��"ࣾ7e�<�A.eN�k�>�����[+Ϗ����r�ϷjGm��"���Ѱ-�Աw z�������~!��@��P�Ѿ=��i�Ť�b��/�̜y"Ð��+���#��b���҃{�q�����!��F:�sn�<M�7%�.h�IW� ��q�����v�x��^x bL1��(MG��_E��%e�v�����fi^��#����=)��O���+���z����c�]@1.W�>��d�2m\7ݴ�T�����0J�~w�-��U��P��X#l
���^k��:�<��g�<����I���`҉?��G�{]�o�1�o�7B��M]��F��C7d���!�
T=x��.ّn��4���(�gzӷ��|�m��d��%*r��/���7�>qr����zwU�,�,q�!z�J�o�C=,l�%
�(�� �dq4s�M�>��x	�nL&B|��Rf�M�_�̈��ӅF� _P�Z;)�lp*�3*���&�����F��H�����M��{���H3}z�x�,���Yz��G��3���N[A��N�DY�v9,�|�i,H�����Y�M��ڹK�N��=�Pȋc,�iDN�"l��(���҅g3��}�r�4!�)y����
>B́�Hm��æ�$�מ/}"�}�{޻]���5�����m`Uv���A�;ɻhH��
TzE�r*D��q.����ǵ�0 6p���@+A#��w��sk�!�:J��t�R�����F����7��a�"z���Ir�2�����K���Z�I�s�G�h�,����lV*���oj��L�\t�dp���x<����D�*������;N�̮=�.�M\p`Io��9�/jV�Ƕ��oW���=]
/�Wr�}ؙ���ɶsc�9-d���N��2�0�KR��N%�3�	�oow:��D��7'�̶!,q��~T�z��̞?��)�0nƸ�laO��х��j�|(v�>����
���,�RI舭��AA,���QM�,��S�2ɚ�I��_Z8����K�\�ɔ�r�[�eh�,d�y,3�/E:�� b�I��`-�lԔu%V:/�=��Jd8{0��+����1y� `�Gm4�}<�LǇ������_F_,=n�D/ �5;�R��v�K'1�2�K�On^E��q�g��RS�Sa4cT[�hֿC�l�L�����rk��R��4�� ��ŗ��͌UB-o'��2`���^ƐP��ĵ�f&�j��}A;
�X5��rWH�(�*)wQ�a�[����������S{徳E��(*N+�쫓�ɿ� ���2���3���ò���5��:؎2 n:��
#Ees\�c}�.�=>�ĥ�P�~�:�e_E�$�[�Z�$u=p�x�d��Y�<[�A&���WǍ��PR�9M'<��Ρ(p��s��<-�p�V� �9ɟ����� ��ry6
�	������ڧh���Kא%���i
M�i���P���ߑ�s-���w���Oz��)�l@��vg^!W�'���@�thL�]��q���Yйë��X1���1*�[�Qp��s-Sd`�>�<��i�I<�K��n�
���.W9҉,>�^����4[�T�-��f4E�F�q�0p��df����qm�݄t���E&C�d,)&>����1l=)�F$c��V�I��%��̓f�[�M9��rto'������+���C�we���t?d�@$�����h �Z�$5�-�Չ�u�i�����r��a'ف�����S�Jk���Ш:�	O���ڬIP|#�.v��|���{u-Q���H.la����u.�ݠƚ0��� �ö���ֈ��.[9)�k�y��l��A*k�*�_�BfO6��rm\��a�9�#P˧��)�V��ؒA���Z�D���(�rS�aG|�Y`��K�sr��~����%������Il��I��G��N��]׳ۘ��-GhR���<[<�#g��:6v�J�p��ՈEi����D"D�M�� )v(R@=��9a��u�?��NB�]�����9?<~�=�WAF����63������w�utq������/-�R�<>%���ͩ�7�]Æ�Yύ�~�t��ɢT���x�<J��p�'��lx��d�Q$��� ��%��<0/E��]5d*�4��tO"���Z�׈��׵��R��0�G���`F1Ɖ��"4N�p� ���txr�����K���q���ɷl��6��p�9���v�Y
4*'����P� Ë]�#B�Z�ĸ)%��	Z�ig�C��CIJ�> +���XI���0iG�Z�8D�bi�<@��վ���'c@�K�֪��q2x�@rz-��ݔ<���=�A�������n@�u�_��ȸ��j�����爞/�Z���]f�P��y�oe&y��8/њJBB%�['(s��Z�y��r�h����T�Ζ��ހ; [J5m�" C)
+5�E���
�z�o��˰D���"����Cz���L�-��i�r&j��n��#����!����N|W��ؒ��� P�[?b��K�/#IV�v�]a�cg�4�of����4�tH���1g)O��S�:�����~o1L���H��[e���,���Sߔ��7�k;���D���8-ax2,X�]�aכw��}̺�Au�$v�ҷ�+�cuiD������ϗ j-\�OL�
3W�L&DLi-�F��*xH�ͳ��!}�������Sꚜ�su1�ON��᳖��u�>_�H�:Y�5��� q�� ���C�����ն�\�Z[},G� n~��Y)܂H��=��C-�ů��a��4���2j�7��Gp�͏D[Lh��n����dv1�W� ����{����4����r1z����Άbg�*ew�z�U� �k�U'&^Z�4�P����(�?��g�@O��,���6Řc�K�Sib��f�n�)�s<ߎ�k�WZ���aC�>gv��j�]xwmu���ދ�@�Ք����uL�E2	�m )R�����rdIZ(a�pDC�4��I�`��
�W����('���q����n�)�n,��9Y���Y�� �f	�d��쮄��{I^��Q�9͌��zk ��)����-�Я�jذ�ğn9�ľ�&'�}K�m�]m��7�z�"�FX|�l��vq rΫ~KkL���â��U��*���� (e�N9����p��D�KO�$��y��6�7=_8���*i>��Uoȳ��k�'�{�e�d��)َ�Ir�E����Vt�K����b4�V�3���H(�o;h�}��t�����z��a#��w9'�ɉ&O�����"�ﴗ�d;P����	?afg���(�Ԡ�.��$�	�؆��Or��&L�j���g��Y��å ��P�Ǻ��!N��=C_WOؔ(5���&`e�0�sTQ(��ǐr-!�I��B=p�~(͛sh��,8g�;_�٬H���eR�����<�K ���d@��:�&vG>��	��SO9��T��V����S�.#�Q�W�M˰���-�M��f���y��ئoĊ�/V֌��:0^* Z�y8���(��cց-D	~a{�T3��֤�_,�1r�q� �ۥu��DU��:�`����X�R~�@#a�	�%&���ϵg�,�]����G����K�2o	R�<0y�j(�@pV	��?q�+3�!qI��%T�+ca�T"+�B/z�p>�Ӷi�.��I��+�B<\ϔ�O�.�*D���f74*i	�����Al�)��Y���rB�{�K�^M�O޾�P�T��l�v�k�VJ6�!ۈ�#�'�=���rC*ء��)UQ�,ֿ�ȴ-] "�꟮W��9/�$(ԏH�|�
|	���A�<�^�yht)��!B�~��j7t�2��Ɗ^�����Bac�ŋ�����d'}�4�O|w}�<��U8�J	k�aY�հd��x��o��U�����v���e-�+�q�OVIV+QɆ�󐇛��Ô0֔-�M�µ�������?j*�d�<" B �2��D�����:����G� �)�-�l�������n��̶���=!���EnXLL�&�u����W1��zd��q�J������A���p�icyrW1�j7���!��R���x@�
xcv] b�+G���F�rS/^�[��;Wǌ"�hbi�EH��]{���ᬷ�BEm�>S7=,�-O��D?&y�	RT��0k��e� V��4oG�q�P����pi��q��4ear,?X��Q?�B�S��_�f�����!V���ڸ������)JQ� ��/G+KtCH߭n�_�Zé�C�Jp�߮�D�GA:~�Z|f�2q(�jwL���d�4\��m��W��t ���
�>{��up�.
(ؙ���3���'�A�BtȉB}��v��O����0FU��Q���@�6�QYi�P��	8���Y�ju�֌���0�U���_�ͷQ�K�9��[T+��d:Ւ��<
:���9,�k���m���5E�?l���!H��!&�������"�s@��Y��<�T�5��ѭ�bx2Ч�R�|29&���V�����q�;���S��1.k�U-�I3k�?!Ir���(��7_�U=���aMk�=Nl�S��XGKr�A��'���ˮY�=�&!vt"M��H"��bہ�\��'{��ѧ��u��9��ȡZ���mxm�&C��s��`�G��S����l�>�9��B���U!`�8�ONd�x��J�/?S;�?4t���(���E�Qɓ䚩��>ՅM�	[��fh��kLC��T�� 3���$X��V�����=vּ���	s�1�h����չ��PqL���Q|�O$�2gT/C�-"(��|��d;��h�|I�t�Ov)�]��[��z�χ ��C�!��U��_��*��Mk�_~|<�PD8;'+%U���1��q\����0$��ML����6�i��ha\QD��U����,�� �nd7�}���C��}�(g�WT�!6����	�<P����/,aҠ��Ǘ�ɨ�S΄\����"�@�,V��[��{ы@)��+o���9�������Tٰ�_{��Ҝ��G�Fw�2��`�b��4X�=I������K�"�]3�M�[_O��߳�Ǹ�f�p�/��|̧�u6zǴ�ְ�<��]`��GG,��ގ_l�+�� �Ȥm�rc�sb!?�p+����-�p��˥q:�љ#�d�f�1�p�9�v��eټ֌|�^l*�Hϵ�����W$զ�K���ۨV
�F��+��� -��O�=i�g��#b�m`��H�tVO�a���n�?X��<l��A���G��?��fJ�-F�fu�x�
��X�-̀���r�*� ��'<�n,,ʌ��v�1�	p�i/Q�5�*W��,���[Ï�`ӆ���s�Y$>P�����Ԓ�# /p/st�%�;f+�ѹ/�0_�n��s���P���_�(�r~�bg�l��e�o����'�K��4��a�W�<�}zS���z�P�lMe��?��[Jɑ���*A�T�΋���B[c{
f��iXH�'Δ��3�~9�)��Y��F�	�LM�Ց��( S/y��@]?D��H/]Kn���	Z\��^�y%���3f�*�kP����7!�<�?+X�uf��4-B%�ǅ�{#���P�|��sKiR���7�*��ϱxE��_��z۔F�IL��|09���ć�'i���yY�����ϝ�]w�{���\�=�x�bK0 �ب*b���VL���B����+kX+	v���2�0���9�#�QD�?8��w��,�����a*�1jL��\=�)�w���=n�9�Y��FY���-Țv���لa���=&�zJbM�
��
MC��8-q����X{lZ��aC��뽘K�+GN����&�d�CJÞp�J:>��|_���Xn�t�\7p��}&ZgH@�>#v27,�)fs�n��\��xz��eW�Z��űw��.=b��4��sh�C�j'���$g~C.3��)U<8�Vs\�^��. ��C�>\V�Z:��gɿ:ՉD
m�K�����6�~�kR?DG|5W�Jf�(��s���][D9$���H��V��n�
g-�8�47��ǡ%r|-<�N�5�<�:��8�u����/H�.eH��H�������n����2
�''D�� �# Ņ�/���)��UD�I,�ћ�"A��[�e(���8)�-R�]��������G莼�8=~��׆F�bF�l��`Ō�?߹��3��Ƹ���[.eW����Q�=�l�x��0�;�P����5恑~�h�	B�Z0qk�A�_����?�èw\�yN�D7�����8��D�
ƽ�0��(�A�9En�q�����M�}������ߦ!����y�$밵��7�Ѩ��2��U�m�x�1p�3��*���}���Z�i�m+,���<U�օ�)>�lZ:³���SWo�z #\ldy�՝��3]�H4ӥ�8�ȴ�}]����5Z�)^���#/V�#x���HUFϛ�T�������{�2�{���'H�\�������H�	�
R���2t �<])�:���ݱY��
C>�`��p=�����-?F�l�]�L6�I;�X�G
+�ͭ�"�3��o�c��vt��b����f����ǫq�"�%?�����O'�-��^v��Hi��I+i����]ݒ�]�:����-��\I�H+Ϳxdhg45���FNd�g�r0�������䅈�}��(��D�뻖�`�����c�	� _��>¾��慴�T���݀"L���b ~�t��<?k�-�/p�$�i��s�9�<� M̝n����V�_>�9��,��oWx�T�D<�b���g֣�m?<��E;��>{r��>��f:e�`����6�uG/E�!*�>7�v�/����I3�y���7^oC�G�Wfݙx�w�WWх7����eՀ�L������5����o�.�=k�h��|�S$ִ7_nŉ���dc�L�+���GO6��rn6�������@x�/Q�G/ji��'���ԗ,�z6�/��}9m��蜔���T�{��yV�ؼc��1�9/�k��!7.X����'¸A��X��h3v���,�H���-F�a��rZ4�e�{�G+���E��L�<�QYt�����xEc����I�.������g{����s�>��<_�3e�����:"7~9B�t��+�x!!og�g�X7�p�@�%O�=��s��B�
 ��2�������a��Ox�ِ�_%/� մ�+�r���zLx�D�'���W�j�NM�SxQ{o��R�7Ba��a�:��v�[[ԅ6�f�����aRb �X~!g�#�?e�7R�pb�Ba����&a[�ӥ@@ѳ���cdiv�&`��������)[
0X���)�2��&4���+>��D�� (܏(:`ј�P.s���ϭ��{��E���λ��	��R2[!�V��H6����b��s�P�kH-�߼�����0��fؾ������:SŊ{�r]�c�c_x1�w�;
��ږ`?�V�7mm�6����W�2���{z:�8�dFc-��&����5�q�?_���{����Z< `\ED+=��9�/�u�}�����r/�΋̡�KO3���z$Z1i;i���'h�C�ҵ"Z7z-�	�A�U�^:�X�߇�H�
bG?����s`?4�����{R�lT�ܵ�F��B�*5��|�O��Gݥ�{� b:'?(~�`a���[���Q~��P�uQ���tu�%.���p��ڄ���8,��X�*x�0eE�2ܙ�6�Z���j\���w��`Y�[�C�@�G�N/1�z+�t��f	�ϩ�6�ܾg����B���p�b����.>���G9���p�ǐ�g2��0>�*ܬ�m�4Z/�D��r��YΓԠ�q��^E��g$�����n�z�&��*4h�R�7��;�*���ߗn&K�*q�/ "{�l���U��[^|�A7WnTmb ΁�}�][Vh$G�SY�Flek�[�J0jP<��?w������v��b3b����k�D����1�(��M���¨m�P	�@���+_E�8DD�/�j�
gr�m�ܵc�`�ξ�S����N[�3���߂�@.�D�{dZy��xЧ��������$e:��؁Ay���k���T�{ֶ_v�g�N��z_��u
��� �y��2�Y�l�]�/:ϵ� ��z�E��%?|���lǬ8��9+s�l�m��������k]�_6E�e��H2����h�Y1{���6Ѕ��E�?�;�Ւ�`�D�]Ek-�K$� ��gZ�"{���^	S��O��dU������>�()�U�>��qM�n���oV&���9�i:NT�$)[�w)����q��O����6�C����]}���6lL��Ԁ�<.XPS����<h��UH�ܓn'����?�_�X# �АhDjp�>���Ȫ��>bU��1;�fw����Z�GEݚ܏�-p8�_C�Za5��,̞v���j`h����I�� ���Ń����������1�&��;���Q��+Q����T������QN��A�U��,'�{��#�4����*���Q�d�
A��M;��&�ľ+n��:�X�OWY���?�N_��!ֺ��s��Z��dJ�C��I���g�2>�$�?=����V�x��@J�qLƀk��(�܄�~���?��q�(��¸�@A��	r��h"r>�A�wy?��,��X��bl8������s����;Q=�c�r��L���д)8=��L���l��u��;RdI/l!ONW����i�FT��^��O4��R��v��np*�r�c�4c�i���0Q�4��|3ݞ��W�vVh�R#oэ;f7�����?�<u��,���k�[
O!VO�	�|�$K�������D�7�$P֖�1�~�
�_�QB"�'A�Q×�N��w�4pf9lxl�RN��O�E <�ytN?�#�bh�!��xX[�9�%k ����1{J!B����0�Xd�R�\�3����P�$��(|��3��<Ki�S���e�Li���_�f��R�J��,�ըW�b�p��4��yK@oK���
�Ǌ:N�/����⋄�����C�����B��ﰸ��	�R�j6�
e��l�G(�����8T�'��N�	��!�f�yTjk[�C(���Z��!�l�'�t�g�T>D�7�ku�w�*�`�����Y�@�0�21����}8?���kY���W�DnE������毼�XAڎII�I��E��%����R?7����D͜E=*�A�֨�շZƽE�Hr*!)k0�f:l	���<i��[���g���	��襁*�}Bj&� �^�O�hܽ$�fc8�P�>��Xn�T�t�q�	�;�5�`����3��q��@��X��Rībo����m2�o/�(���w WG�o�Z<e<���X��O#�5^�]�}���VgR�J����P����Y�s�3��pW^[����4��)kJ�)��0�xj�pgAYE��s��[/�#��F}��y�����*��:	[��I�جm>�V�u(�����<[kw�2�t%�W I?17�����r�/к��E�*k�GI�<�%��>nC�PȦH�{�D�DP�žq�|Nb&�|���g)��~�� Y�^����1��I�x�����6��w�m4�Jޟ��ðz�Pr�?ץ��Y��ݼR�˺i�����%*���|��JL�	�.�yF��U�Ѩh�YU�|v�/��� ���A���c��kn78��@Q�G��n��'�Ė�L��&[�@��;7\�L����{P�g ��]�3&��:u�E80睆緟Z-��
%|e
�O�B.r��TθH\.JF�7n�=��p�+��L�G�W/�\���dX]P�Y2��_�"�Y�'���ӆ�9�[�m��'�Z����(����3#��`,�}@
�
�˗C��Y�B�����(�г5��[[�_��/$z�k��ήZ,�t�r�:~�V��Q�����V�;S`D:<��:ti��C�yb�G�����#e��xuQ��0h��!���{��̌�7p�R~�{m��|h�G����}�L�j�Gyl��n�zE�~�UP��`F��9��GF�fk%g��_�|Ȍ��37����i_�I�ho����<��9�KyB�����/��
?����j����#�X6�&n�������\#.�Q�:�/��Uچ�s�F1Ci���d D%�F��KeB&%�S��w��B�)�,���n\7�O1ƃwX��{BĹ>� ���3�eCƃ��\�v4 ;�78�`x��{����/��2?`&參�27�;?.���{v̵��G)��E_��е�����c޷��?�w���1�D坮�~e�<ɜv����$�Z@���t�5Q��O�Af���ٶ�3��Eu���w�D��
X�)�C��OSy�-'-�7��<ϧ}������P�� `��
.j|mC_^�
��r��M�)�2�`�EzL���Z�y�`�TMЇ����#�*��w�����9M��#����������1����#�����U?�\*_���h��u����=��A��U��_Ԋm"�57�T��֛i�}n�c���)��"�����3a�Y	[��oޣԫ�q�)�j)O�� }��VJ]���b._���)��cx��A���߮��֧���
)^Ѣ�o�&[|[�_|�o��o�Z��&�F�a��@���\�gQFS�är��5���$�r�^������ogLi_�	+���Uʄv$��;���<���N�u��(��ބ�@OL���&�۞b"W:��O���4Kߎc�Oy�2$��&G���*����ki�#��r׶�
�Tݙ�S��sY�H�1ϖ�y��dͻĖ�^��^h�u$��%�[��"`�d�3Ǝ����,x��U䢮���ԎA��;�^�бU�uU��c�����ZM�ӽj���͠�!�6��2��G�����v#d�	t�����
�()��*ε�~g>�]��� ��'��-�\A��*�X2з�A��{�OM��F]{�Ї��Cc���A�	���pu�_�m?Z���zVu����_�]�NbS�"��
��@�ќz��)���y���E宠��0s\�5kn���Ҟ(^��P#7�*�OT�)�HzD�g]��r��T��:�r
�)� !�̦`����`���w�����^a}8ϱ���in@��n�=��s]���y;�D�QM.�����z/6��X����� s�b�`vR�m�<g�Z�� �}���>�č���՚ 렦�<l4o�v˵ r�Y�o��ލZ����P��S�x�8M�m{�}l��� NL�}{�)�í����L8Ȉ��ú��E�����L06;������RKf"�E��÷:�����W!~�e�S_���`a���>{����=5�ſN� �%�{���>�K.��__M;��M.׷��2��z:J���Q0>Y�Q=�|��&X1c�O.�}�9����NXlr��Y��UGL?��d@\n��ˁ�]��T$ΠZ�2�`W�u�%��:3�hܫ�lPq�5�nB���y��	2Nd@i�J{��K����C.����ޫ,�;�}��/*�-/F�����[��vߤ;ܽ���ɨ�"B��u'd��lj��+w��oL��w���ޕ�8O:jV�]ů<g�xm�?;��7��ԹZ��u˽���|w��]~&�{���\b�`,t0L|q݆b<1Hĺ
Qr"Όv:��p�N`q(vZ
�Ķ��=dN>�x]>d��R+�Ɔ�N
�{�5򖳨-�ʹ޾aW�<�����^�i���9�-�o��EzR�#s�� VQ=��Cʱ�ё��lOM��� ;m^i��D��1�	����S��������OC|Bt��+C҅}P���:FgPy�)�-�l���Nt�)6�1���K����jހ�Z���a�ǅ7�X��}��DS\9�X���J�b$LmU.�3�,�z�ۧ\Nu3MJMJh�*#�(e�N�BC:��@�6�q��8�E�Z������lF��`�$gg�^+(bx=mS4pO-\�$�A�������w8$� 0g�+���{�@��j���ɀWGG�X�̓�
�]P���}WM�Be/�s�"�V�ZB1H���s	ZP��i�Ԑ�K6ƫIi6TS������;������nD+m�	p+�n�CB���vX�LE͟�gZn����b�OA:��(�����2��t���r&
ñ �WM�i�A�w_�H�(������a�	-�[[����(��W\�(L��1U@ϚD�p.��t?-8g�����r��i��2M�w�[�f���e�@�.��p.�&�	���Vț�t��Vm�U&�,��u��Ͳ��E�iU咢r�x
���Ÿ�C�O�y�h  �N�V�rY�<W'-�iLAae����n�]ܑy�KgS:R&
+[%�B��Z����V�$��:�͍��e��Ͱ��`g����,������GIh���O���&J�LwLJ*2����B����������ѽPǾ��]����H~�����WzD�c�Q:��<�D���ZІ-��R��n�|I�7P�R�{� _/LY��	�I�QFcf�2�<�9 ���g���f�{Se�nϣ�f��]�sg�j���	���u���̺�U�je�c�g�4�ŷn�]��-����v��P�����ԋ�~4�#%m2Q�8��%(ֱ��E�lnc��o�J��of[�a���ɘ��(�i��xE������Zp{����	�ϸ)�7�J�n��<6f<78�|��X
%4�H�����4�_����������.�d~ٱk�|���;���K�}�oz(�� IIǾ5Kd�p�	(�^�X=`�Oٹ7�@Ip:�
+�<|�@����/c2�Z!���A[��*�IYW0�:	�-yk>�Y��x��hBc����tU: #5�L�ˋT�E�gH��VxN~��ٶ�}��^���#H{����]-��e��",mXIDh�/��5|�R
�����[�H����k	������f�M�A�#/eȮ���q����z�v��E6ؕAd�>�N�&������� ڭ�Kxw;� 	@�@%�Ky���M8��������s��ۧ����7��aE��[���1s�Kp����5��H����V�mw쾀ˣs���"�|����j��{���4��B�˜�Q&����)�_��vh�7@h��x��4pD�M�l��ַS+ŋ�ًmT���a�SӢ�0!�R�
�c{��J�	�o��({��2�F>��M��i*@6�n���jM�Hw_�[-���){d���4\����� Q��GW�&$��aqa(���#�257���C��w��߽�.��w�,\o�����4$�A�42a�
+~	u�:)y���c��,���)um�^
�j��W5��@��*��'h!����j՛ϧ�1Y�r�qD�]=��J���"�ʬ�(�d �[i��Á���dw���sҼ{�'b�]iv�#e^=��.3�c��,. ��
���	�;�-ȍ/��Z�7���'
q'}��v�۝��\�DQ�"�Y��uH,�������X/���(;I-�!�@�U�{�
���w�A��#86��P�1z��]r/�̐K�=���m4�2\sH��Ƙ�;�ұ'GwU��:݌��Џ3��]�I�G����	�yZ���P,�f�e�e��t�M�������M�H!�(B$��ܕ�V��1̙8\�۶����G��eˊ�O/�URRx�Mi���D�I�ǌGqJoгǮ����@�OeOz\�~t��D:z��5K�`P�.���R���Mƽ�7�l�����s��zJ%]���L]oAN�����E��L�"����?�uOFuE=:����a��#)n$K��~y��~����Ψ�]���T���T:΅?�2v&�;�����O'S/�r��oǿ6�]j��\���^�n��r��a�T��xﱧ�b
0��5Ȓ{8�7I�����T���&ٺxMv�0����	�:���s�7����kܞhF(4k����x4�	G|6I�)���#�G�i��~��cC)f�a;�35r�k�c�:�T�\<�G��J����N��j�Y,龐B�O}>ڛ���j�9��[[�/d�%���icT��i�՝�,|�(�")t�p��N�x�E\ƺ� ���?P�
$/�h�@Y���tuHV�Đ/<��U���O�:ᣎ5/�B>�@G�-=�:*A�QK"5kb���9���dx�~50�9�U_R�]���������X�M+�𙮧�­#�JAo�������1va���Rpxi�r��������uL� �?������Ŀ<C�Z#ӛ2��I�o�gv>�*�1��k�F;�|>����l"��y�q�+��~�ی��zL����q�I�`�\n��TԿ�Y�)��~\i��I���;��Ӳ�����-|tǎ`x嵔�F��r�D�B����@,��j�cP��%2�d:����}úFB,���������W_��Q�u]B�2��}�"��k�p�7�~aj�rG	�#{�����J� ��8��^rm"Q�x\����5�()���t҂s�^�X*�����	7�NK^��(��D��՗���`�GQ�J�"f[2^�(8)�� �ؑh�����fW��J����4-���p�gR~�1�qZ��v-�Mu��0�a���cءx	��¬�Y!��v����>�j��+x.��b��ط���8"��H�����R�M�-�'�%yL�(�\����{)f!�b�(�.�e��m�U*���@��Hx�}�D����+���]�u���=��cަ5���>4x¾�bړ�X1�� ��F����U8��oj�*�/r���\� ���O���qc !�9釵�Acx^^#|�T ���z>���amR���`��j��;v�?�l��.��A&J�wԂc����}�~\�p-5�v�ߘ��	�ꁻQ�6�0����_*�����o�P[j��h��ڿ�gB[	���Y�ޑ|������ߠ8���i�)�M�h��ȣ,${���'1�f5��22��:[�����aDEh�dT�l~��F�`���oNjvD��r��VЗ9�7`e`
t�(3��Μb�ݭ���ޘ%�09;�� aqx�P��u-+Ck#G�K��}f+����?���x`?E��3��D��1;v��s�n;R�0'��Uې]�zs��lF?���S�(�d�\?��O��6V���wXo^'���
m �L���V){�z䗉PҧC�o)�nq3=\EI_��uT��uj�@.o�d��%�0-��\�ky�)�o��O�/�����2R�Y�����Ǎ��=�������[����ɾ@�n��"^;	���(���̆��P�a�)3��>*���a�D�˥�-��(0��Q���lh�E�<!���u�g��b��V6�h�Gpt;Q��9��q���9)������������n6q���-&���d�\��^rN|ur�j-�z�m�\�wPFZ�A\��/8˵�N�}&��b�%���c"`VvM�U/�G��z���XLxR��o�s�% F|b�M>ƨ���/����&����Ck���؆�vI)���o�2vZ+���[hھ͖�G,�#)��	���t,~SO�X�����YFW��V������[ɸ?^TlY$��;���wE�Z�����Ë�ڂ&J�M��o��u���I�T��9�� �F&�R�(��w�t�*O��5�W�x'1ٗ�þ�`��6wԦe�n���[�I~,�/�=5�Y�Y�ޒ�+7�+<p7�(�#\ȧ��m@.���y��#�Ep�_S{}h�k�6�����O��-�R�?� 1F��|���	����A�O_�Z�����P�qB�Wpv��8�悉]Y���K�x�b긯�=	"���NV�F�4'H*Y�����B�_��菜)j��F��Q`%��eI�t�F���¶9�J[�ꤋ������̺q}Z�V͜}Sj��Z��K����N��[<��UI\`����r�8e�.���3�р�V��P!Zy�����hf���~d�~�!Ւ/T�氀3�|�7�f����{�_0P��T��\��p2����&�6�1����&AKSj0?V�/M��l6��&��e�po-p��1��%���i`�>���:���D�q�]�q���[6��\�T��A�;�r�����,v�J��/tG��?Zf4��^O��᠊�����Ϋ��3G�`*�/2�g��|�y^Q���:>/�HGe��H��Ű L�YȄT��2v����kqo#����.�	,D��9	X�{V�
�~� ��Ο�PӋ0+������9]o�k�6�������\�l�\,���X��3��g;�t��)������瀑c\��G���}>g�C5Z��YM" \�7Yw��k�����^���fڎ���ƙ$7/�Q��U��8�=f��U��1�J{]J�]�u��1L��O�dp$ID�ޢ��䧰��CA�zSAJ�D-.�جCg���e�f^�	մ��$b�:i}�<�4}CoQn���'ތdѱ*<OT��7�$ �B.���/��)���?�S��9�����Us�bD��'Y$��n/�Ӻ�Vim#)3H*_�l�\T�;��M0�/��B��Y��d��р:q~�#0�%�kAQ��_ l!Ԝ(�$��N
`�V�k�֑��W$�����HC�^_G�>�{|���[uGBq�G]gA8�&��Q���y�}�֝n`�)9Km��7'�Z��;k�s[-���1�
	ϼ��*;���n^^Xu{�3z�d&r��}�G^F��b�E���x�mW՝����<�f{���N��+����mה�F��itO�F�;�ns7+������a�n�ւ�l�#�&;�.��P��^j�ja!�j<�ݧ�8S=����z��:�-o�aB�d38�9�4��6�+�\g>�H�i��N�4�OB��Bwm-rZŨ� �*d�7���:�X�5M5��7>h���<�Q8��V�ᤛ5?F�X!��ں�;��Bn֭�@��Ѵ.L���IQ3\L��d2N:�Ћ��<�5i<N�W��k�Y]�xvM	5�n��(�Q�+<Z �@�v衆����*���a�4c�x���+�j$�O�t�P#-���u�n���S���&�
vǚ�5 ��چ0�'���#l%�Ghۧ�;�,?���s�z�U)7�ĉ\��I��Ug���M�B����2����W�x1� �)�ސv�smww{���i�}I�*L�}��]�3a��^���b���XYu��"��Zcx�`~+�$��\�*66�m�����\��!
���O}Lx>E�^D��>�r ���TF۵I��ߴA�#e�o[����R�(�V�	�F����Fz���g���ɕ�ԑۘ[A	ŭu�q�][�Ο�ѫ�B��M	�/�H����|�	%����8��hW]|0���!���1�w��
Q5
>��2�8�0���s���w��X��}�xN���W�#f���׺�lOG&����G�������8L!�#7|�����լ����Gˬ����u칹tr9�|�Jħ�J��4��?�ܣ{,�{ڤ4����E�P��l&�}o�e����1,>l)�&�oN��&3�c11Z��F�����09E�8؜��i3 *���Y/~A��C����%}DD���*�췞�
�����z݆ŏ�9��]ܮx' "�'�A�	n�#�|���<������-��-���2ܰ�m&#�<��_O<��in�8v�':��ۍ����X�~l�����[%���n�T7Щ=�{��
�����^�+�T�T�N!�؋����;����o�weK+��X6v2Q� ހ[kq���b$�Ee�H?N�0:��]����rp	H��ƴ��3ΉE��U��u���vm��zx��Q���S�8Z�l�En����� v��f�����y���R9��w:YV��VU	G�D���f\�XPX��	���S�%3�b|Ϗ\�1'F�8�Ti�����{׿��}�u6��=�V�K,}�?-�l�8��p�{��.�є���"	��$h����'��On����C���c�:t:t7S�����oVf�*�:�? 5��7ͫF��X')�������X�(�(=�[V�X�6R���I5潗���Q�d��*�	�w�jS�̒6*V}뀺e�2h��:�F�66���Z���a~���Ǯ��~���W�Z!��&���Bˆ.���H(�����h-u�k4Cu+�|]	Ia�����kA�T�\����*�f�p�`!����� ���Tn���<��WHSPп;^���|K�+����W�ߝ����� \A��;/Ҭ��󽬔w�o�(#��S�UE3�'��P~d�g�1��a>T��/,��Tdk�C`2℈
sA}n�t?䱲d�8��Q	E
$���`x�΢@�f��eMYB����Nh!����`�6�ꮾ�1�Ud� J�������3�뇷BA�4l���>�Y)������H���G��$5ʽ�)�)���V:���O�r�&��J+ �(�z�K��A!���`����8b^��Μ���3sR}�M���Y������?5���ٮ�(�"[H<L���Iw�$�eD܏�77K���e�,��Z̸$�2or�����A/b`	\��֖��;�������ͻ���95Z:r)"�_>$�X��b0:j�M�o��7x���5������
7�s�TM��^
���[!������q:�]'���xc̜N��w�u��;�V�s-�M-N	�!Rc+2Tm%0������̽��;10`p8m�5��/Rl�uO�7�CЊ6�z"8��U��"�n�h�����Ϡ�^0PT"�(B��@�P9��s����R����5�B�3����M��R8S��72d�XV��_w�6b�o4�<%sҁ�cs����'E/7�.#u��V>"6ʼ���pM}�T�w�5���ފc��%U$P=���E7ы͌(�d��}3���D����:lO ���mdZ����Z���T�B�('0�,�^�`�2��K�*Ź�A?�����M������\ �hG��4A�l���lZW�!ui��U2�(�b<ŀ\r���,�>ύM;���C�u��B��yogi����'B�=��x��ZG�1h�����o����q#w��ߕ���9�1K)���;	N�`Z>s<!��)4����$���N,�������Р��[5 ��'�������Tj�o0�t0lk�3��ܔs�$"���#
XD�����S�~A�e$6�A ����6����y6n�n�W8�2�Qu�,a7�j7�f�>�[([O�O@���<�I�f��&p����[!!����R���V�tI�g��P��y} �sy�o����g��V� �Ȧ��i?f�(f�S�1���p�Zs��+H�O��~�{[E���ͯ�Tz��$���k��~Y;L�%��v�8ȵ�c�@�\AЀ$
�%�6vv]~T�,�����}����S��������T�%��kf��=b c�(�)�)��V@D��Ϟh�܍ ������ ��m��d'\��u�^_�0	��_HY���ZnH���@*���0Y��xX�d �����j�q���?.��Ph��?ߞ�A���lې�4tJ�u� ���E	������K���U%X�n���5Kc���`A�_P�-E^�R�Z ���N��U���_��LH/�2:��d��5��덇:7�*w�_}^l鴺8-j��
坮��j"�e����Z_WbE��MD�Ah��w�.	���ࡊQ5+F`��j���5��Ʃ�R�v1�=8%���L �TK�Ctݠ(V+T����P��
�o�5����J����c))k?׼UA F��J!��3jL�C����Jr���Hm�&S6$/�^�ł�m"�}�K񾝢��_�:��Κ,Р�����Ay�r:����U���Iפ����$w��}�˩���a�'U�_H�`�f"9d\���k�E����x5��y�Ӷ�E�tv4騲��������j�\S��Ho���ϑ�s{�������A5��2�$����G��-��p%r{�ӡZ��������)����`�����=�|���a!�����>9�<I{��sTZ����-�U�5�M��JA�����߽�Ё�Q�1�WG�5#R�	�j�n,V]��u_ս�U��}ᙤ��.�{^q�s��:I?�Y���K��/_E"�E���b�܇��VW��Q�OU�*:R�4൩T��p�2gC1�~׼�0�/4�e��=�C�3�l���w,�M�
�~���)Ô�Xݙ�T��SV���p 徛�_S�϶3�n�l�I-���M@�9V8g���C�	��xj���j�@��Gt�`b�
���(�F���_T+��qu�B:�6=�����[��U�_bk7������C=;a��a�b�]U����E�1k��c�x����*甖��9gH�+ǎ�jc��]�?+�e�S���(]��-bkhP�f����k��p�6M��4�S�Fe:�p��m'L�e�W4�Y�9�����[�ذ��Xj�IH��ۈx��eaas
1s6z�n� �9�(%G���۰"�����o�y�6����`�TdWuok�e� !�w���6 t���3��o�3��&-�M���?��Q�4ޥ~��$差����k��p�>678�'�p��^�����\q�;��{��B��d덣7���)a{��s��1_׉U=G��.��0^Hh�,�o��k�����` F:q����3%s�o5n���w )�$�}�o$�]�Q��.D��_o�'Q3�Λ�-E ��2�l���T��s�66��4�_�q)Ex��g�r�k!`qT]q�xo�=�򌈫��`"O�kf�X�hf��-�f�q�A� ����Y�6T����F-�}�����p�_�H��k�;�6mn��i~�.�H`:����FʎO+��A��z>7��WX:����8�_8��.�fQ
�����uN}���#3Չ���֬�n6⣓@s2���ԡ�1.]ܗ��Sa�s�����P���S݄�	�O{`]�]���O�T�z���m�P�WW��&9Rl�m�-A�m�榓s�Ev5Y�n:���� F�d�����3�y{k��O���5.9�pT����b�FQ,	�*�P�/}������=�w���ˉ�_,����~*s����<Yq��W�-�⸏�ܚ�Щv2��.��i�6#��~��L�d۽��'$�\9��[ͳ&,�$`vK��ʩ��V�������^w�1;��Ԯ]h�'s�F���'�2�+
��k
�й@ths�c�t/G�(]"/=�fM�s�di��_7���!�F���N4vyK� +�#�w*a%~%�:3���\ڛ �U��}�q���^{�\��bq�~ڹ>sI9�b�}��n'��Osj�
��;gV�H[�Huɺt�7vҴ�5�l������r����_�ڸ�7��*k��
Ȁ���@U �I,
���(>>���&F�̈́�/���Wc�a��wn-�Ugd�>O�p����g0q�^�NW"w�q�ontMw[�Q/u�����pe��-��07��aW"U��Dۙ� �i�3��j��0�I."Z?{���� �qލ������>fx3nj�5�r�t��~J [�	/��H���%�G�ӊ6�� 8m���\g���
�G&�����l��4m꾭9����`_z,����X��S��ӧ&Ҁu]�NvD����gDK��#K�w���K��"6�����G3t��Or�Ej�^�xXig��&{>G����N�nZ/jl"�H���!�\��r��M��&�$��3\_�M v4nȚ��%�
Ve���<N�P�$KN=���F7E�w�<�g��鶯�7m�k�_��J�u�L�ׇ�E�wZ�3�:��m�۱[e�F"Ve0�*/�=�����ĊC6�M�Jxf�����ZLy]1��:8�O�<��\�~hi@k�a�z�L`WĒ^(Y��a��po*Pz0]��/�"���C��vhb+�ۤ��"��Ss�ǻ��V����ӎ����H��i�5ƤE���^��'�}���1�����m�^��	�'��A�0'P�ʗlX:�Wdh[pF�[���s�֥�.��a�i/��� :t��f�4�"}�H���q��nRzИTa,@��Bl�b��V\��t⟿)m.B�V4��h�a��vPr�䕫�&��v��4�q��m�m~Aė�颕��x<�y��+�</�(ߜ�<'��ì�������:�Q�Ĵ�`/dn\��fP_d�7v�YD����
q���^�Q4f����m���>����A�b���ZK�Gme�K�/^�P��H� ��o��\%j12�!�A�W��a���6P4��{��N�߇�$�����C���� �,�Љ�8�3�{cu��cN�؂�Ю������T���3�P絠hRPc�n"�L���f$jO�+6 `*��{-?��y7�O�ܟ�a5:[5Vh0mq����H���ߵzSy���!�1j����G��
 �n��M5�\w�ԤmǢˠC�v�d�[ ���%ms)�R�c[I�����[k_�iH��￻��� �^����|�q�@�����f�L�<%�;�,ٜ�Z=t�h���)��t���!��fF��7�'��087������6�h���a�KRh��<����y�?#�2�@eF��+K��m�

�G9�+a�mY0��&|��]7�[)��.��㯻�*��X�FLȱ^�v1�bv�.�o�@�U�^Ǆ�$g��ʊ����{H��������L�󯬟�.Y�{2'Õ
Ag�> 9�c����)�w��$��l}f�IVe�s���2��a#��tYT˃Q#O��IS��%C�鶇Yԓ�s�p�F�}h70#��x@�R���꭯�a0g2/�+1X�
>�y>��X�%���@��d�@d�Q��*[2@e$Ɉ������HX�Y~n��`�{A��@ҾC�H�-�@�*��;���ʎs��Pd�6��%�W4�x��4?qe�o�U�oͶ�3W��`�l�Hr���YW-�f��S���E���/� -�o@(�iAג)S�B�Hc���s��Z_r�4�l�!�=R^�>�4��@�����a;S!<�|����;����`&�:ԭWȃ3�;)�)bMX`�t-T���l��Zv�%��j�XKN��=��h(a��\m@!�5�Q��s%�i٘�Cᇮ�J�%5�k�S���-p{dBlm�*�/K��G)[�vO�v�r����g%�R*�Ҩ����!D��<CyHebd	:#A(n�"�i���_;�ý�l�
,b�s��X&o�<�^�$l�	�6��T~~�z$���g�㕦6��i�X7z�0�1*XU-A2�k�F�)�@a��y&&h?G���)�w�#�s_�Z�EHTyp_�T4%�g9۲������X�q�F2�O�O)>>h����0�6f�C+_C�oO%X,�+��d��яG�x���(�5�4m��d��iZ d���y��?�[�����u�9p����֤�|X��y�K,��bpjD1�����>�4��TlR�\6ğ�sӽ������s W-�2H7⹬����].�	�<����������M��x�|��}ta���~�ާnn����%�����Y��1�,�Y�뗦�59>��Nn���"���8�I~�λ�In5��y�r�"����M�J���~Dq�֥�zg�f��'����+�&��"Me��Mo�a֠�_ylզw��]��3���D���i�Pپ۳����3D��t�Qּ3e ����k��.�_��>��9M������w���Xݲf�' ��]��2���xt�uzI!c
�/�N	\dݷ|�Ž������P��k�f�û�w]��(�ީh �V��X�1Qb�:�'߳2��Yh/"ڷ�����*Кo�7y@K1�b�&Et֤E�O&����T�>�� �DM����P�6� ����j�YKG�4P��$ǯ�i��@|������2�ܹ�a�W���YV�3��BZc}#m����@���ˑ�Lst�-z�>�鮇�����ߥh���.%��&�1��L��z=�Ȗn)p��ɚ(�.��)���k���S�$x`�q&r��,lnW�RC��|m��e
����W�~��UP��\9]� 娺�;���R.~�)(m&�S{�� �q����gEl4l�>��
\�P�񈞍JmZ���s�)4_����GI���2��ʱ��>Fo�1ف�(a#V�K	�׹�I��db�I�c�G�����>��c8v]t�<�<z��.���r�(�$����� �7��+�~J�$Y�8�V�1SZW�����fdj�٦��$���z�c�W)��F�BȖ�~9��HO� �o�3X�9�����n�]oR�չ�pt�� �+XDk�L�3�rr��"I܂���i�:����s�/�_�
��q���E�.�Zt��g,i�K#��T�x����>J1P��E~�*=ɝ>��v��~l_=zҚ��T�pAv&���c6�����@���a�"�5��D8k��p��D����T���(��b2��Aު��1��[���m�s[O�����`�)D�!�=y,}Ķ���.�� 
HcV���p�v(z�Z��pT���e���xuHʪ�������2E��:�lq��O��8ś����su��(�i�s�;��<l�5���9��������i�"p�}S�}I��Yđ�_����}�!N�,�D�n���X/��Q�W�v?_���/�/�rD��l���]�R}tP0}1d*�����#��'��3��/��rI�� mV�s��g"0�`,��	��R-�gQt�lc�����a�zZ��2�}�YI�&i��~�\n�z�|T�:J�G&_:iS�+�����(gT��C�"�E ��5{�E����y�U��q�.r]�R��0٠7�@O'W�	s%��,Y��	O��w��a'�3 �MJ^(�9�C�'�(c5��x[O��f�?'�d��HFv�ݗ+Nu���;�W��}���̄�������;����~Ò!���D�W�A�O���U'')t]��-�,�f�T}����Y���{�@~l8'ms\�������gW��8�fx$ov��gm���g;�Ӳ��,W�G%�c�}^%T�zw��`wທMo@�q���5-�� eĮT3R��Ū	ȟ���G7��Z|U
�hQ[l(O@u+��Wj�D]{,!�G}S9ϩ�~`b�x�R�k1�(c��re�j͕-���]�׉,�릠��D.��s���ȍ�w���Pz�ƉǙ��g��l ��y{�X~�H�~PI(uf�7���p�w��r����4�<��up��PV�8~+�I��r�4�|D�
�z������v=��y�a�4�1y�b���B�0pt�����pP$?�����z?��M��A&��eR6�s�T]��k�V�Hj{M�r�xή�����Wj�/6ҐbQ&�C1�ڐ�3��a	P�:�1�>��jE��*{��XlÒ_o裭�iD�%w7pU3��RY@l��?S�g�OϚj�x�x�_)p0���R�ۊ�^}�뾻����ٸ�P�#>��"��2�댽�������X��[�02�D\Ln�����+��t3�[5�I%�K ���uض]c�j�!���s���X��
�� �)L#�%&���4k:l�Z�MzOͨxHX��;3�%FގyK��k��$�0&�.8��<�@�L�1�r��`�[�pΤ�{��{&�\��+x���)��|)��:\�
s�ƌɿ,��#7��=�Ёy���#��sG�6W�g��:�|�H������t̀iǉN�.a@�sC��]7����c�>`�_��bW�d�[d���3Sϝd)��I��5 �2�Qά �U���cj��Yoy�3[)��0%�
��0)⠏X��T�σ~��EF��`���ߪ��G��S�����:f�D��Ip'������Z���4��(�9+����o�O�f��?���r�^��S���@�sP+P�Y Տ��dK�Kb����Qix�a��
��.JY���JX���`��V�ōH�o�k���p��mь���K�W������u��Fb��K���P�)t����N�+F��E�����d�6�&@Zh�pO(	,���D����Y1_5��'����̪�dפ�A�m�:M�9�R~`yޫ�Q�{6ܻ�?6�s����!��:�l\1w��c��pͥ��~��V��a�Ö���Y��(���/�`y0���/ {�p~�Np���o�~7`�"_3�3�F��b�����"��r�D���]��W�)��і��ƍ�g��Y�KT�؋K�Ϡ})�4���:!�Ru2�c���kU�
g�nu�ˊ�[m���)�vcJk�$_�
}�����x�-���>�D���F��Pʦ�C)ڿ�M�e�yE�x��H�for"���"]��N�r̅Q�Ko`A��J��G�頟p��b߉dy C���;sl�o&��AF��n���C��b�!����>�ɧ'ۆ�v�!/�=��)�>��$����%,t�斣T����C��9����EצiH�:�����J�ꖡ_�/��� �� D���T�MA�� ���|e�)��z?���\د�b&��N��vJ+Zi��PS<Ӊ!˞V,4���(d�g�rv��_�A�;��O��W#��7ܹ���l�s��!���<G�iH��u#f���-X���^0 F���t�i�z<��o��j��z�KpSS>�>jI�z���dß��<�/��gٗ��ٕ�~�.a�ȕ_d�c)�D�c��!��Ra��	VtA��%���|�,��.R�7X)����%����u��ڤ`��U�C˕TU+�����Z�u̻����IC1�>=7�RZ�y� C�a ���J
�f:�"�rzs��9(w�����)3��<�x`O�&Q��
�����9զ�Y=�D�7']))�V���g�^�2k�����I3�C�~�θau��K��/d�Q�1(��V��OET�cyi�QO5D{Ƅu�_(8{N{��
?j��l%�F�#ʆ��c-(�
� 6�J\��tx���HR��u�	�=.�:C���� ��n�O�8��9�g]')��[���Ԕ*F�X�dq�;�ƌ�--?Ԡ�	�.�Z��eϰk�c�_���Ijfϯ���5ǯ��S������\�H�v�TSʳxov;d ���Qe|в���X��V�ר��<�$!C|��f?���m���.&�,	�$1!fc?�\��[	��6�TQS�4�l���gQ������B@<|��:�ѱ蝕q|�9���c0���R�sFpL�wJH�x'|��'��f�e�2;�K�pJq]�l����$X������kS@���Uq�`�нS��ņ��cm�[-U��v��ڵ\c\=����2Hh��4�#̴|^�i�C���#����;m<<~�X�츸Ve�ŕ�P>79�����BA!��-�/t'����M��MW}X�z�>�\2�'�����Y�}�)��~$V��AIQ�1lz�h,̴�^��!XY�R��������H�t����O�M�C��� �`gJs����͑�!ͦQv;�j����-Ë
�q4�{1�I����cvv�Z��N��/PpXSO"�6�ܧ��Úy:�jߕ�z�<��Ï�mX��MP�.}-4����x@z�m���o�'@�m�a[a*�u1�aq��k�2[-�����	��Cse��|����O�iۊ��F�uA��1�C·�:��
!� ���6��y��"����g��	�u�ȶ���cp�6gw��ǿG?fj#s,t�?ђ��(�?_�h�� ӺJ�h�Y֪�.q� �E�3
Q	j�|?��Eb�8Vi"V(��b@ۥ�)���-be��_v(�*�������ww�uh�o�z�tn���N�Ev��3����Ԥ�U�U�9(9���$3�<BV����lj��+܌�P[b��PK��뀂��8��I�x�n��{�̯+�&W`n�%淀u��&���@�p<�7O"e*��Q�""u���!�s.=g�6L1W�PF�W^FD�)ȶ���`��^h#ls���c_�w��֧��ҕ$c�T��E���$�S�{���<f�{;α���AP��x��ߍ�"k�ٽs�#����bZ׋���8V���ߦ���&��+��Kh�urhP�d�w�X�ѐ�+v��k�X>)�ɊEc�C!����[�CE���ncF�-���	K�e�Q���w_>2�wp��)Wǆ0�kW��Ե3�5�R��9�|�.�f�b��g�U�4���V���(yf�&ls��M;L]'[A}�Rx�����>#� �[�{@C�Uf` Q��̮,�� 8�=ju�d�ȧ�]B$�#GĢ]�������Sw@�5R]�RyS�n�x�,���9�3QxsE�~ί����Ucemj���o�h
�&�0j�o�!�&Fʾ����N�I�dk�<�A	�m�b���^^��'��B�pH��c���ަ|0�K9��T���HC8z<l'T_�;�n��袊��x�����۞��.N��h������G�BBJ#�q��s�Z�_N��?2����	&�_�����@8T7����%Oqb�<{�f�x4:�(�'�w�5f~Nl�Q����AP��Mi��jHB�l�b�h�6�pj�}"�A��$���/�ax���/@������[ΎU���F�)�&F��_[2�$cTD��z�����d,��/v�pO<�P�����#�pk1H@�X���_���ŉ�i�>�W��_Yn4��Ӭ�P���VS^�`';OYK�4-���U��Y.�9F�Ķ��Ya���3_�4�7z�e [C�kM^/�g�V��$�O��hDΛ��,�8b9.��쫂��n'�����R5� �zMlY��@�/�?l�f��8E����T{���;���PHE�Ś���Q��U�Ձ�un�Tu����W��r��6�Ƶ���v���&d��U����OC��X�K���aa���l.��{f-|	*�\�ߒ����.����l���M�~NF�t��$<�@�ev�n���4Zʹ��Y��Ej��{`�vºX�0�@|�G@�&��(�'���#������Z����`6_�kzŖ�J�I��	�z�@�B�h���1����@�2t��@��R_��h-g&��W��dנc��3��FOp�f�d}�S��ek�\I@��G2���ঽ�2]3sA���̱�v���ЃH�`_�%�[���K�Ow�VY"a��Zhl[f	��iQX/^MwU��`�(k6��u�ɯHd�T!b�y7wFIn�%��YP�J$�	�x-�������Ζ�W���=�UDX�w�;����p<%g�V,m��'6��J׊LO�\��S4��g�hW�%��-�߆�qGVI�o���)j�9�v�+�B��崷�ebG�#|ƀ:��GΛ;��B�6�e*T5��D~��u���'��O��nB�� ��4�o��ӽ�v�!��3�WNO{!dL �a�\ڄC�D҈ W�!��'җ�U}��_�I!��9Vq�Z�ӁF�.d	.�c��_&�o�:݇��X�M����D�]��sl�u���KvS��YwP_�˵g�m�;�#�،�j���\�*JX��f�tC�7�zT�f��	s���П�όM���G�9�N�B3�mğd��$1��d�A�&��śگ}��{�/t؝K`�X�3-��Gyr��9/��l)>nD��ܔ�!_�R�j���g��?�F窟ԱD�����IW��Gʢ��?ĝ�e�{�������������'0���4����4�$�[��#܀ڟ���5�/�rv����k�X:�j@3�g���m���Òw����s��*ų
xb4�,h�?d�3[�w�vNL'r�����=�BI��?��-*���]��^�U0�>R�dv�O��`�f*^	)�O�� �a[_���u?�,�{l�8#�w���r�tw����b�e����K�
Qn�b���&�d_n�Z����U��D~�ۏ���\�,�Z��ef7��v�3�mՁ�U�B���Ɣ�큂�hC׌�'��h[��17"�U��*�I'�d#���a�s\XIiT�����R��Ʀh�Pɣ �C~V8�j��3��Z`�%[���߹�r��:ej^O<�|"X���(�������'�j��`�i�����H��/g���x�	�*z�!e	b��$��y�Y8B��vR*dt��7U<�������ibc4>�t^�*��hd��0�1�G�=1O��X���:矕��	8 ���I���]�e!�2:���?�3N�=��h���K:1@�P�
��H��)��z��H��H��:���ɘ4�>^��Mj�;��u��h܏�@ 1k�d����Q�Kp�A×nM��%YF�o
J�lV��b]<]����k7�7Ǫ��-D`�[^���i�Y|,�S��4j_y��e�JM�mS�Y�W�ly����;���ZSժ̎�T�Hq� 1п'nf�c-�<�-���D��;���i�n �2�N�T>����w��3�_T���P"���XE��m��9R.ف#��8n�_���š���y��l.���'�F�hq�L5Ai�~;����8�?I������XG�b���M���k�W��t�Z��k���^s�h��ꕉf:�)6�����<�#'1���ftב��N22p����,(�:�Z�o��~��=	Ɛu+/]�}W���N ���ψ��@O�m��������c�"�@;]�_Շy�����T��7�Th�'gZ���
u���:�l�W�Y?���v�N6[DՈ�_�0�Q�����~L�|m��Vt�,8.c0$4t�y&#�25���-�#��4uC�Bl�=C�"��^����2���]�ڨ��_9��_x�Awo���ZX�a���а�j#�'}�})����.�|{v�$�mB撻�>�4^zX$B�z�2a򭙆�;c�>��&1���m�i���9���Ia9}}�J[��/9�ث�W 0�1Pmx#n�W����=��ġY8o�ꫛIξ�7.�U{'�҈O
���Ǯ)�t�Z�����S�B�(��z�sDOdp�}\0f27��YJj�ڌ`Ĺ�m��GE%"��0uK{�F)�
�g��般��� ���&ݮ� ���Z7�ޢ�%�:�7���5N[�n��a|`K��0��.������}]/����}�����^���7@�%e�;���X�MDv+��'
y_�@?���@�m/�9z��/��0�ܩ@jݮ��	y��x���:��7'S��?�\"�H� �o����8�㝽Lr�_`��*Z}��pp�L��=�ݪ�ı5�X256��b�ϢX� ���4�h���}�Hz�'�^���H������ޱȴ3D052���sA�N���P��QQ!�i����R�0z�*��'���a��hC%*+��s�C|���"d(���+��ă��Y7�~8b�E�M(smD�$���c�Ę�x��M������6����Y�>AyV�Rk����d7�?<�b�ڑ�L���ב2Q-�s���Ǒ��8��.�gڭ�oݩ}���:��O��4��H��R��O86G�i�u$޲�p��Uuփw Ej����n���:l#���vs��!�8���:g�:InԿ�� ���z�%��`��:q�ͼO4^8ZkF.:��I�2|�0�0��Z ��\��l�|��O.@�n�����R�Σz&��g��`���2���?�u�r�&���Ym�S
v�,"7��^G�a]�u��0gӉ	%}h��W���S�UCV�U�ģ���$PD�%Y˽�-����<��^�+�����ɇ���K�м�槥FOUe�2��J��1?��|�_x���\?�v�I��(O6Ll��\Gb�|����@,����Oh��^�G`e����ѳ�$���=���+̺��1&���ܻŖ������wO�c�P�(��1�"#�*)�3H�Y�ό�����f�"[6����JK��w��g�.�"{7�im�K��s,���Jm�*C��F�i�Iw�L��+5�e^I� b5�}"M:9r����0UT�����]Ԧ6�6��b�/�W��ʴ+y��j���4�,��|4���0�HHL��,3������Ł�@e��a��O_��-̽:�T�+s�
��Hu���>Ϳy�ۊ�w�}9V3F���G����[2�x�j�غ������U�0!��J��^���v΀������ c�>�ak'��C�������n��e�JB.�f�s���f�ȑU�1�T�H)�E��C{-���R��sG�K�^Ôo9�^��F��#����Q�W�YdI�Bxs,P��|>��y"���8á��7Cߖr���?O3�mHM�+\�
�Y��ѧ�]7�tM���  }�/4G��,rs��,X.Ur�e�n\���h*�JI��yt�X-	8��j�����wX���ބ��Ŀi�KdS����ΐ�NH�6
q=w���"�����^%�T��F��SI���g	�b��񆍹�����|� nه��"�J�M 	[u#��-��}s
�
`ћ�E��cv�r[�U|��՛~-82��@:K�+hS����Y�ڝ:�sėX�Mbt"C���Y�:C��c����lv��j�)� 5��Cu���xҭ~r�J�֍�Ka�3Y��9u���< �< ��V��j��x��9RA�4c4�֟JƧim��ᔟ͓pl.\9*�`��X$��5��J||�OQx��EN3������	i��I��S��`�A��OA����S��竐
<���&�G�&��u ��\[h��B�UvO��n��m+�"�˼�Q�Ö�N9*/1���.���5䨋h$K�D����g���Tg'R2.]PkE$�#L4H�����Q5K���~���0�o~Kp��&�=܋��e��1O=�{/���D��0Q�[�3�E�i�d���'���4�Юn*\n���zL�nW�Y������Ա��������.T�V�"�Ko��r�,��L��L  �+\];㋳[�W/�[<W�Y,	�{K�x�Mw���d �])�����
�@t,�-����ʯ�H����F��/�� s�OClk\�����%��j9sv��.�h�hKv�������rp���p�Yj�4!��t���wȕ��uG�c�����^�$ek[�����P�t��M=��۲�7b���Y�m!�-��Ab��m���gҰS숀��"�Y{��.39{�e����^�z�<��	5X����&���;����H��a��P��t�笄���V��"�$#�%�:�B��"TҎTWf�3��>�%�b�Q��6�۫>��N��R�֜E���Kv[�c	j��H-�N��(#v	Q%D�9�k��H��[U��1�S�E�hI��~��-E��'~~�	��&�"�������1:�h>�#׌�Nbk�&�w�� 9	G�I^s��My�w�3�4~���Ç����mΰ8$��S��#N~!6�[�(���
\�>��xӭ�ߑ���z/�<J���כ���(do���Şt������BL��'����V�l��߼J��|608�!�G�"�Y����A��V{��&�C���W�QX�(Oe������%qQ�w�+�~@�etK�>�ڛzL���O���[�`����N9�P�������텹Z,����֥�cL$���MPi���P���H0�\����QT�q~��KH�%�ˈ�:������°�-}O��`���ӚQ�.�� �؇
��Ԓ�� ^)�(�+c�$e|l�L^��u��GI��ݦ@��Dt=�=`�����(�	o'"�sʳn0c��p1���_K{N��oQ���râ6P�R�ω���%�9��Xp����Q�wb3�p�dZ+T��+�:E�8\����k,+�ʉ�
Z���JE�6;��-i|๎�m�R���`h&!���A�cdL����W@j`抡Lm֤J>xnpb�3T��� �2�X@(���������FZ���^*�[$�%,���uw��!���,qi(*�l�Đ�o=j��,���$K3�\L����Y�h.��R�>���� ��i\D�h�P`��:'o�	@��Wzv���݄$V-�a�u��F�T�1OĊ��B�v�u�Fe���6�E��d��kh&�g�6USnD��~���{�`D����B��"��� ���H��VĜ��6�� 6�d�Ⱥg���Q����V�	�:!�6v"m)1]}�46i�$d�������Ke'��O��M t̖Q��������H�$$؆ϲ?h��A��XU�аe 	�8qi�^��E�\�f��!�,�!m�Ͱ�2J� 4˩5{�]N��8$r��lw�z8_Lr�H�������8m����R�M�F��o��w	-W�;)���g?&��Yie������	��2��H,� ٥8F���d��%��g[���]�!�64>�4gQEUԩJߧu	_ԥz��L�'��ц��1�o���uIXn�r������&�ʛX`ӯ%P�����Z�>*�.�s��Oz'�T��v6��B�gK$�Zb�&O/���a�f�u����?	�$CSӦ���-Y��^�b�5��Pu�LyKE�׶>��O�ȑ���c�Ş�/����Yh		�i�Gq�,�/`]iRv��f`(d�.�R��aX3)�^�nU H$�ڢs6/���������oJ�hʌH3�4�-�%&�����}���Ay.V�Db��T�����֠�*���Հ���#\2�����O}h�|Qths+����T8)�Ph�l�Xbj�c'��o���4s�u�����剫lj�g��,��Wi�v�]ƺA7���с��3�dڅw&k�Jv��k#���Ha��O����e[�����TE���
���7�%�=t$r�|������nz�G��O_�o�/2n�)F���G��>�=_�����e@�]J�dȵ�R=��!>�d���V]b�^�B�	gX��0}������SP/֢�;�]�֡��t��9w�c�eX��t�Z@$�`��|�
�qs����M��U�׿6	�YYPn)"Tf	<lC]�~
X �3�/aaq{��R��G�jp�{<.�Y�r�戴�����Az��Xy�_���Q���\m׊���9�b%`��Fa�f�	�S�-ߨ��P$K0	��� �H>k�#Mfˉ���s.��t!`�_(<v�=��`4،�C����S���a���B�R/���;�#�9�S{����ʚ��`�S��MI��/�+�d�+=��� 9�E3泞{�6 �-mk�u��Ox����<9��v�i�1���Z�.�����6�ṥ���$�>\]�;�ii�Hyf���8l����d�Y��+�m���^�����W9}�%�f�7���>�����!݆j�R��3D=���4!�?�5��*���-Y�����}A�S���
�R&m�m2��Q)�r�=J���{��a>�t�	5�k��59P�~�F~�~�;9��}ݚ�b�.@�+,g/#hF���x���+�=���M�������E��40b�W#�hʊ�cMf�A圻2/+���m�
�ȼʃ�5*�q�OX�)�L=z$�gR+�@W=$HE�L��?�c�b��d��2�V�M������7�2�����cm�(�US��w�V�qM�1u����	�8Y<Lne��G�1���fg�����t��mڮ^U;�xA��TD��_�"
k/��~n��v}S��ǟ�������A;Β�4�cah8	Zn�@�a���Ba�^v"~�wF|��$�����V��tj�Q1/�7U7A�5���dT�����	��}�`|�����E��.0�'��:�lTTv���C,$�B�(��Ő��4��i8�&���.
�-�����
5Cb���5�#��6��oS��������&hT��rz�i6��D�����|^�^.=X�΂���Sa�8��?�#��޸� �ճK#�~�6=�bg�=@����2S(��*�����cS�����U	Ε�6f�s̓���������i�<_�<f��#X��;���7�;�����N-�Lg�`At�Wp��>S�ɢC葝�`�K�9���Qy����3�7G@�>��pJk��,��b7;V�ɝ�dZӄ@M�3�A�Ym�^��n�@;����Li�u&Le3ل{��v�w�79���s��xl����`W8�7P�gS�L�e\��B��<2̧�7�#��[N!�CBj.���"�Y0�/�4�D���P���G��^�n[�À��hw�B�^졈�x|d9Ⱥ�I��Ǌ�a�� �7�����ܒϳ�X@������ԩ@]>Ox[[����;���|F�Y*+�iAG]T���=�d��-^+v8���ar-���/ ��N�����/f�b��[O$+�K�Lg�9.��<��'"[�;�miۢ*��yʘ·C@M����(�j�KE/*#�̝F��� ���v
�]:�S��8�,l���E�VJ�ػ��V6"k�g����e��<�>ԫ��k��)խL����9�J��ęH��hN�[<]n&P�\0i��,p���‌��S�n�Y�zsbC݈�]�o[��z�{(_���H���7�T�mbd|'�r��>J1���!��O�V��\�I�g���H?�@?��� �,Җż�6ڛn���^=J'����;袎���n��`fX��S�m1Q	���8ƛ�K�����ǎζ���4�}O� ���B̶��9<�k6
K����| ێ	J�7�P�IC�k"eK�V� �����#��>��L����1�|�㽖��F�.�����|�]���e}����[��z�7�H��N��~)qc�L�,�o1��?�9! &�s}Cgy�+�KDNt�/����]s�p�/n$��)v*Cm��z͚���;�GEfբF�Z�Zf��h�	��a�Jrs���YːQ%�蝆ednӣ�����qL��mRT��$�|�����o��$���jƌk�K�QAr/��E�~�J�0��
8RO35'��Tq���F��K�!9qoY�.���K3oB�~���9/�;�N��NBߪee��x�%1y��c��ac�1�ed}5ϩ�a^�.��b���̻)��$�x2�����Ryd�ܼ@W��l���-�ʲ(l��!nVE�h�;A��r�HdX �;A逩��#*��� r�1�B���,�puA/I�k�?�cAZ&Ϯ��}û������.w|
')Ȗ$LD@�-&�k��(˴\;U���M�t�׼�C4�N�J�0�*�A5�sӔ��
�zٶ�i�yκH�^ZK�5�	`�fT�����6pm�i"�T`�\�ˑ�G�_A`�����13��o���s�V�m1h��3i�kչ��J�$ьor,�sz�~)�g2Ǭ6�ǽ�8wڤ��'��� ����B�:�#W=2���o��7��թ�@(�e�o�)�7�X�(�(� ��<8ص7�M��aBR<c�� ~r\}�
��ִ�e�/�3��B!���BL
.�3���@�q>�}�/gѪ�rh\{��Q��&�f^Kfz�ޭKI����`6�qy�vϾ9{h��걄���pˣNР�yZ��:>�n_��d�8êo�;<��h�s�D+�T��&-�ڨ�G_�)$M��1�,NKp��>K�,:�%/��.��^�r���&���g5�7[I�D�g� ���8���cא� �OM�F���^�-���_��3��&Jh�<-�g�z��3�ί�7��i��P�&͎wA��=��m4��	WLG8�}X}b�0�ĈUE���!T܌����@�]y:LI��[yͧ������X:w��D*������Sx�[�*���!���D��8K�,�X����`��T敢�F}|hiR#��,���w
���>��n~Q��⏐�( ����P�����5����?+.�2�@�N�6nK�(�|�9oǊ�.bۼC`�*T#©Y��c���x�'"SXտn'B���fN�æ�zx��#ޛ}8�Q��Y	�o -�k�0"%��y�y�]Tg5X��iȔ�0�\C��<9�;L���SP�k���8�Ιi��#u�S�e�m��Jd��-�u�S�'�@UT��;�@6 �I�G�Q��կ:���)i�����U��ic�� J,-W,'<e�����D�c����V��':��Cs6���m>��#D@�,�T�T]{��ֆ�����2���x�fF���ؒ>�4��?�&����Lc��XI�8���
�2ρ�M�h�����%۽�������Y{%�)X����;�d��V)>&��=�]�t��������0��+z��=�*�a����E0�P���r-L��*K�ŏt.�Ė=+�J���*�e�]-E|r/�����V��g�w��,dm_e��а�픻"=��=���0i��w`c[;;��s�;�T/&��8��[� �JN#L"�廘p\_I�J1�B0����"`�ju=z&>�Ǻ�e���l7ShyY*@�.$�l��D��i{�<AȄ�d�/�z�gKTwa�v7���t�`la[�IQ��0��-��}͇�ZT�G& ,&H�@��\�9���yĬ���ӬX7�l�H��̷������'�6���y��;k�@�Χ*[p�u�-f������#X2)��w�m)���a��@�4�Noz�'���C�X��0t{�[�Y6�m�s����#睚?p�2�J��AW�)�5�ZI�s,���T��	���o�W�b�L���&�%O����b��\u�	r�o�$$ٴM5n�h�q�R?�t6�rA�o2���6�iH����t�ū�m { ɦl�l@�U{���@��9��e�������PJ�(0�08�[����N���5�M�t}m��*n5��&��q�b&^\��B�y}���<c�Y��]Ӹz���Og��M uL�X)�@��5s��f��V�ykOv�FqK��g��J�q��"4�[Fo��ݔ�v�c�Ǚ�|(7Tn'�}�ǒiq�Ms-�`�n+)��[�A�J�DYA@U�^ަY{'C&N�" 9�=o$�~m�*�*J\�R!Ga8�^T�s��?�m~����l�+��S��K:Hd��*����-M���$�B�ɰ�u�3N�	�G
Q�A=�mT��l:;'`ԉ�B���� L�}_��B�ᚶ,IL�Kx�T���U����e�r1�^A#�T���׎۔���^y�~	������K����(���J��6z��(�W�V�Qu��� g��bs�AA����98Ƞ��t����F��CsM�6�^�2�"��d��u�-K������א��F^�o3�ʉS�%S=�'ۧ��s�SK7�́�Y�s����ߗ 8-\�UM��ewW�f�6d��$�D���Yh�7�1�Q�8-!�$�Zc!w:ٶ�}���XL�����o��n��yP��G+2��".�������@�k�I��x��Z�y3�m媎�>�[w�XĽ���q���Eu��p�ty���H�OR3*O�w���_P�D.���=�_�i=�N�aJ��xk.��क़{Zb���v\��#� 6�~3 Q���H�ͳ'����[guvO��YU��Ʀ��y��*�I��{�Kz4�#���ՇD��x>��Z��m���mb��Is��Y�5�|�!�9)�N��� �"�$��J�ׅN�ϐ�����_�I�p5x��p&a�5�RDLɀ�Au7�K������N[0-;<�e���0m�k�����[W�����5���A�Y��߸z!P��f�A�V g,���o�9��_+l��`����}�N�薽6]��GR�����
/*�쓩�o�{�o��$�G�6�y���V�OA@b@��g��O.���mǸ��M�x$��� |!�M�+����7\�9K�T5�x#S��|��r��GL)}��M�C��ل�����N)G��*nD�4��L�0RE������\��nկ&ѕĀr$:�W$���+1�S�'�љ{"�u2��Ӂ�:�p�e�3���>5���2�NB�W�c�[]�"�r�9*^�T��gÎ'�j�i��Z4�P�H�r6�f��3��4��2J�T���@d�\�c��rz�R��W�����QM�s<p�75A�'��0R(��{��3����!��ޤ=��@%2�y �@�r�a��`5���lj�./��~�Y=܏-�1܋��9�3 �5;�l"nG��z+!%��L5T8��5=�
fH��
D3'��P<��e!������uGѶ��M�+�=1i'h��= �ì�=>Av�Bj�p*,md�ޠ�Uz���s!��$�1A"���nI���]}�#O׫���]n�%%a�
V�=��`5��q�)���?�A	�����[�4�/�%"�������b��B�Dk1-  <W#Z{�VN2Ŧ���'� v�0��қGUr�^�7=~�j��#����//��/�۠��yM��Hl;������.ٗV��ʍ᚞�&l��e�����H��B~�����kF��%?i���'s��%��Ј��EDY�0*%�|���J:,e[#9�����^�^x��Ŷߜ�ɀQ#)Q��h�u��4S��X2W����
�԰���>� ,J^!�?��U!��*�,��Ö�Y�6T'<iz��:!������>wM׋��2��q���Z�!��["3�������-��O�?�R|b(�W7�mɬ��G(�g��`(���[�=�	Y�[�����Be�9�Ks����@ĕ �V���^����9�F/7�fL(�"NkEѝ��-�e��"͖
4�$J�4��g�c�%@>	����z�d��4`��"!�&�?~%������73 ��0���4r>7!��R�:��7�����e��B�a�OJk�P��-C�̜�Ǘ�\	���}�#9vҢ ���I��e{H'�p��#����GK. �S�?er�2��Ͽ��*M���gf�~L;����J���}^[I�2��TE���`(�̍>�����7�;y��.U;{&�h�P���uP��A��9KX�Ii�H���Ƹ�^R�y�r.����, ����l�$l�%T]�#� Ҧ�p~���6�U�$�U�Zɛ���˖�R��#
���:��K\�/p%��x�̱��|�N���Sd\l��5��u	��g�m��]p_���z���@8ﰆ$�B�l�q�4\Y�V��ԟΎ y�s
�f�E�E�8S�T�9\�C+����>5w�<?A� �m�o��f{S��gNf
��(�ӹ�`��,��~�e�$� v��	T)Ɏ_�Bp����R����d�����E�Y� ��a,�
�L�P��P�#f�hY�8F&(ʪ�<ߝ��]9� UZy 7��*BQa��1MJ>OJ"B�qO����:����D�:FP;���h�.��$����F^�@��/���hGH���r���ŠTѰH��È3o(nF��Z1���3���r�Ӡ:T,��Sӝ�A�m�"WF7��z^��Gɕ'9u^ pƂ�L�������X��Ƀ[b��WEB.9E_�{<�'c2�Yc.3e�OՎ�g����4+�"[2�r���ܡn�x�ʯ�\5#�[AA�Ր/�hv�ߙ�9��o���kK�7����0x�T�SҴp��6u���#�j�;��(iv�������m�<l$�}����2�L��z>�m��5,�5�������D~V��4۔E�׌��u���Bu�Ȇ���q�P�C��i���R��#-K3��|���9�}P���Bs?����tY>���F=.�̾j���L,���4+����5� ȣ�+`qs�oUy��3H�/J)D��]
��l�v�b`�0���K��yJ|�� K_��Ν�N�f���}T�8ʿ���[�0��20���GȆ���D�`7���fqB��ҝ�!��Ϲs���Sq�j�ˢ��,�:+�]ZZŪ��P�[��.�K��U�i�Xd�z���3�%)x��3ߠ{��o���N�����جf�И��-��G�e6����b�����B�(mU���y�v�8[�Uծ\����%P�`����ܟ�@�l��mE�Xجͼ�j�Q���{sR@�@ib��`YZ��Krp݋̟���wNƮ�UY3��"y����Z�6�H������Pe9[<V��g,���@� ���NǶBj���V_"3#��{z��]���9T��z��a�n	����x�3oL�ԔZb��#�]�����N�.bo�N��2e�p�JXVP���&Y6��t����޾w��3B�	�u����N�`��2��-'u�<�)�i]��}bA|�<>������[�P�������#�f̇��	޳7��POj��~�;��Yd.�2�o�V�D� ��\�i��PQ�z�[�rHm�$�0��3w����
���Ѡ5#�[�$��}��.�58�����Hov=�N ����q#����nĠD&���:��=ʎ�İ9&�D�b��Xo�~%���7��������|f&�1C#~lO���gڋ����I������R�f<bӫ
:����K_3)�{s�3B�����85]T<.N��zoG�`#���q����,SN�&w��C��Ұ"��QnV1��]�)!���J?�oݡ�*��p�F�E3�;�a���������he���%�ɜU_�x[���r��T�p�67X��"\��;��jx�TO.�٨��5B׻�����e���]�1k�E��&����[��R2�J���u� �*x��o���_g�ǨUC���gS�e�p������� c�5y���VU�������L۶{��d�+�#߆�Q>�_�\�2E٠Ӳ|li��L<q/�8AAG%���i��fsx7t���?�i)�z	��Ц૴�~��,�8<h�Z�<�� ����I����=~�*8
���{"4�Gi.Y���W��)���'�ۚ�L���o�u�*P]����������	�oII8�^���4�f�[O���)�54RR��ѱ�-�	����ؕ
L���漴1%� y�����(lv*j�`*V$��W�����f��[F�c�I��!��m��r���Ǹ�˩�~�%c�5]r(����ӂ����ٟ���'�~q�qS��O��d�<�����-qܞVI�4����=
A0����+������j�N˖ɦ���c�"�=�7�kDX��?���n�p�b��=�uz�F2�"J6������k�TPL�t�R8����I�Z���3W��|"sY�C�"��eqrp�ږmf��|�Z�>BO� ~��i<��J��٠)�|�����X�%6'/��5?����� �Z+}$鼋-��YS��B1��Y� %����ͷ$��˲����H�ld0��HX��a�`���^.���ϟWf|3q�2��!�Δ�ѵ��=��1�c#MG�9�r�^���?/�v��dŴ��te��:�ǔ�*Fӯ�c��(q�9�s�1&\����:�l�x�x���b /����S���`�A�"�i]�>4� z^�q����ɵ8U��h�(Yv��Z|������	���yt���aʚN"%�Yq��Y�o���A����d�nF�"��Ɗ�
:: �mp7m���._W��}�ψ�K�y�:�U ��0�y��:!K�Kh2�MW_Z���a��I�n�UDʾ}���H��͒E��ׯ�[��#�R���B�
�4'���� ���ڞ�,��3��9}�tZ�Đ��H��o���6u�ˣ��X�ܪm��؁�b?�X8�&͐��-�~���>х}/p�Ț�V�pw#��P��N.c�g���PF�B��~��xu����
S"�t��ʱ�_9��b�~
��	���٤'y�,�.|q�
��rS;�6�2�OI�3G���L�~mԴܢW���s���ozۯQ�%���E]�V�߅yD�����Q�&�!�!8�t���^����p�#�� m�6���
�z�2�+�)B;�2�3��F4Ϋ�}�C�9�ϥ�9�
�,U��{χ�9�U�H�O7^W��r��#�a����bK�Wf��.c9�&��9���Uwm���=O�!���I<����{3�D�EΎ��r���:u��5�?/�����:O�n�\�4�wճ<d�E�l����Ÿ{�ky-cE� ����t��>� ��CzԔpS}&�Wl�
\���r�����l����eJ� -�z��$>bӥqM�5",�ԏ��?`����ˣ��,x�d�F�H��/3����dF��e��X�:u�%B*�V$�{���BbK�����	{p0�1�?!�|�V@@�Q��*2���>��E.-�2�5������[�
�q/����������c�&^hc��B��G�����n<"�)�ޤ�X̒�x/� �֤�w ?xR����\����$󜇉i��,"���3m�7�//6c(_���Z�Z���p+V����$����{DI��÷�L	2��Z��������L�)�D�<dM	�G�rR���ݭ=�4�vN�]�AZN�k�!�ݍ��7�S����>��$n��y�p',�B8&w�4��zU���k�����'o:�#�����43�����������\��D�gDT!TP�J\d�j&��h�71�b�s*�nQ�rC8��&Y/#��(� ,���2zx$�C`+�_w�O�ŕǰ7"�]f���Ag9����kT�H�ŠQ�J	�Ɖԁ�p��[�=3\F��cqB�z������ʇ9����9��-���E��(��"�9O���񌬧;�)�Fĵ�,�Z�Ɔ�:�Ԅ�Rb��m@S��/���ؓ[:�MK��b�[>�%YTN
B�%�]����g�����{41bQ���S��8�xSq���ݦ)�k	=6�$~3�lA%��z맕31Y|�S��mnr]%����+��m�:���ƴi�=;Rkw�@D,��4a+��
10M9�ׁ
'uD5�S�����&Sq^�Y����q{�\97��mP�u���Y�d(�oF�z��Dn�;��
�Z8�-z"�25 ��@�R&���o����&ɇ�gCfJ$C��a$DO!�_o ���2� �a!氩�Y��/���טҡl:�v<Ѫ�5+���O3�$:�+J� �)ߪ�$O�8J9^��2���C��B5VڼZ�J��K|)�/�M���oy��k�������
�f����8</��j�X}�t5Gn���Eﰕ��5YFтT��� ��=��f���V3���a(�B�$�V)n�����7�n�V�_�h��A��[���YZp�2�xI�>B*�j���@����պ=�[4yG�ŷy4!h���V��ۙ��
+�'-�����7C��� e=^��u��.��go����up�z�2[����;8$B���t��X���������`�����A��[<rp����@���dx� +h�kD�8m�̉�\�.����Ex]�Ŋ�yl�,�&��+-G��}$�g�T&�?��#��1��!���9&(}}3�>|�um����XQ��(<.:8ҫ�a8����[��yJG��}������q����J�7j����z�:r��vo����a��e8Oύ���&�JjM~�s������E�6��sp���Q�����_�{'�fyP�L��V�H�D�S�L�����1�<iU�����ڡ�8��;[=�c����h6�j�H�'�K�"���s�z��ZߞI0��~���-v��~�a��ܸ��PX[S�ܨ�XaN<�V�}B8������g�G=����Oۢ��V�M�xgx�{T�e�|�'��_O����<ut�*(<�x�EbΈ0�U"Y(b�����bZI���<1gQd'�2^�6������N�����0��ވ�a RYТ �M5�������~]�����p7��xg�r�Ƶ�{��y�!"ӲJcqCJ2z��s�0p�>Lx4[y��xl�����!�9ܴQ~�����佲��L��=W
��&|3!)�����7�(>z��a�d�[��7ϡ zx��<��0������F�B�(�� �\V�춬�	߮��8��zZ�o�pέ�N.r�*�\#�`gR���9�}� ���B���՝=��ƚ����h�{# �6��8�f�4�0���4�I��*�l�ޞ'Y:.5@7���L�y��"Q�<B���ET��;����+� ���Pt��~bdt�!�ʙ��1N������� /Kܟ׈-��¹��L
Xw�}�O�f��	�9��Pb�.U�\�HYZx�IC��-�*���*(������*[��b��~希�Z�w^'
:6���g׮��������mp�B�)�Ym3�,�eq���O{c)3��E�0�׾�_��?-�2��������j���+�*8��w�%����{ە�2c�43�Z��y����!��h�\�?�����i��7nN_j�x6�T�bvQL���%9���x&����}E<��=_y��t�Ĳ����n���s��}pn[���?�J/������E�2:@�5dte���N��~�]0AO8Q�
�j�g�87}Y��  OguH��o� ��5��Z����I��_wc�M���&�E���o�3�Ռ2]���e�P�e���`��w�Mf_4X��o����xZx��t2����&�F��� �D�d�5`B��e�? XB�z�h���_@J?��`u�O���e� ����
.#Ԟ/[M�|��^.�~=�^����g/��%�(�]�6[�`U`�\��N�l�l\G�P�����x�H�;�	�/2eN�	�ޒ/�f~����/��ԇ�.E� ��m0�����(}Ir�eH]�y�xqӸRq~J rW��?��F.��^�� n��H4�F	ȝ���>��^��J(�ޝ����i7���U<��7�����c�{V�
�k]Hh��n���G��3�꙱�(��U�0�� |Ҝ>��*_f��7A��z�+	�ܷ���0�nȽ(t�j����'�k4-�U	e�K|sm�}Q<"&���h�^�d�����_��Y���<�F>���)_��$�٩M���"��JY�����?�y�7v�9 �h�����D�F�o@��l��~\V:�	��}�QE����C�]��f�*[E��e��%�_�X�$�d?�X�|�*i뙌�:��;�ܹh�i����yRUۂ��U]Gθ��zf�s��~Q�5�����L���.Ob�ϰc�N�kB'!����%���^�-1��ۉ�â��?���f�)H�������5;YV�<0JȲ"���6�+�Gy��-�>�	E���!��v�efq\��?��^G�t��o�L1���6�*�w���8,�F>�{鯃��&w�6%��N�3�{��+��-����&�>	Ք�!�D6N��[�h���b������v#?Nm����*��F�UcmZr�1�J[��۲��`����O�{i�u���H�"xYb�4�0�k])Hk���V&�J�FX_���ڇ�<����7���?�4MI��j��虌N6�M�ZS#&(z=��E:�&��	t��܆\OVQ2�>�t`���;'`'@��ݟ��e�R����2_�x�/�B�%-+���÷�Up׽"�<<N"���72Nʓ$ΥeK�B�j�j���Zܧ0�[�?Cí�-�{x�% K��U���U��#�?q��S��blTw�,`��ԃv���D�q[�Xv��Y�7���3��YL/����g<�X����I��ξ�j� )���~ �K5��.�Y&P��PC�D���Ap�l�n�m	��|�<ʌ���]��0͕(�_j�`-r����
���g�1���V�?��K�JI[{��	�&��le/顕���M�aER���0����X��뫢��K�:.�ˢ��5��;�ag&\Jg|#2A;3�-X"=��/n/���ID`Q�=��7�ڴ?ub��,/�W�EAJH�c`}��5���>�
-:.@M���\Ysc*<�4��Vy~�Wi^6!��瀏=1�tz�lQ�s�Jc�&��_�_g�����n"�:��e�k[gٵ�͊�z��.��/�O�{}N���g�cu� ���c?Brׄ�r�c�'��[P}��[Q�ة	Zm��M�G^���B:|k�X���B�^F�xRGY�l�4���W^Ȧb��}�w�=�;�:�,zI��ӟ�l�nߘׁuB�����m���㌩}:nl�y���&y�w��Kh;ZT㗊sAb-]�u��� <�P�
���b P��D�b���p�k�I͹�l�p>/OHM3�ס�H3�M'�W�E<*�Y���R��A��;Y�w!i����)JD��LY ������r��n8$T>�S��b�j�u����}ö?��������ۀa�ڢa���2ˌ-K���-�haږ���5*'1�D<di̽�sq`���[l��C��"���p�й����)"�����J�Uڢ��t��f��KG2r����� q�C�-�A]�^0��e>��y�����3���1�6�2�e�"N��ո���4�?\��9%�)����_Ę��=Z��s��~�����i�(�[m܌�V�>*WC^���G$�p���9��9�F�NSA?t<�|�g$&����T�00�g�����,��n$��&�?��6(@�o��+�	��B�v$A#"2��H��G�5  PQ;��l���+�ݪ����蕎�:(.�\��:+ _T �̶f*ߜ��)1�a��'�l����Z�S��<~��#����P3�#�y�:.�Y,��]���
nJ0ua�o2ǆ�ڢJɆ��x���MlG���E	M�Q��j�%q��,x��A^��1��^ ��K��?YN��)az�N2��Nk�[!	�a�P���r����A�oH�ؼ���تx����,�t��Ǐ)h����E��9��-�nsHU���\ӏ,m�Ɍ,�ى�t󵁻�ҁ좲7�ׯ�رRi���d�!�!lŦ���ϼğ|���dD�.Ź��&�]��)��ٴ���[��A����C�&�TMF��O��.�"}Lc�+M]F����x��֬��T�������Nc�6~�9�P.�qlI�fg;����)w��ؙ�����Xj��v���CI�x���)���39�Cl4lr����D�:Y�L�\t�]q��؉k@��1��0�]ʃ�W_�h)�Cxɝ�u�{�E����eY��9	��8�H1�cod�z-a!*H_ԏs0�Q.�:��z֮�o���o!x�hY�~{<��y#����JL�D���QY7Ȩ���'o�a�g�\���u�'߄.{635��KȨ0�h��0��p�$��M�"t��7��1<�n�x�eY�6�5�|+�F�ĳ�˓Үp����00�m�S(S�;�֦p�^��6ݱ}���k)�@��} ��������J2��h&��2���;��P����|����*c���5u|�a��Q0���������"�mׯ6%��^�5�:��^S�
�����;І2�C�N�x��<ɑ!�
��\Oy�.�W�M�4�ݝ���ϙ���BD&�@SǮ��ǑW�S�i8oa��P��+�ޖ&A�d��P�gH���^�}ouY��A�h/R����{�?p,�c�,�����x���ɐq�����#V�J�U�0k����^��(d��8n��%�,���w��h�z@�����tk.VTr/ݛ��E��<�J�ؙj�G�I�	�+�zV�.�K"qQ�\I��͘��h\n4?(��*�7�pf4�7�W�����j;:���b��V�C|6y��L.iSQ13�ޤ�C��rl�� �]S��gCi����/-���al;Py]Rk��R���c�2�1�� ̬3��%�pm�I���}�m8�\�c�*{��M����PA���>s�c�ޢ9�����wt�Ȩ�
��T`վ��#�JE�8*��+���،�ȧ8V�%����)Be���Ts���e^+Pk;� ��֬�� �/�@�Vf���Q�F������8F��n��iQ�2\!���W�`Xh6�D�����hc��8j ����.��Mg��Ffaw '���|�a�Ŗm��&
X�,ғ��R	l�ɽ�_��!�,�|�#P_rq*���Խ�Kt��
�$���Am��5��8b��0���n1�,��٥�a`H�$�K�b��k�U9i_4!�'R���eE�H>&�$�A��:�m��
<�r�voq2/�40aNx�7�/�c.&�q��a�0��Y_�	���r8�N�:�8�t�G~�x-Af�0������~�	���#s�Ձ��iN�t�k���\$4�K�����g�;�Sw��w=A)0%iۮF�6@��� n^I�Az�����U�쌦өc�������A�E*=;$��/���i`����"�Hįځ'��/�ٚ�0u��g}�>&&��k��j�}����B�a�S��YXh����O&����|�m%81`x��ߍ�b���6-���9����6W����3[��T�ȅ�O�R� ��<.M�1X%��f%�Mt�g�B:��u�b�蟓N�Z���l����h�*�B�����T���6H���� ��'^}\N�Dp���%��k#�
`��j�l��^?,x��V��a^�A=����O�>�ww�O��ʡk�����@�K?@��C�M��"^\C*�t�l��8�����R��{��i�[��􂨵y���۲�����$�~`�jb2<{qf�v�5��SV"����>KHek����N}_���A�}��k����+��@w��0�zzǬg�OО�ݝK�� ]nz���ul��+��Z]�.UE��b4>K"�!A�ͻFj�91��"��Gw ݢ���[fgt�Rc�n���n{�6XE�<a���E��	δ��}M�,��<(k)I��!�v��+v�/H�g��y�����H�1Ќ���=�|�x��T-�v�k�dǋCvP�k� 4H���Ut��y�3�:���_��^���A8�{(��ԜG��Gg��Tֳ��2`o%�@��Ȓ>os���jZ�hǧIWm��hʂ�?����2N�eo��^uNna��y|-E��WŅ���?2�E������6�O(��k��v�g�sR�ݕ.�D	+���d�I9�m$s��`�4T��T�u|��`�h�/"1��pX����u)�h� ��ĭl�!Zv�t��M�!�b�|�P�|��3Lc9��h���)�:���S"}W�S}�_�sg[~��ɨ���Yǲґ��݉�f�����1���������H�!��VU1�s3��˰���f�~�r�O�R��Ԫ�G]��._	<�	�={wfgX�����u�.-���M� �����23� ���N�cvت����F����#�"�v��4�v��\s�ъbI��x�PC���t��j6�ziHo.y�L���Y����ݹե�#��u�t�i	n?,�Pl�I����%�8��M����kp��T"�� ����ѝR� q�7���Tcaʑ����{�f��^ņe؜h����4��;�B��nRv��{P��!��pO5�Q�ss�����}7Ģ��`�_�}��w5���?��# �#�Ԩƛ�=a�E4r"�{�D防�y������$jX�WW�ق���_� &�"��m�]�a�UU�5
A��K�)a�|�Љ`�O�}�.��;i��"}(6?��`nyQ�IR0�~��O��q�B�V�u�'l.�������µ'g�6 P�[�� �ms�|m%��]��#R��Bmλ-�P�a�xw�$���4'�U]�뭀SʙOdz�Z^�}4�읒��^2���9������ �b�lk��9*�3�\��P}d��p2�e]�B��1a���e����I�����]e\� ��8.@:}��� ��g���I7��n Rd�6���v�&���#�MHC�U��m����X��}��ӽI������w<�'ی84yܜH�J���
""��P_-� aTw#�	[��.z@������Trέ�>;d��*6��k�	������9�١ӡ�O�� �8$�p��n�K��7�gg'W��s��ctu���f "C,Y�d@�r���)+ #����R�ɑD����`A&|���~�y�d�d�{K2��+d��4��3]�;����(��jZ{�q6����h�q6zi�y�Xf5����ǈ`|�Ʉ'$A�?�������7���K/:�-����*6�����Ř7'Zh:�ǮI��=�+��&x���W�*�n����b�5'I [�bǤ�Q>����K���H˪* �<�w=�IO_�7�tg�֎~��e@�0|;M&�r��8����we����{;��9��G����t�J��
0;�{��S��������Xc��z�S�V���/���:����g0��l�eb��r��d'.f��Dƞ��&'�%�.�	��{�ى(�A��?>��U����饱�Hx�JZ���[R�<���-C�is��U|u�Od��STm����Rc�R-G��\ҼK^���������4�ܩ^�h@yl�Hp�	H{��'>����z���򳾢�N���m�/5p��o>���X��,q�׏4r��b�Qm1�&�Z�ys�jɑ	���-�&�$�Gh���i����Ml���B�U�O7��P�_�8���/^FJ�^L�5�0FweqaN��q��QuEOj�aB/E"�Gl.��:y�n��ے��e��>rJ�R���f!')��T�Y�B+끐�)�-{W�S�}Ţf����y�/�	�u��'��eC0Wx}&e���$O���?�W�8sZ<>Df���;`Ǜ1!/6�ªy���$�!˭Aߺ��ނE&�fg�n��9ι���ע\u4�L�<�V�������pn��2NxӞ����F�|՞�`q��C�A��{�m��NJ;^�$*��Ċ^&�J�Ɓ]~Ge񱑔LȒ�{�p�eK�'\b��9Z���w��!�=��0�y�ũ,�{"�Z���K�XQ����B�b�

���=��."��#X���p����P�(�&[S� y��YJ/��b��K&qV��/C�r%��W�%�O���3�k�~�xƆ��8�
�v�ȡD�t��$�o�֭4E� ��]��Xd�_)/��CuQ�	�]�>��J/9Tˈ
J$�^�EΧ/�-�>���X���M�~�8�Q-�b�=g����e�[��(=�L�qWHb��גRP����sD�T�I�fe7��Sho��8�	��P��Υ��d�
{��j����A�Hكm9T;��o̟��Ꞁ��}1;Ě��;W���S�1�P�i�3�z��":�u*u��L��rN�Σ?D|^�tW�⡌�f<Q��4���^��f\��	�U��P�C! �Ę�!�D=n��֟�����Cz����$�]��Yo�6vY`r s�]*��B���w-��\c�0�d'���f�n�*E�Tـ/y������%��^��Q5��}ͦ8}:�kڒD )iK���o��<Ks�����S-����zʩ��亪R�u�Ha�[�1�>#Q���O��v�+�p�~�a!��de��T
x��:{��0%�[01�t�1�V����].��,-ǌ耒Q���F�O�����4(�ɭ��NA�{&0B� �	�:,��D��������a������3��s�VD��Ze�W0O�����μp�l�N���[	�ۚ���v���Uvz�A��-|����, ���<�P?����龩����qa/�@^�>����m�T�^�*F���*)��L�ݺB���T���@�-֥p#)m�5�����,?Ý�*+ګ8ڊ�>&CiE*����&�G�z�H��9Y\@� ���[�w���R* ,x2�t���2�*�:��p>��8oj����tJp�x�/�E�7�w��}@�+Y\���L:��D|�^����:�V�f���q�.���єWJ|�Q"�(h� 3{i�KR`.���%g��k&x[�Fɛ_�+�{��e3�������
'Y�ŭ�"�i�_��5�S7=����J*�7)PL�j92 �`�.8_��PE*��'z��n�WL�c������qG�g�mrdv���( [�I��e	*x�۬硤<������{ig�7	<f�=�P����2U�a<����A����}fR���~YU�K�ˤӚ�[s�� �X��H��}s�ߏV��ܖ����YX��g,y:jB��6��C�����-觩5/�O ���uq���m�|a��v��8�e�o}%�-�b�M��hN�!����0[.S�Xyp=�w
"��/�N�55i	�(��������C�ɤdȄ�`,���eh������$,)QF=��%��b�ȈJG�	���w�\�B�[_�~���NԦ��.�2Qa����f�('x]ol��J����ڥq�ż�������mU�����[8��5Op1ȃ��������7��h"��	��:\�4k�'��k�Vf�!vd�}
��v�LD@=r4dԋ��� vS�y��lG�f�����//b
���,*^��kB��GǷl?
&`)e���g���}S£K>�D��s� ��9�q7ߦk�V�LI��ic������B��),%5��*|����SyR��Oڲ+d�[��P��B($ZƄ1=?^��@�9�z��C1�r�hK���έnC�y�3݅��n�M,o�,�Ŵ�U�e���*%d�[ˤ��yp�� ?�^2΁�ʕ�ʌmÄ��<ı�0"��G��5�n`ʫ�%��Ā+wYM�W�i^�g!2�*~�$�3���m�
4j���y4�A���C� �t�W~�Ȏ2��z��z��Opʸ~��۩���ƑB���qQ2p��9������������.�ӫ�K���?Ks�
tũ�&h�e�*o#vr&����;=�E+|��i����)��%�a�Bц�[��!�H3�&�or��k�Q,��� �V
�Y��cq���0���Ӯ(:f����d��Ȟt%�
GY2tu�5���� ds����6�_Le{rk���K,��l��-��L<��ׅ�{9��Z����꺁��<ȯ��W�5t���*fK���-/Qn&^�sWν�>mE+�+IC+������v�S��L`:�����h%65���9Ï���#��������žo�5�I��n `_4��R��8�o.aX��ݬT<�ў�a���t��- ���9�8��_u�w����j�3Q�T�Dh��,����-I�_�lBP�C����##M�Wr��4�z�Q�+���ؼ��V��������C��/m�U>ք@
��`[T�Э�C�	�̵�x�X�*���������\nUhh��ðxoM:��3�q��-�7u�Tw���g#���lv'�ɟ��v�U��8����ǲ}�
`3
^t{�ߩ'�q��sR
��|��ӑ�$+ "��9o�v�������e�S���h%<�o���g4��9�F9�b6�N�M�g`-���d�'$UfE�V,6�� ��ì�-DO���KsY�a��$�b���Ɏ'��}-%Al�]��~��ll�X^�)ňf5��R��d�OOv���"�b�LI��*���z �J&��;8�e^���q�w���Oy6�:�3+���5 ��n��� ��%�m�Y.�Y��B@I� �g@�9�6���{r)��LL�'V��BM�e��bT̐�:S*ũ�g�#�D���^�����3;�4�[�<E�"mIU��ܖ� ��D㶇Cr�a�R����
�%�;@БP:b۰���	
���dih(���r%I0v�h�̍ �#�ʋO�a$�0�����9J�����XQ]2|7�WI�1p ����*s���֩+h�DbF��Ԑ� �M��Ъ��oj8n�����w��܊h�9���wciP�,=�4j=�ܞ�Y�/�������2������⃮ �;���)��#��6��nй)��+z�5�u�.a����2�W��.\�5 �²i3��R{SrF_�\[f\a�@@��Z^_��t����)4SxS&a��nz��%?���ӞF����Hg�"��X��S�s����y��E �^�pg��#_Z�$�p0|/d�0��A�g���Sc;,�8�G�Mp�48��ƙ�f�v����~ݦG1�.����A��TEnR����!��ny�F�jZIZ�\Z����ۨJ��xy��,���e֤�X�Ԟj�$�J��G���<��S��âdň���l���y�
��*\�'<389��̘h�]<�����������]K�΂C$���<��j�;L[/�y,����V���n������Fb0�1��\��!���@xv5ue ��Ǌj���)?|�u�y�ϙ+/�F��{x����RY��&8��5ur1I?�6Q�˔8��:ȣ�����T`�����;��uN�E�����S8��B�ٓ��������m��N||�ƞ��ps��xKҳ}�����+Q�n��KL]�VYK� �<���d03�9�.'�fn-�l2�� �!.٫LG�ktX7B��v���3���s���-��I8Z���`>Ҿ�����?q�����bf����hr�"����	�8.�3MK&���O�}qW0&4�e�0S�;"�)�oɲ0z����2�Z?�
/p����(~\<@ ��3:NZ*�� &� �UO&���H�^����C$�h�<�u���ق�2��W�����k����+>-�X���xw� ���	[?D+��D`Q��ܷ�Īh��v��}����qh�
;LC�o5�u�e�4�"KG�Ɏ�v� �;E�8g��ɴ-�~m]��Y�l�.r���:>�P��+"��V���l�yM]b\��e�WTu��E8,��:�CVW�9�����4
��F`)�������~��pa���-��Y�M��J.�讉|���o!��� ��O,���;t�+ ��� rS1�������&��
��C��U����Ϝg�W8�Y��~�;�e''�x3��U[|q�RRn�V@�.���s.�&o����1�ke���J���D_I��z~H�x[i�F��r�yo�/!�f^��L�h�1c���~��$^r|�
�Jr��1��R�/����N0G�)�5�Ā�x�	����
�>�	?����8�VM��X-����| 3���K�bl���O�]��K"��֐���$�pكũ3�w��\�]/#�����(3�q�����u�K�o�E������T�D����9�_ZC�}P� �:$ׄ���޺R�%8Tqkbm:�n�T�r�V~j,�D�
�N��s�n�1[X�ۣU�+�,��'Pf�.�Pv���y�y��T�t/��g�y3�4(蟭
p���}h��(EI��W��Y��-�3	����ھ�}�2��S�`�潲�DF:>uWH��#
��̄K���e>)a��`���Ii�Y,2��F���Ŝf�����U��E���ڀ���Y#�cI���3��+��jV�ǿ|=�Uu��@��G�M2ڼ_]�kvc/H�	�����,����FOIs'N���\)�6����;�3�7��&�N�D�+�/��ŐA�hz����􍊋 ��
��aj��:�s���)/X�W6`��,�V���e�O!G��^�~��	�Զ~�Ϧ�V� � �M{�1J�[;�v��Yn��u�euK�p|0+�@�\����(A�����OA���
�\���Ѽ�ܸ���c&���1�J�}�8��?2���u����Z$�8"v���h�]mO��~��i��)�OapsLbO�؋]���+����6�$,s-���Zyda��oe%�����eiB���I�#	�N�,��B�^ԁ>a��hn�������zr�p�^�ta���|�sN�v�����
��ʆ��+�Bi��]w����i����%�j��`7����҂Y�Y%Ҕ��0@j����R�~������(".Ă���Y��H��U��#��M�U��/ezR�Sy��������,�$�Ʃ�W�Q��
~���Wŷ
>0��*Ak"�t\����p���
.X.��=
�Q�M�#�&�EyhsNbQ��� v��o�Y>��5��d�T�|x�N+�8m���q���~Nr��XYa��eY3	����[ə�-��:bGx���O������c���ЊAN-}�zr�ü��!.�ā� �8d8q8����t�l/�D�ݺ��w��ފ=����j��+e��=�X��Y��ry��N�������.���]�fF�����m�l��B�9�)*[/`G��J�̟�_eCd���J�h��ɰ�����Bm&ؿc���_��Z���|�4qqsO�dn #H�MC��^O�����#���S���#N��ˮ������讇���Xc{x`�\�N���O�5#���:[#�������=3�pq0��p���Z�*�����<�y�.l��,����2��r�3�w0O��������:%9�A���p0Ȼ���UAP��$����#�'��h���klt�(g<ʖ��<���4�E�=�d���<�G��˯��՟a3�����?�\a�+�*1�,;Y���n�'�Ђ��<ݣ@ʷ���ʛ�鋉�?�l�k��a�5��d_}�'Lˤ�SԒ�kM?r{5��'{H�A����W[ܬ:�[�Za�j�����6 �����cv��� ��oeԅ�P��ϲD���?� ���Bp��r�-�6΁�z�:xG��EU/j7?�t��	�_�<X�u��42�XaH���V�ƱѦ^S(2���X�,'P�#��'�@�V9K	fv��;�����!o���=T����|s�֕���9���<��������E��V �3�EP���&Ơ�;�A%9��Mj�+�I��t����d���#վ�����:̌��
%71�O�F\���dn�t�n��%�(� !����$�8�2����`y�V���������t�o�EK��Q��"�]�z��w��F��.�s�>�"K@nhFuT�M�JV/��pO���.�P��B�-�C�:��i�;<���(eq����L�r���\ZJP��;"���{> ��u����������Q���^��B5��MXD	�`Sc��\W�H��B)s`�Tv���M�W�T�W9���+�?��ܮՀ��/����v���/:� H��[�3ir�'Li����p�1���h(����?���;I4�K ]&}Eq0���`DΖ7Q݋<�,�w���*5&�cK˶rv�5�x�K|�w'0Z��D���>^{�a���w�	X��j��{0[���xl���ƺ��YBG$l*�:����)۪�e^h����.����A�4�h�da��8�X�(C������,��з�i����	���%ƌB�OP��W�N?�6W$	��Ԧ�$R���M�]���t,/H�z�h�JR�৸�����]�ޚڮO��q�t!�r��'W�pY4��W+Zi�̸�б�3��}"t`�V��Rq�5��އ$�F �#*�>�&%nL���L�Ѵ�#�f��:���8p�_�b:H�U�޷K��u����>����E��]o�j�{�ڟoYH�w�����tH���~Q���k���/3ȷ��M�$���)�L�H>�����mBJ�>9�>8(�V+��X8�,����#<�\�n����8G�?�?���+��#��M��BW����M=j�����8TE�	'��c���ۼ~K䲼�Ԭ�q4dУ@mI��A0��ZU�v�HИ��q��I4|��1.�S�p�9���~(���B���	�b��p�P�ԩ��Ro��F��;C������Λ�ʺ+��6	��$Fȏ�xR�8U�"�d*�&b��p���UVW�p�W���J��I�A��v
�l�*��];���.��C������
@�b��`�&�8߾!۵�i$�c�唙�U�/5�gfM�/�J�����,��ĥu�ȵ�TmP�&��>���I?�U����-�����D-S�e?�~�(S���j���	���1��σ���e|�tI7�E����z�Zڲ�J�Ų��Y�M�+� Mot/}��� m��$�����YE?K��$�\`ݞ?��f��(�g��M���3IH;~"��&���W�K�B�� r��5�|�߉���fz)��0F��!��o�
�D������7�J5� K�v'dὸA
8g%S7l�x���ާ���iC�6ɸ�m(51F�j�wZM1F�|���fqG�g	�����#/���`�ҏ1U�U� ؀���5��.GI��H��]�]}6Hm��9⧴�{%d%W*����ԙ<6�ac�ϟLX^b@X�@�
�h��F�*���d-;�@�`��o���q�,���q促�+��ӭ�)�MK"�b��*t03�Q�j�L�e��TI�<�/&�.c&*>��S��L�c:����QL��Ivwn��!��!y8d�H�cɭ����n�n�@�� "A̘�O��v�ۦ��ũ*͸��������5�*Q����X������}��¦��)�o��Ь���һ�c����)/g耴e��'�|f4�b(|��!ծ0��$�o���3��:�2A�q����jqm��¼Θ%k7c�0P��q��������-t���JE��F9�P�����1�O�7��C$���,h��tZ�^>�J���wF�FSs?�Ǣ��S�$����r�`*�q�
�������ok�id�FO$A]����S�Q�di.��g-��	ZN^D~8�����+wsX: �d<k9�N�%t ,�>@k����.����.����!��#�����3�G�
3�;�ǱǜAL���G�d�S!V����'��#���jFdIq正��(�~��P�I�n˞Ս�h�j� �Kmja���`�=�]�n��Kc^C09���u2t����a�Q�bp*�����6Ė�ꮰ#���9��M\�z�^�����R舄&,ѹ�J~�>�1؞��7�Jx�J���I��|�Yޅj�Ͽ8���ȃ����l�ү��e`�5!�H�
��['hvz$#���.�(H�w&�E��3�n�~4��^��+4�Sq�����ջX��&�y��}�P>��0��ꨠ�k'��}V}2�&jK�\K���InR���#�����ixJ����M��fh��(D:].^�ΰ/�!�ht�[#��z�O�=�m��}2!�F�,/��m��PQ�N�֤g^UsV:S,L��p��G��Y���9��ϺߩW�c��$m�;4�{�ӗ���"�����p�~�WIf�=Yк�!)iH�j�_)�5�>(�ƍ�|!#!��|�TL�3�X\t"�d���h�L��p	�vLD��F%cYގ�X%��O�~^ ��(����/�W
���xK}�ĉ��w3?�BJ8m�G���MUk��KϜ����e���e�7��dy���|��-�7j�؞v�'��}K/��"�Yl(��d��bQ���j�����j�`� x�&g�>*h�?5x���Ng�۟��RVʭ�"Z�I���^�=F�� `��&Ʒ>9a���X��O���}��k�^�R�-���2�[�׫5m����!(�џ�Ez}��T�昤��>ճ�/��f�<�~Wc�!��{<n�C���T��iy����Z�IjJ�|���z9�Ǯ��2A��N�����$�V[[w����K�,���J��p!�6RǤፅ*J�אT0K�_ ��I��jr)%d�3��9���2�q�V��-s���� �g
M֖Vc���m��w"q�����3�ۿ��&t�;�Y����W���1C�k�(��i��vӕ��z$�C4�e0�ݥ�&��(P��䞫n�w��F�Gv�	���j���#b�/�L�Cx
"�Zp�&L��?nILWKdT��mo�J����8Nt�L_үhԁ�4��q#�ILh2��<�@�*e��j	k��h�e8;>��۝�0��ˢ�|Y8���('��)j�1.���^�bM�F�T�E��xUqE����H�3�����L����=x���F� \�˿�ۇ�d��+����?A+J�>��	~1�j@h��p��.$���mr�՗t�5h��4�|��MNA�1�7/�a`���=�m�N�7��S�5c���N�r��4�
���e�_�O�Zd����u�A�5j�.��:��iy���Z#�䀶��|R���4o�W����Wj-/W����]������>����c���kTe4s�5��&�*+iQ	q��L3s�C,&��`��P���y'9M�ӻA�a�����^���,K���C�w�ı���ש|��1UM'�%R�w)�N5�U�y���I�4}nt �K����g��fqf�_K+%��)}0Y8H��2I��Eշڊ�8Q�
�Nv�C�9闄w� 7^���ֽx�@W{�������f?�#`<h_�Ǝ5�)\�TҾ>����ݨn 7�;�L��A��gN�~��U X�&(H�?נ1��T�=�-̑.�&/%�S���۳�N��� ���)<
�2?����~J�;�X���f�`g*&��R�J),�*�:��47�ZJSI���W_G����i"��MͰE�y]�Q+����U$+1-��mzIX_�rw�'�%+ȼ�G��^`~�fߵ��y�+	˂�*yO]�������Gn��3mX�Ί�� j�YVs^�p|uX)��En��<K[w`�)C�+yW��&E%C��eX��؍{�*N������\�`�b ����}_�#��H(��wPɏ���eP��ŀs�����(zp
�`���x�4��bʵ©Fo<��J)�i�T����>*�]&��a:Q��f�z�Q���v2ML�������w~Ң��=|��M�ֶfM�)�ڐ��bb��T�ٹz����~߲�&`��K�8���z��Jwk�2�]Ab b֫(��
~���[q)\9��u�	�"�:�@�-9�8�}���6���4P�o��zKٜ���	�+g�k�_-��8e�H�w�CD���4K�TD@`�Ql	���wSFB�\S�Cv,�� [rO�&)�����ARJ=��E-�!y����cKPi����x�0<�P<����:I=��È!�;_�FAi�8�,g��ۿ0� ;�ۅ��kAVc�kjc�o���a���Ϯ���[Y��K�]�r+i	�N7���'�)U���L:J�p���i�� >��j�P@V�ci�%����x� ��� g͕f|.5��^fm���3%�k�
�4/�v~eʺ`�Kc���ԖG�2B�lm;k���N��@��qg����O��'�w�T�WvTi�&;�&C���L��e� d�~��5&�����՟�� ����ƫ�(��3�������~0]�U1<�L	+4�� �g#�y�Y�5�����=wW7�z�1�З &>r<��K�D�k=
�ZP �q�#ܴ��r��;(	���J�ۅ� ���a���_��,�I�X���]�h2�CI��}�PSEϺ4�\����H�_Ȣ)_�e6�S�/NVB#6t�]йM�:0�� H�ZI�m̑�a�f�2{vHT6�7����z��v��E�;�� ��\5��Byv��n W$�t��ݮ*t��\� ���0	jg����&z �O����̞6�n�� ̑<��9P$�\��m��S�����^�*�h)�O	��:9(?�&y��u��7]Ya�
�����s�/��>i�,©����E���⑜MK66�C��|��[P)/�w�'���,���Z���ʴ���La<�|si=o_�Ц�τ�A�Gt�0$�v͋�b�T����0t�����yQ�t�JE�Oo;=��
@8߮ב �y���l|4z#:x�{R6:�N��0jWT�,�o��k�z�����Ā��y��B��@ԋã����U��;�L�!Z�����x@�����F3Y��51�7d��G���]?$���fg�r��Qm�����:*k/\��B�y�iG�h�S���OW�dM�,���;B~\�w��w�e�Vy��U�!������	�h8e�+�j~ɑ8݄a&ݱw��-�%�W��`^{f/�ypyy S_XX{���D��:���yk�<���nT���]���64���wX6��#�I�̚�����P=�?��[�&д{�l��:)f�Eon���6�N��
��C����ص�)+$��8	=C����TB�	W�m�@pʾ�RL2� ʿ���Λ���O8tN*��'�����:3��֜����)�B�5nCa[�x�1��L.��`��L����n10�~{�����;��Srƍ�(mÒ�gb��b�x�E�l��"��MoZ~�KZ��"�F���F��cX��p�����T��O��@��"���πж�s�E^f��z����J��K�����	5����${�~5�����;^�C��.�0,�M`䩈w��1PM�˰ǝ�0���ҧ��q�(
�Q�D�ǡ�cD�ڹ���mm�]�ɢo'�;҅d�����|k~�4Ye��yf��m��q�b�y�3_�����Z��ȣB�nʢ$�	�Һ��
\8Sp|D0L��A�i�������U��$wJ���w�uNf���>��Kp���j���Q�M��yD0L'����n�����i��p�x��҂�����Φ����-����Aݾ���iV>�bDM��;��p�!����A-xk�uE��@f�ͷ��E솝��߰���|J��ٺi��V@;��
gN�r���2wS7���뤓�ߥ�R�J_&�䈽U�H��D^IYHvQA��[�䑭���4UY��}�	��6��#k��<��"��uO�p��!p[	� Sk<�>�i6���P+����`�Q�J@�������%Z[hNg�hx�<��M3/�
T¡"G���HJ�Qۆk��A�gW4���C-�Jv;��0yv@�^�M����w� s㑇�m�l�%����2{<870/��8�K����{�)ɜ��������ኈ�8(�<.V-`('J�E�'`����s�A}>(�� ���vD�21rQq5o\�x�E�As��i��*���k�n~�T]C*���c�Z:�n�D�����
ps��T�u�����W>�ꁼ���ġ>��ئ=&�l������X\��e����rC�~b�2���Z���qw���I]�A�
��"db�Ǽ�G��e�%�k�I�~`˘Z�ǁ�kJ���5ӥ
�N}#��	�dzY���b5T�$���v�?׷��"��OߏR�=�x��쑅/��2�lQ��z�b8��X���^}͓��1L�����̫2�S��˜����{�ʶu������c��M�1-/�C���ymĳ�Y3W� �7y�����e�$:����lQ�ҁq�8�F��d��2��D�R;ʀ�ȕ��Dn����[s����J"ٴ5��R.o��j������ jȉ����1ݼ�D�G���{y8�)���D���m��$_kK{y�p/p���D�~�"�48�t��Oy}}�ӿ($T)��p��b�^>ʝ8�ۮS� Nڣy�i��=��8��Y	�rZL���e{��*k瓒:�Ɣ}'�t҉ /<�4i�#|Rf^��(k�y`���"|�r���pF~��훀��J��--��
�(�� C֡���3� ����I�_(���������q���<��ߛ44HC�RtpRM;c(3
��\�"�[��v�"W�k(��&>�:�'�2�'���@8&	be���a�hR>��dm������E=^[����0�М��V�_܀�%�TV��vl\H�*���%=҈Z:���'���u�f����ʟ�tg��J�0��Z�v��+Z-����?�w�D��V~����\��UH
��Źߤ��Fw뚙�ݢ�\����z0]W>������)�ӯ+z
���hpk!UZ������O�]̩�e3}n��=�ͱ�[�8�3�/�;��L���F�!/��������.c'�%'��1�u~�͗�����@u�@D���-��o��FXX��I̺�>�t�e�R�t+��7���]���;� <�UN������l�<�F�$t^BW���ϦDd�����ꤤ�@��P�4��/7ɣG�!�ǀI"��:����YUrs^�=��_S�$υ� ����q-�![\1��hNB��ι�}I/��^$�S�n�⊧k}3qw�t��E^7fp�/�������l�jɀ��5Gsޛj�r�^����J�|Éw����R&!���q#e=���o)�&?�DǱM�\UgF;>+;�VHR��h�As4��=����QN�}��,!���+xBC�I�ˁ-?l$�����:��`���'��m�jn\��%�+��
ka
h�]��_LJ
Yk��
���}��п����f����Dᦌ�������;�'v"b��X
��*U哻m��3��Pnw��`X�S�N(�ѣCY��-/b{с�.�f*� �����qR����;��ذDZ�K�:EP��ӎ9�ū�S��XY�1��2��޷����!�z��̹�[Dt��L��k��6�1����-���Y��M�(�̟\��@6��␠����nB��r�(��k�A9R����L2YM$�Eꎄ�	p�%���vS�,��c(;�5�q�{���YjV܄���*�M'���k5��5�r�/
|��|w_2��
�,�@�~�}?B͑m�c"�����
��L�����H1~Q�Kx��$�IAy��L�%:��V�����:
�P=���F��ncf;��*����e���XL��8R:O������2:k.��"+��M��Bw4G=����H�>Ɩ��ud:����
��
(Κ�*�o�ֻ��7�ԌA�R������)^�Y#��o{S�-�ݓ�99��LU<M�쥴�}bĺ�b��>'_HM��5���r&�v?&f����#��=�o�����F�L.Mk��8q���.��4����l��OX�d�	g�H)��M��6�YF��'�D��6���[��H0h�����2��m�%Ӽ\&T�.7���Ǵ��t���v��T�e�O�0����s�{;:������ ���hU�@�� *�n@� �\��`�Os}��#��~��4�a'��k2�~���o��,]D�l�#�c)�P
��CpDZΡhF�
vr&�A��b.���3؇ߍ��r���dN]�� XU�{��?��nl�1b��Xd���CVW+�d]���l�N��ݡ61|������X�|�мN�k���T�8`F*f�_����?��K*��8M�۞�й���k��l��O�bU�I�0G4�w�$ߐ�"��k��ѓ/�*�r��(� }�r l�GE�MȎ9�X>�����F�7���	��L:=�U[O!�vJ#aᛁ]�����.Aj�
����Єv��r.��X!��jǽt�z�
����[�����V4`�� q`�Z����	��@z�q}l�.M9�ZY���~����Y.E�9<�p^���m���yx���"��l�f��zq�+bS�LK:-^n�m?o��c9(�2�?�hK�Öɭ ��c����D;@�d�����.��b�a<"��I�Y0��=p}���-�HR�"d\'Ҋ;��Z���@�2Z�<2����lc@�u��-;v�L�)�h0mk���o�9�O;��uHz����R�@nB$�tHU���d��iQ�p��r%so�7]�;�A(�g�`t�/�k�CU�?���T\�b%�=2�����<�;_`���!��<S�S7	�*��	O����[�
WR�@���:@��`��Rxe������C��{�&ѕ3�؅-���m��
�?ۆ���rI��r� Ύ�Ӛ���࣯\�I�D��Y��A���"������&U-�]i.A7bgu�Ϙ�eԶ��l
C1�ȂsA�[a����٥������y���Jv�tL��T���*�B�?fޗx�ۿ�����$�z����f�S�jj�6V0����GA�	�wd��C�7#[4��n�BYvtb^֔�fp�P2�owѱ�ש��O��0�����dc������BC�.��9�N-|�6/��*��)9-wTY�����]6��X�O����|M�w� 3Q`�Y��`iV-p{�)�R�j(����O{����(a � D�Y�E����P��s����ϚҺ&X�T���3��*~��jf�XG|���K���Wh|�M4�׶ʵ��«1y���	1�Я��K�oq��BV�EN&���mD٠K1A��˦d��|pe/�;��B�p1�Z�Ł�9H�Y� %�pB�Z����n[� ���A9�E ��ƌ(�~Y�C2U��j_f��Kn}��tB��i�S�G�ؾ�o��!��&����_�]�e瑝%�9N됨�qnm�n<�Ċ5f�i��ٔ��{����� S���"A���:���n��x���@I:	d=V�K��)߿�Щ��g�r��qv �"����Q)
&l�Y�}E�B*o�:�7��W5�5
ӯ��$���Vi|�J�Ԇ���S�
�_y��n�]���Nj�: ���]<-���f����*������%y�UC꛳���}���in���CR�P+# :�^���0���J%�U��y9�OpX���<�{����	 蝫�M���8���&a4�w
4�C��JG���.��Y������S�֥'��/j��mh��U��� �n�睲��Y��v�XN�A0�HXߞ����1�ME��y��Oz�Z����G_��,���+)�]�]�7� �w�\όQdf����c���=.�'��s<���Y��^:��*
�������&����<��a�����K�I��-l��.G>��-O��ɪ�ϣ��OI7�m 6��~�KZ�?������R5DH,_%���.Vc�5��ؒ�.�~u��W�<���q����/���+�̜�_Mw�̦��\I��6��*����¡��������㥾���\r,�3�td�W ï���w�S��y˛����>���f���#���$|`��v����wuc�Oc�=_\����#��A7��u@&Z*f�f�Q�B�G�)C��6I���*6C����ףs�αYcބYmE� ~"|z���^-��7�?�eFw���� =9S�	��x��D�p���^�+���=�g���QC���9;Ɍ��`%H+O/���H�4?��:�kޣ��vk'փf<zs��!k����WZ�	��ei�=T[��\��{L荳��%Q�Rr�'�l]}��l,���� uH�e�k���m�v�?EE~ܐ�4��.<�Z���bX^廝����lua�F��O�J�H�]-r�j8�Z-v/QAc��)���\��,����H_����1�=7ۉ�h�K޻H�B���ߩ2�y���\��Y\��d�<k�P^*�]�|SA�܀���M����t;O���%�_�b�c����a���w����'��ʮD;��,Z\G�ؚ���O` 8Z��bu�`@Y�ID��r���hT��d���_�6�;u����w {ށ�ě���K�XI��*����,)�I%y��f9޲k���G��0j��������A�<m�Ԩ�k<���)�R%e��h.� �C�Ǐ\��M�����)�{2`��з�u[!k�=�%H��[���k|�<#q+P��7���?��?�Vv��a��%��e�t���r'�eH��j��Q��=I������*a5j8,g^��7��'6pHq�# "��Ky��t<tL�]�N�Hܼ��h�)q��0�j����*����:e�̓��#%hnF�󂒥��zu�U�)	q��S�mhF�G���.���5�-��xO�q�L +��m�{.mOd�=Տ`1T��V"�Md�X�,���z��C�~v�����X���~jW��k��ș�������uzd1�蒌��p;��.b��� H����dY��,�	b�[�3��eh!å/y���ȿ,�V�]�g��3j�{I�{F/p|�}��<��@&Y2��(����u�톼�U��<�x��S|Cj�Pީ��,���Q���~������p�����}W��ᩣ��p+�D?�>���4�^Uo�����W�����vě�A(���di���J9�qx�6�I�s���Վұ�����ΆƋ��� &A��_��q���"��)��(�їNJ*�$#��ٛ�v\��)k��9�$�+���Q�(�W�ׂ��D��Jbt�b�Xk�����E�e�}���}�#IN���U!B�T�ܺ�:�w���`��ǔnTě�BD��e{C������%��8�A��o���5���'��,]D@�#
t�N	]'3%z��W�a�\��p��D	�9X/��q3���觞9�����/{���^ο�V��U >s�K ��W? _gC��������dF_�-��vЊ��?�J�Lvr�w?^�Җ������&%�e���� f6�s�!�hR�)�j��Nxnp���O6��6�5��uER�Y3	��}�;�$�\[҆��N����1lg���{?�]���g5U�nnF��Mkw���{m���<����6àH ��`GX��k���7_��jj\h��猇�~.��OC�=\#�s;��H�#*�!F_�����
V2�4��'i˧;�
��h�$�����
�&Ky�o_���9����ڕ#�c�d�0�Br��PT�9�BM�6�7ƃt���}��w��^|�W�m��-�1�^ط �b�L�u㌢���l?ɑ~-��0�f�B�����q_:X�`�%/�Q�C���>�p��0J���'��Hz��̸���r�ЖIL�ړ�Do@��5ũ�ib΃�G��wTɭ�4��Փ�B?h#(>��ʑt�����N����.H[7"n��C
C(u`���<6�vD��P�ƃ����^I����2��֒�;O���(%u�Ќ��{i�'�ORnT����@��3��Wօ%l�**��i`+}F��$�ӿ�$�a�5TCiD�V�O�mIH�i���<�7[��B>P�������"�@���E13\m��=Xy�機F�߮/�FZG���ޅ�CT�K���J��4��>����sa9���_������s���PCWwS���
�|�1I�V� o��ڹ�/V�P�/TFI��֪6��s�)�8<�c����z�z}v'.5d_�{���)ʊ5C]�+�6p<A�������<�+/g��/�!��h˹A�kץ��C�c���m���%3�Ts�Y���!g$)�&�����Z���qRDJ�Q�j�|ss��(�� ��2��)�'s\�23��N/�[b�t��ᆊ#;W�V_��n l+�B��r0��tA��������W�R#�x��r��ݴ�4��)�a��پGT��Q�2�E(�W�#L�LmgHA�B#O�=�|����㰬B�����_���}^(��&�'����->o ��Y�Q�r��V�+�h.�A�,�˴��'���P�-t��T?x��2N$��K���B�FՀ�)����]��t̙�H�gZ�a�A`,�ù1�VBٿ�O��-�
���3��[�Q~���o�"�k= �k1z��Y]�UqQ/�؟�_<#����)�ߚ�L��\�ߟ������k�s$�0x���r�)�TV��)[5����_���]�G��H��u �u	�o � �.k�[<�d�It����CQ�������{�k���s�ɖ��̧��AE��K�%"ȋ/��H3hW���A#��$Y2�<<�µ�n�l�|a?Du�$=�PǸ�����e�(v�NE�E{c$f~O�J��ȧN��=��b�^Y�Dj9�{.�$�֡��7�W�Č��e5zi���ޜ��9��@�C�eG�=����I	�x�k�;)D
�� 4�ϐK�	���ܻ誉'��B���+�^[���!r��p��h�%���؊[�c1,��.�P���s��N�����&����N�?s���yw���)"H!��;E
`�E�K��CJm�=3O��c�I�n�7ǰ1�׸=�[b���%�6�;��or���7eet"\�G)�:P�1��h~u�c5Y�0t,���-�M^��Z.Z	4q�cc��� 0�E�O���{ʣ@WMc����pބv	�j����C=�fg�N}I�D��'&(��|P�x�4�V���OP��l������b7�p�i�W�R��1����E�J��m���>np�$&t98{�k�F�P���p��u������P�� :H#�u�qqr���Yt�+��	Rl�2#�Y_R Z�j	?N	�#��U��+��%F�kr��"s�b��s}��IP���f3�:�E��Z\�i�4��S��EhTY��F��&�dbÃ_�A�k:�s�L���"tjpNt�TD8�;IC|G�=�M�őT�_�,f�
�Go哶�)���տ�Tm�Jۑ��c��ڠ#-�����������W����(߅j2�t���(�O�F���2�P|���k:t�u&4���G�&J7�{��̢@�t�j�gd�o��B��s�c��^��h;�Z��a�VT�^Nw���;py���1��#zɌ����Ӹĺ�kO�Ѯ�hu���	�8�;������?�i���&/]h�+ЂyC��43Jo��o�E`��1&k_V�����*���,�t�Ue"�`��%�<��?�S`�[���5�z��>��LoUV�.���� ����w_��l��8,�������ȉP�xL�<|0HK�!�^R����5j��*���b�ޯ+~�����O�9�Z�3�p�RRX!I���R1u)fD�#iV�)���Z�hrw�h͟����M���4I���S��E��p�[�(?*B_�����&�S�!�#���_<��Nr��H�7p̧%I���\c�f������F v���Q�&��Jj� ��(�]\���<���.�Mծ;?I�C;�-�H���x��`���J�R��͗DN�j��yYgݞC�#���q��p8<8�`'�*DT��@HV/�1�66��q�@A8�S�����(H,j�x#�~0���ѶW-����F��z�݃��1GE�t�wx��;����c�u�<ڵA�U"��'*Ca�s��������}@p�M"b
:�@G��}X��1�ܩ@I�L�-��{�/�ZVz��D��zU���&���A�<4,���ӦGx���_ᣫ���G�"z3V1��5�O�i���,�Զ�R�F���~�J�k[/EA�S��Ӱ�U�cv"]jtb�9S�L%�v�o��i��6�gB�E���͕�;�`z��=��}�1�!�{ģ�U⊇����ީ$1_-u(�XL`�\��ҟ,��s�ys#�'
����A�������7��8u�A�Q��;Vԧ�=eX��P�)����~2_{i!��Z8�И�� m���⸎�$*�L-��i`���9w<Ow��ػt�-���P��Bgl_��F0�����)�}\�Q��j���~��g~�
d&�h�.�pY
��]�9��mʮU?��ӋbC
N����e���~mc��ao����J�/uz���	�rY��,sQ�0�ɌY��j��=�¨��p�	�I���5,���( p�q��eL��4M!��ʿwt ����1UƝ	@�h
�y�N;�=��J|�z�q'�DN �r�)����b�-(���F3�+�$�lf��������w�� `@7�6Jg�hI���)`�oR2�4��"KM��.]RF��Z"�;��y�yN���wiI�)���<k�dt?g�j�ݨ�QPn��+�ɩ�.�����A��"e�\3��ʖz��`*߹<_��b���s�4d�h��l NGg:i[=N�=i
.�@l��x���)vKZe�s2��
Ժ���$%v�?�ښ���3�B�NS���ғub���D����w�O��N�F*HT�4��B0�>ew��{6Y���/��f�-�hSj�g��n���$��PN�3,�Մ�w2�z�Ь��k	W}�At8��d�"�4��A�jzf��vѳh �T���{�G��j
�%\兵��&w�c����6\�g�d�{�3Xp����T��k;H���|��o��9�'9xe<�� {Z�s���Mu޿/:[a��?��-Ԛ�������h���_�j	%o��D�0��s˭(���I<�w�H�.�	�ˈ�����-ϳ���dF0�Tʍ�����p��1�6�H�Vq��J~-&�ˁ�Ff0��kqRQQy.W]PڞZic`7�%L��X*�|����PB0��L��6H���>n$���nl&7v]ظ�ơr��@(��:jg���l"B͘α� mܡ�b��ﲑ���\��L?'�J�/f��2�����\+H��QUdKʨ�n�tc�:�p�.6����F� ��W�3��4z^��<�OZq�-�f�t��d��K⹐��
���x���*�0���j<�|���G�5{U�B��r�9�F�����2 f�}�_�hd+������O�TW(%����&׿�YI�J��f^��ܪr`�����YZ��
e�c��]m�r'��eقT�$�Ze�����Q��oWڲ�aS@��H������4#�I0�y�z$��}.�p�n{�A^|��b�����Ӊ+� !L3�}��ŏv��=�trTܿ�yj�4����+�A�ebs�쫋�P�"��.�k5��W�4��`�S▄'��/� ZI��7��fv�v4��*�Cd�N9#/��z7ܟ���b��r�N%���3�=�߶��"W����#�%�?��(�d_��Zq������gå>�7
x��+�A:�� {�O�eR�G`�RߢU�|>6*]2�ji��n���4 _-xye{t��g���3q�砫�;�J��3�'��3Yn)�n��&���O���X4��2��*'���Θr�
@����p�cAA�^C�bX����%J؃Z�	�+t�żib�H���4@�⬪��Qt��-vG�$E�ں�,g����\��*"዗#w�E�;�{�ʎ0Rrk� �*о�4
O�T_
�lt���A{�ܾW�,�uos��Ƕ��zT�u纄8Ce�)Q�B�ȳ��M��,���8$����o���xI��X2-�	�����h�L�,|��h�M��ޗ֤�l2n�qq�O��V��=�_��P��P�t��V2T?{�㤃X���Q�-��C~��BM�>�=.��˂�3?qX
�:���L�<��%�\+�r���_.%��j�ȯ�xe����������R��V,�������c�u���QH��(C���bFsq�awM�{6[E���H&W($|k�����H|���m(��u	�����v����H�n��AT�f[GzvD���a�5D�T���ŝ5J:�	@�0��X�}感�#s�T:a�m|�P�upĒ<�uL�ce�3%KVy%��K-Z���C��<Ҟ�TX�WǕ��
 <{w��8��~b�i]�#����-�#��~:��:Ce=2�QE)��J��*N�(�����Y�8^����`��"L�q[��l �0ԇd#z:�s�e�#��W��_y�*yP�m�7 �v�_?lB��ާ앭{����n~�η`�ll+&��s��N������|>ƚT�>���\�d4�c}���6
v�KRW�en4����O����?�۸��0�8�ׄ֗�s���1�V%���P��r�U@Y��a�L���4֞�b�(���P^��
��زM4i�"'�S$��U͞�U��ۙK|CF�x�l�{\�GAM{�l�����y��:�il�#��G^fs��JD�<���*���ú6�E=���ے�;��XS�ʹ�l%�Ax·�ѯ8;����Mp�9Y����N��#�r�p4�t�ajB����K%ltgS[��(D��$�Ɛ��p24���0yy/���9��~�HM���C��J� а	t[�ݷQ��/��R0i��`��y��U��:�Zt՚~f��',0��-#~ws2�e��?2�sw��+�N!e��d0۳��'~/pJ����"�`[���� ���=x#�=�Y/44+�V���##�h+�}8���И�V�����˷��Tq��s��鎒�!,�V�I?�Ý�vӿ|��QFC�b`5��,	����o�x}�ox� :��F�n�$[`G&�iw`=���@�eـ�Y �T�=�>���y�<�6�U��w�KP#��{��sV�	� qEq�j�[�������NN�;������]`�\E�f������>�ϱ�Ԏ�6%��@�n�l~vL�N, VؘPz{�ܴ0QS���%���I-���YS�_o�f��QY����)�8��p�n���8�M�	�7��nW~��;�X��ڠ)ֆ�P�Q�YI��[����U�Q���nۘ��6�{iv�����on'�d��K�AN�'�;s 4�5��=OdP�E�`+�	��,��j��������$�f�3\� �G̤��� �Qj��Ѥīr��J�g`�/�4Dl�E�����#r�i�<�+��j�L���AѐuށKh�敍Z������:[U����e�{�$��ұ�	��F���ipH�a�``v�t��o��#�(�J�⨯UC���q�B��������,������D�.��bG�ev��4t*���ӥ
�N{i��~(b�0���
��QSnM�T5�߸!��2�v�L��qZ�\���Z�];t)�3w���ꛉM��FI��q��2kH�6��9�s��3$V��5�%�fͺ�^vi�;�A�e/Ć�!�O�TM$M�k_ݽ������n6��J�ȃ�\л�B[��S�2���ז.�g]�3�#������SX�OdF��c�{h!S��]zm�b#�Ҏ9yr{���&L�$EBƴQ���$d�C���z;OԼZR%������[�-�Q��|<���tI���C����o�&�	ʤ���Yc��\���I'�t�oU�:hÏ����\�C��OC%�9J�%�d2��"��HWל�}^�}Z���.��OyK�2{Vn�'�2��}./
<7מ+���/�`��`e��u��*�m��(�L0�r�91k|�d��0S�<��5,W�=��4��d�zZI��Y��ڵ��ђ��EX9�/�k���k�����oV|J;r��7�ݸ�Y��e�ؙOD;��HB�/��5_n��Ѣ�J��,& .��[~��^�%�Q����xKt*;���F7�6��p�Bw~��H��S�zo�HO4�C�b��%���D��"�n�z�"�t�Ձ~�x�V���)�L�J����SUx��=��/�� �/�W�)�5"�Fo:3���I��S���`�FM���7��#��� b��U�u_�S�t����M�˖�ݾ#ֱMH��-�$�`kK��Use�� �9��S\iՁ���ɢ�ެ�����ç��Z0͸���7&؎�[&���Y@�d� Dw_�$��ԍ_�9�@�]<'��Tz�~�A{4�uj�#Uxn�:YI�ŕ, A�]�K&@_�HP'n�:�)�@��4���*��ʱ&x�U���dB�~_8��`:S�n�^�u/<�)�iͬq����*�#J�L�.hH�g��fBf"]��q�;f�D�P�հ`,�5z����� �"���ˠa[�ڑIw����0�J/8��6ub����o���<fVK�b@r�����g$��F�v��Z��Y�����_6�����T ?�'S�������J�� ��	 Z�0*�ord����]�Fa���j5-�=e�b���k?k��"D�4Χ^Q��<m��e6l�	;߳U���_V���ka̡�����fB�����4�E��'���;���d#&��6Ae|_Q���C/G��R�߆�d��@(���-8p�z�}B��[���
�R��V����z	�/
=5B��q����� ��0�֞�z�]�{-�ٵB�Or@ں�Hwv��h��F�@vf�>IYd|��	]w�u>�n9�s-���(���p4�*��ʚyͬ$��Ÿx��[2j������Xcd�W�Z�� �v�W1��*��xV�8 �ZS�+�	��p㻩T�F��ih�����	��
F8�E�;�%Wİ�m0�`s�z�G�@.�#`���:-	f��3�O���ǉB�E)����������"�-e��H��*�.Y�Q��6Q{��ٔq�6��"r�<�6���н]JbfE�����;3��Kdw�e���(Ӱ ΖH̱q�D�auL e�qSφE�������T�*"��������7�p�%�/�@�+���k���~rѨ��T2ʈ��o��ϻ��#KMCqs��&FqB�"GqT�����x?�4e(���)��c����A;%��y� ����wꚪ�k�a��=���6��4(��3����ƌ�'I�`�E!��m��I� ��2F'�hޟ��L;nS-r��d~���4��J��(����
�K��L_d�^G�SXb%ad��zt��.�xyEu)z8,sxH�P�0al>$��!wAϚ��p�v���9���
��|�/�ȣ��1i�#�5{d���b��)�΀f�̜@!�M�C��Xpd�hg�\��3dՓ_�Vd�x��'0̡����#g�Yu�x�Ŵ���D{rH����D�j�w	����}�ѵ��0���%*��5�u4��!��B���ɵ�ݬ������CO�VbF�uҷ��*	�R:H
s�G��W��2	�.��V*(b6�����G���\������p;��*R�zq�+�)�@������ŷGa2�d�7�z�����۸���֬>a��*�&��e������{]c&Z=z 
/Jyѐ�v��I���ȷ%/`V�!��Lx`W��ŉ#��h�(K�=q���nxAF���f��u�+C̰�����
;<U�:����"�O`]��.#z�	b���-�k7z0�)�#�/*q�5���TW��oq��`���q�a���V�ٟv��CNg��l��ɕ�?C9$�P�$�X�%�g<�O��0|������J�O���Jk�[�����-8C^<:c���L�Qy���ӓeN4�A��P6��0���|�WE3T��(g{~�9#2�c����,�޶�K1�s�')S��\��GmoU\���48���z��4�d�^���No�ړ�!��,�<�|��6a�D
�R����F���C�k���ʸ�u6�ŭߍZzAU��٨J3���D�t+�����*(�K�a���bN���1��a����-�Цk���'uqN7���$w&����)MD���*n�XD��o3�@)��|��Ǔ��9*����Y��F>�G�vUDa��3�T=�UI�E�Ƕ����E!{g�h��|qޖ��!0].�hׯ��[�wp-],I�D맶!w���EA��Վ5�RY���w|�$L���	��0r��NT��`-�K��Y��Č���*<�iRI=Ss�hk��fX������U/�"\� l=�	�.�ZؚA�6٫~����k�n��[#o* �޿�'jU�C�n�4㝫z�XQjc��t9:g v��h�e}]�#�b<��~,n���V{-u�j>@A�E���m�mv˜��R~"_0���*�M?v������˺zb[��5Fڢ&�����b�h�a#�)�����`���@92�0�UOӻ�U��K�E�y/l���� JH�o���V�|�P���By�rS� �I}
Լ���7��Q9�����Y�w��$�w�x&.@5�g:�j���Y v&����^��^Ϊ�M���ㅣקΩR��l)�l#������n����^�j��-Ǝ�����JY���T���@q�M0}�<Y:V3郝x6�[�4�M�9��cJ�|�]2R*�T�A�}���9��9��<Md��؃Ty|:X6HN��,���9c����!���c��9�	�_c�+qmH5� j����"9+��;;	e��O�S�w�AG)�����𮾹;Wm��
,��~��jFB̺z_TѬLd&S�2�[�p�5tQD�2N��lٞ�,(7-�L�﬒���m���LhĀ:rvT�le�+B�u��D֦���j����6PD�w� %g����:��!9¾n��jf�� �œ�5���d�^�-��J�������(<U$��%��:�	j?�]ɭU��3R�q֛7�Oyu?з��(<�K��N�p���~ڈ �^��%��A�zL�`��'j�E5�9Yn�"%ݗ�,��RB����L���$/��=浄��my�3�0-�TB�� H�K�c�+٩Q�w�^�-V��,����v��#�-0�r&y��./U����0���䎽��H�K
����pc#�_mo������P�ǘ�=F��I�c	^�N�<�yB���$���݀���]甯����$>V��
#�Ԣ}��|ϳ���a�tC�K��C/D�@���Wv
7�f{�o��"�-��6�e�rG8�\�aq ��]�x�ӆ�#sZ����>�Ws�tjz�2]���C8�+2��]n�h� �;-?`s��S,�h���i����D�n�ev�����Cu�x�� @0���c�*�1�N�O�ur�w�����1̌;w�JS;������la�#�d)����q��׽�b��n't��U1�,  �����-i~h6��Gk~sOq���sA�&qZa�����<U����=Hr�'!(�{6�L�j�����"6���T�q���U'�6O��j��h\ z]D�;cy_�#�-{�n;�zd��[}uk+����7�����:2�2��Q������
%p��CT��w���B4 
��	�΁=n�m�	�n3M� �׷3m�2	��S!�N
��P 蜩#�h��1�{���\�{o�("b���v�ǘ�$���O� ����܆�G�.�Y���
�.G6MEl�����/sv�0�i��{����˂����� ��a��Y��m�����%��G2�1L��ތ�A�9,�0Sc}U��Z`���D�`����I�s��Ez��	�f=�J���Q�%RDu�T4�{D�O�K�űΌ%K��vO5| =	#/n�Q�Sv砾�z�<�'��9}����g,���㪔�����N+Hw�`�jf�6H��u�;��1;�/R (��ZuA�4��i�a)O5����f爐U� :v<�j�i�<r�mV��/G02����?]v�4#�Gx�v��f�g:�QT-����P�Gד.�4;�S"�z��\�f�T�Giٴ! �W:��Z��f�_��rq��n]�C5�����N��u���(_��5F,N�����ai�nC�������=�=i����w_a;}ꅕ����8��♻W�E�퇩���)� ���w��Z�
�١�a�6�+s��U:7?��G4�aN�n�"�M�� S��d�G!g���|H�6����ͯ���hn�W���S]|zq+�O��}�&M����U���+��ҝ2p)���k����c�ؕ����3x3��/,�Z9�
ݰG����k���@ȁ����C�j�,
p0g�7mɡKE|n4R����o	(A�~Irw�Q�s�J"� �a��5�灏�D*n�O4�����ʯ���wN���X��Ka
�*�Q��J*t�J�LvߠԈ8pDQ�Z�H�F=�$�i�Tic]��"^��طҿ�6�8a6����`�őa yb% BN7C�C]��ZYz�]�d�O�̬���G�/�[(�8P����CRI�ǲR��Te!	�<����`�J2E�0I�`]�� �Ua8����^aar��4N�~�Sn���0�����[�ga�Ջ�9.�-(�1�����o������D�D��^-��->�����h�ѐU�MG��O8|m�P�v�:��g��\$�����[;�C�Z�h�97�`��Ӷ�qO�.4m8��;�,�+��+2��zP�?ы~��f�!�Gdv�����jјc�/����h�:z�T�26���l�+��$��;���"���S^j�e<��D��^7���{� � s��}B��6E,�3'H3��\���E����5dQZa��2��AӧΣs�܅��R����H2{��w��R}zv���p|."o'���!�� -O�T��V�<L���L��=�<��G��阸���>��yF&���|�N�˒�,2ui��
:.���ȧ�b����ԋ�ծ+P^�+B�q��W(�'דif�{��by<}��k+�h��6����������9�F1�w=�n����;�ݢ�G#�?�Џ��.Q	�Š�����������(<҉������2�5�d���ğ�hyQ��Oy V2`�t5%���E��Yq�����/�}��s�L٥�r�B2R��b�?��u�[���׬�W��g�R	O�V��)z����s�g�A�$�)��r��(�>/�I�=� ��?��+RP5d�����)��e����]��w�n	��+��1:#�՞�z�ћ���Ypuˍ�7�K�o~����\��񔓟��/�}�랧�ǫR���bB"'�b��'�
{��ny���#0�m��#�	Z����:J��u�Ph�FL*�m w}F�~�1uMnXDe\��U_��$v^]�zf��ĳy�R���4�N�ï@(?Qz�):"#kq��͢��Ĥ��˨f�s茛T�K���m��UГK�)����g*s��|��c���*��q��=I�5 �Zm;u�V�<�=H���L�WOő��[ 4J쾰��g�����J�y�P��Yv�^�df4	������Њ2{�$��`�#2�� �O�܈GW|u�y궘�Cۈ�o���k;�nJP�YWh�7�IwV����x��Q�"�ew*L�b>�EYc@�s�'�k�Ɂ�<)�|T�X�CMǵ�&�����2�6l��K7R�_�� �Hvpj�� �g�J��<���|��w[�8��MhO�h^�ڥ�J�Mɬ��|m��&���Ø�#�hi�61�~�X��&���6�O���^��A��<1�{A=n��r�7�=5�����XO)r�Jf�Jb�Q{���\�@�x��_��
�JZ�e�^4������ N���4�\|��^�&e�ݐ�WK�Ob�|\� �4v8�G�mU�n�S�8��
gb|�A����C�-�����BT�" w�c��@a*�#�hЫ��Z�[蘿�ǟ���d��h	Gߓ$Ť
]�Bxf�S4g݅����� �l3�6��E�	�����r�	�vK:"\�_���Wy�U���7���\���_ f��!)�9��놤�Eǂ�"�|	��f2��@��prJ��Bt��D�^O$��!}Ƀ�A!��>lh)�1�9�xv��|̕(�1�W}�[5.�g���޻�`*k�,���W�� G��Jm>�!�N�Ŕ]Yଐ�!c��k�IT�2J˲E%fdCƤ*C�SM��]�QD�B����o������+)vՙ-P'���)�!����Gы��*En���tq��^��=B�����f�>���ꙸػ�hy����S��	(_����]��{��weڴ�	1��Q3E� %���2`�����r�_����1ޗ��`��N��ˤ��_`��c��ȇ"��[KU�I�Ay�4���&�Q�����F�r�gd�u�
+����W�se_�
��n�
���άc�>L}�<?�y�����:r5m�`��1�h�\5F���ǫ>=uu��F�O��~"�S����=�)2r���<��85�	��z�g��Չ>����G
9�L�)\l�fC�t��������~V��ױ��rP�!fNo��.3���~W�G��=�n��X�Z����&��_#ws+�S۩@5Y:"v��?���8DC�ʝd[M	MDKJ�}�S6.&-S�GS�{��jɗV��@��@'rO{��a+��O�'���j��<�[kǲB�PZ�e)�Q6���w�U���V�R�%�������_�D"����F�%�)8��g�A�>G�e�@��
T.c\Vm6�y �)OY#�Bkc�w	����ǃ�7QT�'�f�_#_A.%Y$UDWћ8�M0i7Pť�zZ�o���J�����#ߦ��=�I�h����>����q�QAJ:�^���3�=�7籜��wƜ5��Y:�90X�b?1�w7�[�N������o���43��}a�;Qc��@4�Ԑ�Q�z�t_�s�&�Ts��֍�ȁ��J,O�J�;���P�jLD@��CZ�O������k1ޭ���@!pm���Xʍ7[R��ް0���/�-�/wi���.�=�>�ZL=r^�$�pDh�kb?��ƌ�����(K_�06�٩��?��Y_܌����w$��]�>����8���I�0�$��yr�fX0�v""�g�2��w�)�R�/!�Ԇ���~��(T����8�w)g��|.q��MƘ4Q�,��+f��9���[d�m^D�d�t�b�?w���Fے��s3�a��Y?4F��?�����̤�*��W�c�P5g�۝K���ܙ����C�Z�=xM�Ł������.!h3�y��o.mf{����!�C5�aJ�;���A�U�tX���х��E���HcM󫮌�����}�.o�����d	-HX!.|x_C ��Vu����q��_�����=ɚ&%e���˷k�a��$�DV� 1�q�7�ť�UvBѸi�4m��7�_�p�����O~/ūN���?�;�\0��������������ؒ	@b�H��ͷ�UPزӧ���33���3���y��;s��;A�c��p�꜁M���1p��v�)k-���-<�Q�RJ�ſ����"��L&�ԘԹ&��fX�tO ��~�8�)��ɸT������ޔ!w%Q���ӂ�̧amh���vʅQ*�P��1��/(D\y\�"��%�qE�8't�FM�����gHp�i��G���c6["����@@��ӯY/�c��i�:Ɓ��x>kV�IL
�O/f׌�����'��~����Q����6�vH^po@��˦�!���3�m;��I����[8��aAq`˃w]��ɦ�����פƸt��cJ��¢$s��Rrux1����P��۫�
^L�����?;��o���v2�.�ۿ:�5o�(�翂}�ӓZ�?���1��������,X��R��ߧ��^.;�g�%�k�O��h�����������V���^Hb�\5��|�ѢU���Ln��΃^���9'�Zj����j��2�@E�8l�(���x� ��z˲|�e�T�s7��+wvRfcH�I��̷���l�s�PG\�#G!�+T@zޒ4��İ��3�S��|�?��Xf��_3{|A�>[U���g7z_^������h�1�X���5�b��h3-�;�i4�:�S�W�������[��*dtY��|@��4�$�<˗��U.L����`oivj��M�O�v�Z��^x�0fv��	mp�}��1�0��NxE<��<���S�Oئ�Z"�\���
E{s�W�H[9+�%�Q9��u-Z.�4��=��cS5zT*9�cJ$�=ͺ����=���K̬�������{���	���@K�	9���S�qi8��"�6� !.~

m��ŠQ��Ⱥ�����\;��ĥP�W�����r��xX��
�x_�y���7]�N��]`_�����)��y��ƈ� :JP]%�r����5tIΤ���쓗;h� ��ܘЕZ������ҹ0�e��M���v����z��(�NY,�^�_B���ٌ�x�t����ۺ�<�ň5�a�?L�ɗ&�z%���d�k;!�`t�Ը�F��.�&E�WoD�&\�|�k�%z!B�7Dr�z	f$�!���v���d�uH�PK{�&j��O�$�˨�ގ?t�-�U��6=��w��,0�c������0	�_�H���ec^�*��i?�%�2�Z���Pף�0��?�;���KK��{V�����z�s���F��9�nS�5�G�����b��(�B�k�ҡA�O��p��<�F��F9�O��A�������yrM�s1�m�8�#l׼���3�خ��0&�N"�0�}|�h����p��$֜�1�K�����у�*��\9CΦ�QG9��}t�ʾ�w�)��~�re"�-��u�a��կ�$DR�Fe}��>��L+v�w)���j	�̸L��M:Μ}+�N��������(��c邊��{[�~*}�Ouk��:�N���6*W�gq��J�=�@m���������(�~���f5Gj�0~4<>X�B����j�hj��_��X%�"u*U�ٚ8q���2��)ˡ��kQ���5��mֈ���48t�2ޱ?��:��b��wZ��:��m����e�hbc�߻.��FM�k�J�V�x�-��3b�h)��O�f��5�UР榩T����\�;47]e�b�܁:���g	��O��S���f㘦�$�ye	�㮍J`
��U���@I�'R,Cb��( p���}
|�#��/�!T78�O�����x���$s�}��$��!,����󼌏����.�;�+ѧ$���^�
��˻W�/(p1g��Y��4fl-J��N���QՎ4�n^��V��`@�m@"�%�{A�����V�7Ve����RP��7�)wCЛ����$j�zf&�1�)�K����×W5h3��ⳗKf�r��l��BJ�79K���x��۞���L����w�FȒ��7�s�GS��8 2g�g	�Yվ�AGч���M�Qd�c g!78�ׇG�m�7�!��<J$6w/w4fV/�ckBR4A���5�o&�<���4Y���05����D�Gz����?��DՀ�>}������\��kE�����1~������h�X�Ѹ�13�ڢ�N�p�NC�
ۭ�� ��ĠmS3A9��˸�.�z�:�pc�(|�ZB�K?�g-ŷ�g5�}�<a�;�+�ʭ�x�$B�1��x�Z!�RW���Ɏ*����9-�H�l5�C��<DUv0}�4/�ӣ�$*�)�tw+�u[�N�l_V.�<��[�t�)p��3U�2e�HpK��)��m������i}Q9����qX�Ӑ�Or�>�m�X��+�`��!�ߟȏ�产P���+ǚ=zw'��s`�aS�,,�}��xi �{��d9�xw����2��ٰ���a"|1�s���QB�D4Yz���o�v��a<��)�t�����ظ�hO��Q�}�� �8�֝�-�f�t��l�`��3�R
 |K)vkC|}���~«�J�-�75?�)"?�X"��<TR;Ф۠��Fy� �Z3@�G�[�9[X�m�����<��Bh{�I}@��y�}N�d������w������t���ڛ);��-�L j3k��צ ��K�Y�ł��"K�={K���6Wo��Iyz$�,ĳ�I��O3��d,^3d�"��KO%�o��i�����TS�qn�E
��a6h��t��`1���t�ݨAD�1+�Z��A;�w"��a��+�H��Y�%�Mm6-�(��R_L��h�F�>�tR�m]q}��_|#�|��Z#�Y���$*�{>H��O���=�w��	83,�R���y�EG\��~x�{�闬�c����Vw2�l{�Y�Uƶ?"{�]�[�|�kPj���rOH"�r���#y��YQ�g���}�O�D" �6����X�6{���%�O��u�Ex�c��P�w;&��JQ�� �ػ�9�쌝։A�ʹ��,ˤn������ų�p�u�����7X X�����(�	�t+D��>&��u�pϣ1�M���{y<��>�5�^IL�����O�N��wm�&���ub��3YZ&��nK(�6� L�9�����A?v~���;t	w�T��Wg�U�H�x�fȕ#Ƈ�&�!k�%3��<�oLwԒL��Sܒ����Ȁ����ӝP$俙.����m?ޭ�dC�H>�YM���*�M���~*��u2�PX_�Zx=8�x@��Aɾ�����`������juCM�}��ç�������e�<Am���0���<7.�3���bd@��+�0!=-� �,B×���"vJB�:"t7��20AFx��:2�du�'|��Z>?豲'����	�����O	�:V�:@?�{y5���r�.��dV��dG�"R���d�B�ͦ9'��B�|O�q�s}�nш�&�:��Q��&�`�S@i�������N[����ӓn'���y���2H�pN��2�*��ت6�t|N(��D{ܝ�<��!\
�T0.=��وNG%��]�d$�2�Nْ��8R����:�������b�窱��w�<B >��Kv���KAU��ϡ�SMߖ����t�d�#ʹ.�u��}�u:9$�k_��w�ٗ��m>�yI6�o{W�ǆ"�/�T�����8O�`���ƃ� :��yy�.�j���C��}42#�᾵�И�߉�z}���J���`;&���Hq�x�ֳ})�R�����1�l�q�lΧ"�{���#�U�ZC6���
�g:�`�x�%X��������;��3��~��m�f�O��V48qfz�P�Z�z��J��*�#�Q�T@q7��8�$�� ����CL����������r�vbFVid�X��_m;pVWk8�dvB1��?�?Zj�r1�±�[_t��k��N���%���8˪���/�E�pZw�C�i�x[}�N�lE��K���~�U�vܽ�0~�0��/;J����9%\��'��P�ȯ�5�Oi%{�Uci8��W��l�|ZK��j�Ϛ�[�p�-�9�8����S�*��%%6�[#���'��`�х�l�[@D"�I����s�c�VcY�M�SY�S&���G�kh�x���o �= \R�k��ؘ��һť���Ϳ��H�΋D�v�Ѭ�"E�I�r��S��6/黓���B��~��AKYtOc�M��
C��GL����إ�z��s��8-����ڐΗ7�L~����)�`����0�iӺ���
�[Pğ��`Ka:|�$X�L�
���S�٬���ο�Ʀ�O�������^����\��uK1M��=fN(L�ǫ��Ǹ�PzF���X�gbaOʲ̉O|Șf��qX�a���q(�T���pq%�o�;#�4����'��ܫ��e����:;sT�{e<�4�l��`#���S �`0p�<)T~�O������������&�ز�+�G��=���Q��I�B򒖳��*��}�2��>��Ⱥh�#��?��g4�~+ڱ��:�#7�@�m�����f����ly�Ʋ�w�B��U��,_��pY���!�f�w�(+^,0�;p$��A��K�ٍ��![���c��޷�2�Te�L���ŏaВe�զ,��QA���_[ht��˱�v�����ѯ�3ܫ�����`В�[�h�j
zٯ�>�x�1!%��˟|3:� ������tΎS��=#n�x呑�JX�=��I{��Ǵ�%f�x�f��W=GDe�аN Y?�MI�-3�R�OW�󌨩�I]C�ia=�A���4��h��<lU�f+�@��U��0X����
ʹ$Oo�*r,����w&��wD��GTC��7⮸hQG����젅�?I.��X���5�fx2��.6!`�A� �uM8�P��w\���r�]��t�6��@X�gn�i\�hh
�&�BG�6��<*>�l�}��hȽuO��8��3C�j�����B�혝h�0FZ��G�z4#���Y�%�i�3���|�J�����&S�04��L ���
�	����Ć=w��7��{:������8n�X%S]���3�'�P��lşw�e��8�R���z+TPp4F�j����U�uq��]��Cy��d^x�����9��<Õ��l���v Є̷x��Tzb�W��4v,�cDF�D;�A�	��iS&��RΎň�jk��1EL��:�	�3#��.��� A�rP�f��V�2�0�SOy.	:��+�=Q�����0b����Ls��;k�����P�/(;�4+
�+�j ���-X5�!�O
>8�ܪ��O]�����3$�(�y������f��J���s.�����ȟ���w���z��L�VZ͋�r=���u��e`�֨��h;`D�sj�yh�XEt�xt���CK�����R��b�VR�X����`�[�yT�_8�aw�w)�d��Hu���5�����H-,Ñ���*Ҷ3��l�/�	(V:Q%=�k��}�*��΄Ja�B[�>�m"�e���9��JU�����T�Qkf5t�N�Jx���Y/3��_�t}V�X=��U�N��Q���l�q�/1���F+�X�E��+�Ԭv��V"��7������H��0z�`��= �ʽ.���f3��L4��}�����,ł6@����a���r�A�B᩟i1'2�NN�16ƭ�iC�b%���_W69�9<o���V�DH��mq����n�T��Ԙ���m��Qf'F����l�,+�#f�f�{�7�dݛ��\��c��k����X�_�6��>R��/�+<�̶SDS�	�1�D��.?�
���02nS�	CN��f�wó۽�{�>׽#��,e�D�C;�~ޥ힂���s˛a�dGL�����4zJܯ�;c��4F�c�!���\<��Y���Q�p����ď��8���:nB߂�"E+!3o�R޷,�
|0�o�dBHS�J�Qz�������d�+��+���
���[�C�6H�k�j[D��۟ϔ��F'����!���8{Jj������H�Ȉ���d�w ��0����*C�yA��ͤ�o�޷�]��e\1�
JBH�]H��6/J�6p��r.y����9 �a�)�����Z����]��T��ޙt�>��78��#v{�p��+V��J@z' p�&0���v��%B���9���nWw�E����L����B��D����O�\촞���Q����P>-s��a��%�$��B:�_�pP1��֡���#*�*�l��1$"�#v�7�	S�t)�q�2�£.�\�@9]4���y]�Յ��Y/I�e�$7����SB��Q	����z�� Kߤh��hO�}6B�e�g����#DJ��8Î��P�12	*�RS���S	�q��H|�'�ؠHp��Ky{O������O�{Y�~�o�β1�H5�smG��rA_c!"V��U��lR���xY�^ ����*4�]���f�9O?��M��aCL	�"�U3t�9�FB�Oq�!�0���9�k�+8J�Q����~�X�	Y�3t���{K�pQ4\J5ޙ�)t�//J�����4��A� ���mK�Vt�S��z�B+��/���zr�ϥ���u��&/�lP&� �C���+�|Y�G�fL��c�C�>VbjcE	�vx)��i��o�}X�����L���F�LIu� gu�#0���\W%�`�j�;Asf|6��df9��Փg����\�B�ثe����N�eL����}�*��@���F�?}��N}���32.�/l*y`#����T���.�@`�x ������q� �p�{���f�����h�E���x���4B�@�2%T��!��J�)�\W#�Kh�Ee���{��]�ZF�v��r��n}`��;?/�9�v���ҫv�m�ha�y/�̈�)�#%jX[i�~� 0��g��11 �!��W �w��=����_�H^�e*\&�&�u�z���O\���g%[��,���6�vfO;���VX���%y�W;:�f����0��.R��2i���m �X�N��*�"ܘ�W��OL���6��p᮵������a�c�B,�$9�zQ���6��Y������<��a".���M�gi��d����*��3��짫�q7:��tU�������m~ȣ�s���$��՟�����P6�"Íaϥ�r�4g����[i8����Y6�'YO����W�eEB*ub��^�}B��+�� Ʃ�vW���~�gc�"��Y�-�ᓻH�}Uh~
�_�ߒѼ�_���[?�� ����@���.e�U��|Z�!L��$'��Z�[e�?�ўĲhpW�!���_Eb >A�e�1*�~�-�	#�����_��p�Z����*}�i�0�H����8#�7���~!  )�P��+8�n#.�,��TB��l��t�ԫׁ��,��g�~���ޜ�P9f9S!� ��O��K���č���'Мe,Sm���!2��)��rO��в����)ՋS��j�Y�������@fXl�o�i�O�ծ���B�̎]N�x;ψ���JU���]g���q��.MH��ٞYI��q����7'%sHˋv%��XT�8�@���g զe�y7��6�9i��`��J<�_�՞��q�P[��N]Qo�FI3Ѵ�ܛo�'�u�jtZ�g���NQ �M��Q�F����&��tE��RBPO��~����z�/�n3A��j,� ��^�"���yleçu`�}���J[�D8����2�N�!��(>V6/����GI�ΰM����{Ǧ�L��_B:�j�[��g4�1���L��8$;���lU*�x~c�0�i��(�,�S�X��)[n����} �g4\�UǴ"�����~#]Mp{cwƨxY���jq��)CT��ԱOB$@f)�,��?B��r�<�y߬x8>�hMzE�����x�z�(	ٖ�B�ɤi~8�o��.ǻ���OK�DnF��*1\ ���e�_��^��
�~���"��6z�6aW�ö�mz!��G}��MV�s��>���S�Ҟ;����,7�mM�[c���8B�dM?]YN�<�Q>�ջ�`����n`�p�3�L�\	:�V�s[>>kyvާf ��зO����1�i��`��MKfW��
�8��]��3p�(~=n,�޻'����=&F%Y���3�1�c��:i�G�ɔ�ڐCaeWRu�&���i\��R��V�J�q��b���% �&�F	)|�sa�6����7$�p�~&�gv�C2쪁.�x2'!�T�E�A�]́#Lu��(�g�6�<?^#���㹔�IWYo�(U��������	��]���}�j*��ߧ�	Mf1}���xoP}lHs&R�J�W�R-�=�6k�����ZO9�mn��{�I�/��{�6Z��wўɔݭ�v]�/+7�f���.��@!s"�\&!�:��6��ش}h"�'���X��e�`�X���R�	�t�8�ϙ�\o��Κ����/$����q��-&��n��X������� WK~����ޜ�V5��.)A-���0L[[ ���Ug �b��aϵ\X�1�[�h� %u9��}�g% %%���Ӌ��8�`R���22��&���ND�ө<΁m�w��#A%cm�!|����/��WjiC��+�V�"�ĸ?�QJS��~�(#`��l�o	$���,�)EG�KֹԊ{�?��T�-���E�H��+g��:��\_er��� K��`5�Gq`#(+�Nr(z��GtO�<ء�u�R�&�6�w����2-��UR�db�
*�=^�D� ��q�YZ|2����# ��v׀c����Hd�Z��K�z��:U����~R�a���C��Mie���c �w=�����.�	H��JQS=���ǕF/!�.i���Z�c.G��l�>Ҁ���"B�eǧ��s5W�����a`�A�uA�F��g�� ���߁����3�F�����������X�ܰf�6��l�N�����xK
x������hH~���\��͠4�j취'�"W���Ը蛾;~�e��M�<e��9-]��:]۵�r�����h��2�(�)�m\��2�2u��䂣������sH�=����Gj���#N����Z�<�CTw|k��_S�*���,3Y0w�pǼ���y�'�GEETnY���+5{����ي:<��x5/p<�ȁa�=�Έɪՠ��l6Ò�J>J��O򿘊~��{:+"4�^�R��Ųr���W���Z�7����8��|�b�|ez�z�}ȕ:��tf��M�>~���g�e%)�k1!��4����}�L'��5�!�.�##g�K�T;q�=�Y���72[�<e�FPZŹIۯ�涇���5.m��0�';w`�����**�N�k���9[%�(�����wXL��d�{iJ���&a��)��G��$�� H�Y��~�}�
ڼ�E�uo����mD�lF��TFo}]]���hVNkݷ
�c����'�O^"���MBH��B�H��)G��k⶗���tr_t3Km��ݤ$-����]w��=��j	<��mI��Վ�G�I~{���]�;��hXC�!�v�%��/$�k��0\yK�p��^vrVw8
�����+J��r�����]ؠ���~���g�(tP�0m2џ2i��
=x�Z��6�J�;���鼉� 
��B��	�����}�
������cĩ>��:h?f~V|��ԏ���%����v�X7��B)b���5U��p,��fMC�.7#OV䊸�4����jGI
�P��������+�{C�N�!Fn�:�f�-=�r��X��&]<q��V���'���텺�zϮ޴G\�̓"m}�G��Y�6=�A[=����2�2��&N�؁�?^���=&�i�N���z: ���~�2D��᫙W˖������3���ۋ�ĳ�n��,S�� 8�ٺ.u1�8t@�� ȓ�(vڷv'�5�A��,>J�]Ӯ�~F)����4 �rP���O�c�9��9�ns� *K�j;u��~R]^jkK�˼�n5{!Y�dO�bf��D`r��(��c	�	��l�����ma~'�c�M�w�A0�g8��B�b��rSu����k1!��do�I2�R�<���U��t� ѡ�ih"��V��<���W-L��{m0j��~��[[��s�һ~JHEY�w�f�M2"�12y�XׯnDk���������b�q�����J&�3{=�~MSm�cK�Y��,A��X;�L�ü�ұd1����Y��L����/̱"6X�����۸iz)�^�S����0	��i�1b��A���6�;U��Է�Φ.�6�B'�팱�*o��O�h�v�5�,�%7c��hN��	�߯�B��{�떔��A��Ĉd�p2,��ʝ��p�I�Xɐ��b�O�����M����VT(���k�BN|&r}���O�ũ�?*���r���#�/9؊ ��T�`��}��Cg�܋�M� 	h�º)l\p�OߑFd�$,����@e�.�i��)cT��.�Ά�`�E��:.Tj�ǜ6��3��h�a��R�T��s�a0iWjs�10˺�(i��n�������9��߶���!"��Q�]���;?�˗_~$N2���%<�܉0��pW�����j��c�$xN{7�4\sv#��F]�(�t��z���&�W�:��?����ao;�i0�Ӎ���vM�:�k��g3cm(%C��/0.�l�V�<z,������A��d���n�m�Y=�_'$9ٛ@�ng�)�q>�Pu����&M#�Mw��E�������o���h7%T�'9a�>�R!Z,��æ3q�1'��p�!�w>ۺ�ǃ�e"�fu���Wd[ÖC�Ʈ5Wׅ9�[;l'����rh��^�̿���
L(��i��&��`$����?�~�W�i������b�#��p�N��F����O��sq�<.�%rMna�F `�а�c-�gx	t"#a!�_�54~W�����i�wQT���DT����'��H01��Z��0��:�
/�	��B��r�Cg<��J�"�]��[�O}����u���VU�l��a���9�H$8�=�҂�ے��{uX��re �N ��;��#������X�%xF+���Qj�!��F�+S⯛�@����/~�J얬�O�`w��mqC�cX�W�D�VS����-�8��D�gω2V�MAZ([����5���ಕ^Q�����z�o���HDƾ��x���aC�"�c������%3�Ӵ�����Tk�5��i�Ò^��9�GC�鞊&fX���b1�լ��?��5)ٲR�1u�_]�_��g�\���ާ���=��NC6`�7���s�O��67Da�5�49k���We+`	e1��4C6=XhKb>9�V�0Ӿ���{�J��v���w�b���+�s}V��hێ�2X�v�Կ>�r��O�ޝ�zy��`���<�?ݑY�y��$��թQ0rh�aG�<ǚ��d��W2�8��*��Ő�a��l�6.ww��F��|�����t\��S"hw�	ճ|ѽ�(�n���f?� �4�͚�9�1�N�k%fb(#ܢ������ആ�	ẃS��vϫha�N�G�ωߪ�^ߥ�aa�W��|"��k�B����򯲖ɻ����`�6� 
BJT��U:+U�\�.�.�9x �o���޵�g\W�%!hZ��)��������p���G.үjK.��+�!�X
�/���ņ:O-������u���F�)Q.H3"��E���	q�	����I<o�;L1�t�<�v�]�+K���w	�$�u�a�ʯ7$�BW�pV�E�8�w���Xh�4�k��<d(F�|��dЋE���)K_5��ȿy3Nv��z>&�3��qN]�������bH���BB"P�����fE�#�%	�)�/��A3��2��VX��˴�M���j���bҿ�է���T����]�|����/A���
E����A�^ۨ���uj�̝i()��q�Վݺ�����E�h��Q (��uF�����/�D+�v�]6R��*ƕ�l+�皀��=�/U�羇��t��kTXU͌oW|��(q��)��"��Q���y��άԝ͞Hej� 4P�7x��I\2}�� \/�\�lN0��x�z�,|��Х�ƫG[y>�|�r��*�G,�h:��<3���r�V�ܮ�X������J�5[k%��4N�Y+'��䂚�Aͧ6��q�f�����ݥ�X�Xx^�<����>x2��1T�O��W�H������1O��Mwv���9йN!&
�s��g�����Z�������>�N�fƓi�M�����|Էo�J��D#k{�G���D��J�-@H'1f���>�벪7���Q�t��_�����[ڪ�0r8P��d��R���2�:�kK�"4��g{�,_���W���9�=s�n�9� ���g�k�9��R8(�76ޕ�缵�I�3�ܩ�z�J(J"6�-���?���c3�Z��b���Y�yt3�g��b��=�m�4���w�	��{���T'��9��=�3�,<���� 0��ǀ"�|����Gn���Hw0�]�E�ɰ9u�%-��b�ܵ=]X�j>���i ���l�v��^ld7~�*:5�Bg�����B$�t,�a(uMAB?��c����G��/�>Qezv�f�z����"5������ZF)�"?�V,Kk6[X6��]�.�Z��Zj���y���Dr�ř✓�J��HR��@3p	EO�F�L���r�������Q��Q�o��C<|�}o1���ҏU9I3���{2蔖�Ur9��=��c���6�m�X���uIYJ��� �f��d���u�G��:8���P�qGm�@�x(�&�ۥ}������̥�r��f�ɦ~��c�'������$Y�<WA�!�[GR7a�J'C��c}pT{�h�0�����ސP��U�."���3HY�҇O��)������<9���5�K뮐��x�Ɗf�L�b�ھ�W8O¼��
>��p�U}�>�ԍ��,��]W
<n�l��H����{��{�=���Z�ʠs�>{��j2�8בY$8>D�3�$�$�D�b7a��ˬW�P��#��,e�����U�9>x8�D8�bm�N�	H`�/� ��zݗK`S�oN���ԩ�� E�G��+���y��ל���a������p2\q����7���yy	�ho�5���M�-�Ⱥ`�kj�FfhJ�R�I���N��8 uZ�,쬜OE ~���j�0������9�-�@0n�O	h����l�;��Y�B0��W���N>���	<�Iɰ�_��s�$�5��g,�ƍK�9p�T����,�����O���j^�o�s�KlAh��h6�ɵ(�������9�|<;n� ,��w@�$���&��>��%1˒ࠉZ�KA��x#� ۮ�j�'Ǐ�Hԏ=0?G�������Kϯ9�,�X��2a���=�ɋk�]��Ӊ+���#��3�S��[;-T۬z�
 @VWp�����E��ϲ5.�M��LT�ŠG�����բ����'�&���M���ot�HD��up�gW��8�����iH��u�T�uf���������B��l�A���̤�~��|�B�n��μLP�g\�,4��rf��,�|�.���G��ӊ��б�doϚ�:em�Ao��a�����Q,��-�s{Q~a���%\���}2�{}�U���Xj���������
�_~d~�u���YTm�����±�֣Im�glޞE�Ι�{���c9"�����7oU͌`���O�s��T�V�� �He�,�K�2���y�{���9e|_ݮ����vA���]�[��� �6�K�~:�Ө ƯedΕ��<dn�J��*m$d_��"b��~zƙ
ٚI.Z	:�+�3I�nUM��j��b��KW43W�v&�[<V/��oa;`�Q,%8lɸ��*<Kt�-�Ij��,�NA��� /��ԅ�A����.��,�EW�������0O�Ӷ�	�8��T$�����5r;x�;�s����#y!
�H�G���jP�*�f�3sc���6����[ĳ��`"�2�J�	��zY�0u�|�UV�����Ӑ1>�q�;M��(+��t������a�:� ��d_', `��w6+��mWM���mL�TX�F-�J�����*�=�c`�����+�!x$��G�H;j��?{q��g'!��_� ��z�|�ץ�`��3�7��B��ŷ; W���^TV�ٻ�
�����읇�E��F=ry�� �V��ʚ���^s��z����	�䝷�t�R��o��y�~�E���	B{��Ԙ��;���|���
~d���������a:���:5���H	�h*��å�S� KD�>F4R���l�t�������K�ZM�|t�|���E��)u,As�Ҫz�����'�p��`OF�n�>(�7�|��N<�	�� ������C�g�u���cR/F����ŷC��
AY��m��?b�'/��5���Ѕ�y��.�j���wa=��{�=��jw������i�	�v0"K^y_"���Q�Qh���;yܭw&A���͊���!��$H]����0k6Z������ϸ�;�cee���Խ��T�V�a���ݹ�e#����pYp�ux]���,J0[�7�q����m��Q߶��wU�tˉ̢N@ϰpҜǒ�V|X$�����nS�ib.�k@�!����<��a��نZ�dv	����V�Q�V��^�$����"�^+Ę��������+=xؒ뮥�I�g>ʑ��jξ��͹��{s����ݳK�e���� 6����F#r�=�.�j�����!%$�*Q{)O�q���
���?�6pk@��N'�Џ���n�ɹ��ǡ{��%97T�2���02|�I�~u�
Wp���T��7MY�P7����t+�e��L���x�W��~�;z�]wM��#�w�|36����h�&�� �|g�"_�1l@� e�?gJ�N5
��F�df��+��^�u�S(�֗�<A�YN�֟�����[_?�K�Œs��K��O_ �>G5W߳ ���>>�FTcq����guS���WǊUXu宭!��j���0z9����/ �y����y����m{��i U,�筼\͎?��p���p��<ѽi>���s��B�\q��'�Fs��Qa��LQ�l/�#�R�� ���qn�=��*Y��뭙�?�qbTdx��NYސ��ƍZ.o�S$��#��|ǯ�1K����7o�V���ޝA�[@RF��v��l���z�'G���a� =���{ii�*2z�H�t>+jF��UjϦ��c��{�W�����o}�Or@F5���A>��#���L�z�Q�Pᆶ")��i��N;�ɶ�?ґ����Ŀ�JcͨY�9���Oy���M��|⓫��t�x���Y
����5�fo�UT������ i�UM��Y��%�Wbd'\���o�;��O�;��h_!��݇e�Hu=���@ӧ�.���Zz��5��Z�h� ۨ�ֆ|4�	�uP��:a�]|��n�����c'%߉�>�Hx�
���x�^i���J��!�qZRv�<\)�b�w���!�
y�@UF��V�^&H��{��a.0Ӽ�&�#a����N�XN�,����`{;�D�=�|hb�K�b|E�Dx��+��V%���4��~��ʾ�)N�	K���M�s�ʐ���5͡��R��g�ͨ�ԺGj���j\���k��%���*��4�NsDb9�� {��4��ٛ�Q?��L!�:�����2ThޱUP��
��ް#�F��Q�`���jW�8G����>_�?2v��A�t/�-&�n�z\��n�|���i:	qFSc5G�6�`�H�vpI�En{��q\��s���'q@_�,�!��b�3�ˇ��2X]�թ��;;P���G�V����rFt�7��(���!�9���q��U�?�e�*�#5��XH���d+k*p�sg>G�;�Xs �0@�4���>Je3�*��F���}Y�8�q�ʭD	�J�]��C��l��m�����X-w�`��A�nj��uG3Eꐐ^lؤQ��i%e�?s�k�pF�&-1#-� t`���W@ń��8��L�]�T������û�罹1fFin�@�@�C:!��=
;V��U�G;�4���?��\|f�����#S��o �/�Aq>n1�ѷ3Ue����a*N���)��,(;��ZzS��K�j%Z{�d��@J�����Kve�ݭ&�^�}o:��+VzԹ	�Z�S���ūd��2{	�����yNӽ�B>�T������s�ͭ�qRC���@��Q�VCew�A�Jq��˺L��~�>���?0��\<�/���X�'�T��`�z�F� }��'z��ĉu���2�T#޼^���9��㔣v6��5|�Z�{k�P�g ]�ը6��3:��4|d�7���"�|�6{�+��E�z�u�"az�s�1���^tu�����!��)al�l�Yx�}:OĖ��&�`R[�(��(�N8끗{xTX�t�����N���y�ѐ������	, Cׅ��qS+�	{+�x2%+O�ڙ���VƠ����*&�H��VJU��Aw�4��|7!�_I_����}.Ş��OT��ʳ�j�˾��Y�P��~ܶ��;A_��UY����}͛���!�SB��׉�[�v���K4vq\����i�ס�3��YU�rq��v�o#�iʒ0��u`�� �
�o�W.x<V��T�/rm4�H�}�#���X6֖��8;,�ڎH4�4�Z���~v��s_*sD��5+X �����������b~�E�����[a��!����s�~c,E؀�M�Y�|��#&R!+�Ľ�Y��8��x�%�
PtF�9	}��D3WS9��z���e�R� ��"���%Φ'�� �6�"Uv�Ʋ�?��܃�m0/)n����V������wq�� %�++vR?�jC��)1	0v%pAچ"���>�QԿ��!�]�O��}���~h�>�f��i����2��C��2�C�����h̫GD��}H�g�o�'C�~�(�w8���j|�"�=Գ�����!��1*��_`�߲�?��pF�H�z��ik�9˗��8��`ҚF�ks�~�d~I�D�6)�x���7�UP�WP�����A�7u��=*���rD��(�g�Aā]�-�z~�	ك�J(�YV`�y?}� 9�N��b��o���Òg��L��%��K�|P
�\��A@���i��w#<`)���'�N�<}D�)�r��#�����sm��,ƭ�Lvvp��2�f���i�~\�p�x��_�ԗHl'1���l*!�~�1��*�d�-c��;��qGx0�Y�9�qQ��?��!��s�2�����|�^��H�����cz��OkCC�;�Ɇ��x�f� �Ws,��s����R��ƚ>���&�;�SU�M'GGC���1wi�7��M8S�H@�ݩƥ�G�}N�	�r��AK�RtW���>@.Q�޷T���"�~�G9^�8���k���,��5:!�g��{����[�4�
�E.�<R��V�(����_p�[�S,�?�I��d�$Kw8���z~�>)�Cl��{,��E��3ϱ���=����=�
��bv�]���S���.���Wo�?n�\��̽�
������b�	�0oxs���8G |<Ү��
� �@��.q�T�\�H�'p�Gy�쾰��:�.��O�~��� ��S'�C&Fq;!�g�ˑH�ͨPTz�������o,5ȍ�$X��j��꩟�q�j��K�G�ηW(�൴�9�����I���X��Q��&��<x�Bd�!VY���_M\1bn�BI�:�~t�~�R���_�L�B�|�k���4��-�|����>���K߅�d3MtgLe��?�m��g��I�7ttW~�f8�3�A+�]G�����]�ُ##��׳�u\M�+º�� xUՀ쓁�����2c��֜�}U R�Ӣ��5'��i<X�1^�#���ב��T��,�R;�nyBk�C>A|}zsd+�['1���ǽ�'b����	<��`�[h����6x����U�NSW����p�M�W���f���%��ƜC�d�Ǖ�l�Y�-:�4��wYi�s�`̕����/���A�������I��Fb�I�|�X/�^`\,[���d�X�m�3x�nCț����mr4y�ƞ�@)���1���Nv���7���o',�N���hE��+�L���L��/�z��Eπ��)�S�����d"h��&z+z���������'��=�DV�9w�آ��]���`1��o<c����~���8�Xu$l�������MR@���e����Ħ<�j����ߩYY�}TLE���v���� Qj-
����.��������uC�p�;������9L�����[42	��6
���=)#�tޓ�R��&+ٝL���1�pe���)��G�3�l��\u��9�|V-�tH̔g��Ak��n�9	���&�v
K
�˧#��L���b�W٭]��1�AF����=X�?u&%"Gw��=����T���.~�|60�|���!N�����qH�/���35/�E��^6ZN?�g�^Q�s�B3T#޺���n�)��ռ�w�J���Ьߌ�\�1q�Wɮ�<v.�X*�dil��}{S+"�6
�@Q'�pj�:��gfO`Fi!��~H�ᝈ��,���?Ӟ\Zq��sY�*f���$x�R+83l�k��(aE��y��Hw��j��/�� ��m�"L�''�������ȅ����M`*�˪CvՓ(���l?��f�.ݓ�5{O�����wX��9pb��T$����P?eP��NG|#��0�u��L�&:�v�F��������1}(�jy�GF�~�����\(���k���#�A&^Vz�"�ʣ�-�*���e���Ɔ}��Iܗ����a���>[Ҟ�I1d�V `�L�H��Cd�ւ�Z_v��89R�E�M'��j+�M<q齷��s�,��4��������@�N2���B��n�8d[���}}��hm�>��������7� ka�J6�v�,w�`�>.9l@^d\�j��خ�`
yH\�:hk-̓
 }M`�_��bIב�j���f���Ѣ�t�h�%�H���?(Z�+\ټ�_���fn`��ֺ������v��:��(�lo<8�>0�SP��oSbl��c&7!�<z�7��o^PQE�Zx7"_���?}�,WZ��{���\�b����];�4�3˝֙�cx<ͷcg{�ZRȍ�؞q��ӀuL�%�� )�2���k:Cs��ǼJE#�_��S�O��}M��L�̛�^wy&.��{էb���ĝ� ��YӘ\m��ҡ�m;�B01�Z$<{U��xaM��O>�8�Y�M"<�{ow<+��L��Z�eiA&+�&���;i�p�(".��5M�7��L�Vb��d��O�ظ�Җ��NI�i<g��eA�̾�̬��驛-��>Pnξ �c#���u �=>Y;��)��s4p�~�+��!�-�;�7,�)m�WxC���.��d"��v}*���#�IP�PR��UZ����D%�"y^jv����Տy���i{h���t�E��x��v���K�=��y�WÅh���2�R�D�+s��:�!n]��G��Q��Sf��j`�������~D=�^����AϹ�Em�@U�ZSp,=�ɒ�"C-��(+@I���ʵV��Az_e��mRy!��;S������7���
"����, ��琋�s��3��4�_�2���ghW/7l	U�M�H�\�׋z2�3Wz!�GN�e���^0l�V&w�{BM��q�s����{�mk���}��7u����jh�С_=���|ȿ�`@��S��=ɚ- �_�z����&gg�=ϤL��c�N=(���3tJu��V�
�����@8-Ȧq
\�Z\����c�F@1���O���j{��ܦ���PB���C�w%��GӲgCC�j������7C������rOtT�@WS�n'څv�O�~D��,��A�Ü c��tۚӼ�s��J�!���+ u���f�݁ ���X�ܶ�����@�{VaW3Hy�#�N�����*Xg�ƻ҅I��Ӛ�b�{`P�d�IA��^�>��&lbI=Mlbq�e���P���Lv̱Lcj�ҥ������*Sd��+�N��tٳ������!��닗0��R�ac�����E�L/	�C�Z#oڶk�����ڃi	 �C�,pFR��.DY�8�4�N%��/��Y��Ώ�!����4g�ls�s�mg��^�<����qF���Y�˦������:�;��ql��r'E;H���V�o[J�'?�Z�R�pyC��)-��~���Kv��Õ�Ʀ�XNt`�]~��`	���/���=߮��� p�b�C�
�Ɨ=�}<�:�~�a3�3�b�3Ɠ"��V�����������ȇ��5e���K�ր\�f�eN��q�4,kuc����A�?L�5Zښ�C}�g���,� ��t���T$`/WI��}F�\��}|�g�~1�Dؾ�Rp�!lR0�;A��jZ6����-���s�1	y꬚����Ҧâ�b�`�YN��ܲ�g��R��-�wBG܊f]?�U��u��V9����'��a$��2u�(�sQ�+��/�F�����^Twn��/��&�U�1��ϯt���z/���������iO�Ұ�6����tRW�|�3%_ZхJ����9S�Y�:��K6��O�>`�EG�l�C��:<���C�A6�u6����������7Ҷ2-Hg� ��!��}҇���1KRt:$S)���Y��F	��x���`?V�\y(������9i�C���5J�T�̊gʦ"(n��Z��E�!�+e���q�
��884=w�
Y������W,�1ɤ�ީ��<�qN���q0��(��VNv#��1��J��Vy�)���u�j��ԹrR����9q^������bc'�d�,̘CJ�S��H�1�����#��P�d;}�ޫ��m��UAH��ͮ�z�*��xWH:�<R��!�ēY������R��g�'��sY��Q�|��{;5Q�~�rq�Q�/�:f�G�몘}��w�3�Dbh�SQ9;�_f\�y����!�R������*6 �TB�>߿[�BmZ�θ�М���B�>2���F�	����Lը��0u,*0~DiF��4����v��e,s���-�㪀�}��X>��]��^s�(f\ڳ��X'�.�Xwm"������v�ߍە�M?������\Gsv�yx�2p��f�f��>e>�Y0���I�,��:WD�5���D�t��>�V�_s�{A�-�WoTt��!|�j��ls�~��e�E_r.-�����e�E����`W{������N�
���`CPX0�D��;����z�&v8C��|��V��8)���(�|��ђ��0 ��˯��U�D�F��_�p ��:�?��ls#7�:�����6:�ON*p�?f���cm�k�����w免��3�2M��6r�S��o\u��I���+٨Yh�]����w?��1�G����F:�<b��/��	���9�����9�����:z�h�|e?���I�!�eَ7�D�ĩ�qo�t�|rj���U:S��Q�`��E� X��A�NX�G&���X(�*B���h��{>+�M�2��+����{z$��$~N��\(��eäv���>i�NC�<}�4��?�C�������q��+K�+�T��Z>(ѐb	��Js�m��v��u�|��C�5����&"!6~R��g,�n�������KӨ?V-�h�^�tr���.�2F{`qy~=���7D��Tt��<{=�+fX��5��I3$,ܜ����dJ�%Sj��L�\7~��}�wl+�d9�	�$�!*K�z��� H�L:zc��'�7���*��(CJJ�G��#ӂ-�4¾��K�~x|���Q�6�������m1��+A
N��s ��m�ɩ��淛r�F"�_�����:�Pp��(2oZt^Ʉ�E�b�� ,ޤZ�����j��\�
�k��伀��Y�s�}��~x-4�����BV5o#0�X(5�$�ׂ���Q*TU�'{m�HT;zX�������x����� �]Y�Ľ�C.c�b;wZ����D�<<�9(�.6ȡ�PT�}ȣK��wҥ������&."n�g:?�ƃ�b�ɵkW�� A������/[���)a����<0���d;cH���5�5��nTƇ��*ⶔ�N{3� n?)> /��4�6Hڛ[g%pQ1&�?i��7�%��K�J��J]�� [���21{�yE&i���H��j�O	�F��'�E8�O��5U��	(�u����7��Jf�7-���@P[ћG�4�дʿ�ը����!֕@=�t~�yN��su����'2˻&�h�)��.�9
��lz�<ed�?[���0)��e�UBx8�=�H��/��$A�b.���|�kjԕ���c|46U{�̲_��Up�����$�k��+\��r��fA����g*��u8��g�ؼ����,��e�!����cSMun��h[<V\U�Ϙiؕ�[��T��h+i�C����R�Wg(��Ŕ���k� ��,��>�olbs@�\4�8�?,
�1t�X�.��y/�޶xl*�-ъ�<щ�G[�e^�$� �7�ž��漦�7�A�4���Z��I���J���F(&(��L��ڝ<��>��4���N�< �䏫���M��L��|6'aO�Nԋ����p p�(��H\�ى<:��P=_p�����)SL�l*�8:�-�>ZT����Di%��6�v.M�Z|�i����r����.w��f1�j�[�7��y(2�;8H��Ժq�����/̻��1w@}�@Ǣ��Ѹ��_Az�'�3�몪�3�<���&g�R>m� [�[k�y��2pdzP#:b��V�<�ٜ��~���N���l�����^����i�J{ ���nK0'����Ұ4����I����*�|v��=�/?��Rhw�K���1�u�p�%�W�_��ګ�?[�sE^Nv�V&G��� ��
�1�n�2�ʵu?�Pw�fi������{�����a}�V�' FQ��+��A-�W���5D�-�fM����=݇vbBh�;��=�\�e�(o��:P����:˷/�PĐO���j�mJ�"xs��`)�;:�֫Z�=b�<S�/n�o��e�NѰvf�Jb�6[��4?�����.v��L����5����ACǷ�cC��j	w��w�ŝlTX / 4��A!k!Z5�R�W����Ұ��q�֊���50Bqav��"�c�
d�����F���-��s=���b;z�I�����7�/@�N
zS&��w"����)�����aZ� �أ����>$Sµ�'#6���/'��_:6!�Vk����U��� �kCJi���`9h���jz�8��"�����Tߴ�Ց�BF����n��������4�bL���}۞�?�<!�jn���J����{$��b� R���z�$u�������Nx-���*�����S�r\���O`Q]�0"WM|@c��3�P�*��u�e4.��o$C�롉�q<� ��on�2�
%�	��}��}�u�y
u���
Y��g�(YoQ�*��sN�h˫,�Kv��{�� ���O���q�^�s^���
ȖT,�OA�Z�ƽd0���J���_}��u/l�ӟ�޳�U�-ѲB�`(��L-�+R���cG�K�/�i<�S!�T�����ݿi�{����v����P��ن0�ςe13]Z��H�zz
�1@�ۧ��������Qt�A��۩��l��}j}l��4(X��*��,�Ȅh��n"���ӆ���qkE�������.ӱ�Zm����I�����P�p;?0@&�:U����Hɾ�D�1�sK�W�M�;ghf�����f.�l�b.rd��>�Q�IeS�
�:	}c~�;��N�wL���x�e��>'��{ �"|T]J2�K �cH�[�'��r,$7�|��F��0���������M~���o|� X�f�h��
�G}#��qe�e���BSi̙�`�d�X�ŝ���O2� U�W��w<�{�p�2��͡�$��L�K`w��My��)3�ש�-3>�i�b"}��P�x�0�D�S�������,�r�����隤j^�z���Y9ԢK���5�q_����c�s#������,�����,H�e�J�LB,��8��1�FI�4�Le>p���O;�}�ݝ֦�"&�N�3n4 ������-|۹��p���-��!�;w�U���.)"Dh��@V���lG�=[�MHa�n�/�����;~֮���r�G����o��rhH�%��%ؔ���[ߓ���u7��=�jI*�B��fT�f����&r���][����5���^g[X�%�Òü,Ld�E�PG�E��R�L�6�'}���:�v�	����nL�ǌ���y<�\�Mܿ���)5~��M|�=��XSr�퇳��F����Wߙ̓k^�9����͔� *�FAZ����]U�ff���#��oJIWPh,��*���<w��|��(=e��NN�-�m�+4Ă���	�3?~o*�0-���w0�+�e,��C5H����
涭��
���Ep�o1�$\�[��d'�����*I�ѷfc%��먆�y�t`��][Y��G�K�0�^9�ҫ�F����p������7$�(��;��3�H1�ݯ��N�@݃'��ao����u:pKϲ�u���&����:Ez��t��'i&����]��1��%�K��6Kwm͠Cv�?&��9ڟ��0-�	�-�Rro�-ђ�n^aQFN�(O-â�Oa������.��?�"*'H�f�a�S��bğ���\�d��QFS�5s�\�#V����)d�~W��`N6MNO-����.R�c9a�>E[��(*�`���H�t�:���_ "��m���1��!�p쇕���Oy��~6{l��9k��H[kCV2H�����&/2=5��~X�[^`B߁	2�������+ �A�Sw~31��T�H�4�Yr/���}�G=$��|_l����)ܽD�|�{���_ۂg�]�����	��]D��v�P
.�l]I�c�S}<��@�>^N�۳�I����d� q�\,/�T��3�H�r�����y,�t<�Ғ=(�zCb"�'��YQB��wQ���v���5�2��u@�8�G��~���+sUray�d?��uw\0����1���W��v��c�s�@���NC�������|�Wɐ^�E������B�7zIgՃ ��>�y�/j0�+4�'�����k��,���C�<�! '��j���d�X{(�l�zh#q$�"| ��d>�m������N�f���@'��w���������J�4�{;�ĖF�:J�8+�Va&J��L�f|�)xҎ �U�S7�P�+�+�l����i�*���u��xHl�֔oy��LY�����b�Q�5��o&�t[��F�{U�����v�T��B�oɖ�m��@�Ϊ#�0�b���
���47ZN q?��
�jF��r`(��
�������%�}�j��T�0mb��>�_��>�|-ŋ�;����Z�sE������i���a#Ǵ��m���R�b:%��~}(���r%�{���$2��RI8�̨B
b�_ЯoJ5ܖlθ��e�I+z%��ju���X3���q�ZHZ<��a^V�D�/�%�*
p&�'�>�x��N!���<�����&v�:#��`�7��xx�Dyr���DQ�p2�-(������x�3>m�k�y��ڕZ�r2�"-�~b�����.�o(h�񎕣���>;��(�h�<�T@��!+�d#O��OУ�o�L��o`�Ss�&VW~̨� ��8
��ѵ�X��'��KK=�-]�k.���Iq����p��Oȿ���p�m���j�>�9�{ˠjj=��%�ו��4��̛�K�hkg���٦V�ڍW�Ys�-E����(
z���r-��.���*W��뚦fįxfCӐ6�N0#���a~�.��=���FN�H��K��]�q �g���f'2���I���Cb�3瑄��e���p�y��5��P��J��q>~�^���"ݛC�F���HP�B
�"�;�JO~�ŅPq�=����m����x���\�X d��q;��|���m����El�;�)�b՛O�3�>����M1�����CEXZ��B�N�'2�����q=X�ѧ��Ut���е_��HE،��C�����Z�O�ߒ��Q�}��u��z�)�i ��2[�$Ko*�s%�s�9qU��Rg���J�g9����7�S��X��K)���4g.��#���g�����.'��!5�ah�jZ�=�GpΕ���IY�)5)�����,�pn���ƂZe����p�hÅ�G�f +빮d�쏴�Jx$�,����n(^n�_��ke��5{tS�ܿ�8����J��>`����C��M�=`d�1}?p�A��n�3C	�<B��~a�'n���`�����)c��(�r�6�O���vC�8l� ��P��QC�>�UJIN-p�!~Z?���3N�H�_b�����T�H�B�]G��L�_�ރ�`�0������f��tqXp;�8WK�	'�glv�r}��o�K�5��X;�Oa8q�>�#
�����;6O�A�+ny�tʱ�)��oԥ�t�����������I���os������z�7�.4=�:��J�$`�Ca��x�[o �i9�"�i�j��`��-a��Ӳ9��b�aE\\�P-���5<"�@.�"���߰�0������,p���Յ֋_�n�	h�*��>��w�F�9��\����$����:�`5�,��>����6b��<�.ƨ��؊�<����"��l�ʩw����K�U���;ԭ#b,�,V��Lm��	��xu����(9���n���{��_|�OVX����)��SjGa(�$��1"�K����835;�x��x�8���������>��]����7��=�ߕ%����ֹ9"r�[������ �����bn� ����T��?�u��>x�a��sp� �/�$Jj���{8�5b`��ѭ[�5Ė�h�Ε�3)I����d��m e]��A��R��F�;ӧ;�cG�'�e�� �e�Ou�!�}�|zq|T���:!��n��㛿��PK-���h� _+߼�,�p��5�4�:�T)�O&�� ���c�迲J2Y`�+|�#�[� (�>e��5����~�]a�Z&�È���>�L�	�@�	i����ԉvLi����j�����2���l,΢��N�T�����DG������C�Y�2�ֆ2*?y�4M��=�V��L��j�e�?�	�}�9��m�"���;^���G�S�-@p�����g(E-e��u|���$�p����ٜ�ҽ[3䏁����� ue��f%���4��"�K83�u�mB֑��LD��m�Y+NS���d
���<��	M�k�D�J��e�Qwκ�䆗�"8������q8������" ���7'�
5r�=��(\ͨ�G��&fnE̺�?<AX!u��M����O�CM�E4�3�C8N�'z���_�!��ݨ�� ?"�m@I)�V�E��5��s_�o3�g�UE���/k.��;o�Q��F�N"��i��{�S���?��K��ٴ �&�J)+�.?dB�	�CX���!%����6�Q�&ʵ��ॷ�AZ�]�cp~~l���S\t!�j��%�L����ː�9$��*���i]!��ʣ������3P:��xR����x�F�q@M�)�j��K�Ӟl��xN?���#D�_�ˬnv$��A����� Nd�f�]����9�2R�L�����z�V��ۙ��aܨ�hQ���}BX-�����s+酺�R̘5b!fKT���B���f�"1fo�
��oUj���]{�<�2��A����rd�tM��I��1���
�9�W)�����~YD�'��	r�	���)}�,��Lu�d]c�j6��.}n!��W����F:�T�IPT� �~HsK�J�2�[���D�G��˖b	r �M�m	
+F�y)�G��⏋�P���v]�_4���k
�!���L�]�՟��%�v!��{]�1�VA�4bHL�Yfx3�e�O
��J�C�K�J���%|> �#u��0��h�,��C��+� +�M��%��0��St�իS�,
�}�����K(72��}�-�ּ�m�q������w!��[�'"f�Z�_T
�����:_�^�.��[�	�3��̓����D����&(�>�+ITU_ HX��
���Y��DX��+q�;��)����-8�����j��DƪP`��,���v�����'K�]m\��L?lu׶����g�T���?��À���I���Y�
C��3����j<��/��ܛ�}_��!��t$�eO�os�(�Z�rFu����&VA�4�O����:+�g.^Sйb{k�Y�W�8�F+�|܂:�~��+_TQ�I����m1����C�Q� ��h� r�'���cW�$O��eA�EfEn����]ܦ;�ܜ���]:�'j���>_��s�[H���LwTT�L�'�B)�L�ā
�7OGJ���>�{��pٺ7�]���C�Z�G��d+�#�rD��=��������'�"VSL>�IBQ�I��cW�[P�Q§�N�}/�Q�NL�1��+oRz�qĞ�r&�:�QT��]�v�4c:��0�����d��Q�vd�sc�����G����`X6�����BUpwmx��Mg�`P�&��yF���[iT�R��B��u��J��ߕ�
h�zM�R'����=0�i;n���{�;[Ni���^�n+hI=�mWN�$">z��[����p8i�`�zk׻�8�9�Zq��}"r��T�������6�F�X�_]MN��l��ç��}/���w��Z`݈��0!&���Y/Q�'N�������J�]kD���3��y�y���;�p"��2�)�ɷ�o�$F���	-�A�v�aC��=g��I��o�y�4���G��i��F�fUosC��^ZE�ߓl �+��(ԅuqa���b������qw�n ���JX�n^�s.)��h�&���,cX��g��v%w��\��e�N3ޗ�]��؝fS8�^Q-�!��;H���T�D]�$�5� �cRA�T:��{rCU@![��TQx��o�����6oE���g�$��:�ۇ��pHZZQ:]�m��1.�g�%��J�~.ﶹt�`�Bd�î�x|�h�ɣY��#�z����E�3Aղ��ز����&���)4�*���N
[��A����͵�D}��IQ�P0E$̉N�V�O�$�Yģ>�j����ٙ�H3L����z^2h��oB��H����G�ѡW1�:�X��H�S�n6*�o���J���@ϑ�b��}�e8ׁҔ?@��@BO!�0@�
�jLa�F������|�7L��kl�60��тﱄ٤��ﯖ�ڀ�?R4&-�UAQ����l�Iv���yZQ��kF�@�'�3�'`g�b=TQd����~�_�O�l��Yˮ�y�d�9��#^-�!�3]LZ`��-m8-�`��e\��0�pS�F��������1���SR�������謏�@$��;�R�ɿ�%���ۚ�h>Z���a���Y��G����ib�3�t�~d�Zv�3�~�"�v/�H�D�� ��M�����|��տ@�E����cK�� �f�:�Y��)���;,���K���9K���O$s+W�u$]�|Xu��KI� Y
((�%�6Ο��|D�[�b$O�
7W�;�5sB9њ*����d-�NMW�1)�EǄkL��qu�]E��c5�~S_6�X��Ţ�磣v���4�M/B�j��T�<OVQM�o&�V������F�)��Hv�)H�H/��*��HX�S��T�bdo?��8�'��T�+��9��Hd�I�G��{]L������l��0D2��ٵoW2�aϟp-����s��H�b���N�t,E�
���>��L�GW�����}�/�|�b���mnB��ez�E1؇�]j_��=���3��̣�4������5͟2q���?�F�:��.���Q�4��հl7�ֻ����Ǚ�^J񠲏�Sl�#�;�C�{�UTB���B�˞��4&�u������&=7���MK�Iǽ!�zE'c�b4N��+a�Ҏ�c��YW6�V���^�0HX%=7��/́G=Ҵ��	��n�3��Q]m��F����Vx�b^�����|�"Ķ�c��tm�Ӏ��>�]����Z�&$�V`��XG^EW��m�_���?
l���ʕb�Պ��f����r��Uvi�'8�Ro�gJxO<p�	&��.�ӫ���Q���L�}\� �>|w����[vֽ��G�Ι?��O3o�m�&�u2�� D2�&54H{nPG��7��ИGz$t�Y?�m�Z��K$e��Hu� @E���(��.�����,�{�*,h�G�.�Pa~�}v�C�G�[�I"�Ԯ��r�';3�IOm�#��L�b�!j�f%,LG�0�o2H�S�*,�N_ɢ)���~��o����"*������*;*X���ݩ��n�sg{=bY�% *�?sh�����x�)�7����y��h$��v��cr6��l_h"a��?�:����h���f��u�ǳ�8��jf5㕰�J8��a�b
Ͷ�/#Vzs��@HXr�l���R�Rv1
ӡ�J&y�q<��xxy]O1��4��u�����W"x=�Ӈ}K��4�������H��Zȡ��@� �|QA.���w�-�
"�z���V��Rh���b�;� ���]��a�	|;f?ۍ��*#_.�t��1U¢
ʪ�� qe���A�(/���~�D�V>
P�9xB���V���D`'�w�K��4�q�-ic��&�j���,�f�m��:�N�M%a��H1��4wz#�

��6�#�������V���,C��ǘ�1rE���#�w�C�%x��sg��f��̭���RP��.�ε��Uk�̺ƺvY��]q����n���a0\�w���ϵ�Κt��t���aUV�@�=6Q����8 ��B���*}k�ކ��3�}y�|	�п��]tgg��5I�`��q�6lǰb!3/֎R���KB�1W�/oɉ�#]���g��,v���E��W9;�_��Qi�!�Sb���E| hؼ#,���I[Q���7���{�TY��go�7I�(o����?Ia뺎H����������Q�N�=�
c�4����;H��c/1qn-���G
�#�|ʗňb�%Ť�i�Ar�\:A��8+��+�����2:��-v2*��������,q&5��fv�a05�W��=�1
r��bǌ3�����&��X�E��Eiea�@���w(ߩ��~�Zw�|G�!�v�!�t/��bXp�[G���P��z1�C{�$��H��h��"����X�t2�x��x���1���Fo��WhZ'��{/�?�;>���	�x�F�#�u���sX�i�i���f[U��B�Y�`.�y���9��&����~ڋ�6j$��q��2��.ȋt�n�k^	An�)�n$�9&@�x_�����b��~0��3��wu���Q0�[�t�&�;l�~�n	���g�ack��[Sp�Q���uog}��2��ɐ6tJ�) E~� �vͶ��jk$�RS�U�V�-&4�Z�4v�b�{�Ú��8�j�`�&�D�'��%�%��H^Q�x6ύ��/��*�T���9!�W�sn�9fk��*��?��u.�8�����>Y�Z�hB����K�j�+�A1U�`m���z���W
 �R�(�!�Ut���ܡ��R��Ƌ�#�w�!o��#��:�U(T���C���ڹ2L|l���d�$s��`�F;*Ǫ�%�u0�j�&�����P:/��[7�$�nk���C��@S�Gw������+�
���'Q���Ud��r>����f��m��-�{��I��D�
�A �y�W�]�"}�������&�A��+��E����f���O��V	9��>��)*>o��.��`H0FQ��ۭ^��3�XԼ͕ͮ� ���Jl�G
)��_���3�co�A����F��ȯS�}-u��Y��ן�cy?u��]s,�G�N<�]����w �6��\N�P
_�o$(������Ȓ`�	R��?��綿�Te�a˛�x�E�|����NP���l�����9]!ر��ܠ����y�ׁ%��� �Y�㜶�Ok]�_s��X8]"���o�5 �T�2�JX���ց��^"��X�D/%I��K��Z�6y��Tn/aZ0�#��n����6_�]B���Ŷ�T=�$ ������Ū�	�b�ܢ;(T��_�h� ،�5��ͻ������p�N�Ei��s��WU&oaf�ߔ�}-(��~f�R~W%�pZE��B���{�pҝ��g���D�l���������=�@�E�T�K;��sI�[�hC��X�ASv�:2�ʀ�:�6�8�J�&��o������3T�V�{���X�;w���������iM��h��=P�#�0u� �@g��Kώyӓ�&������h�x|�-Ei�M��t��v���ZUO?�Y�(m#.�I�ji-�r�u�{�s�L	r��&�fB:�5U{�U�A�}[���<�P~O���,Ğ1�jh�f!e3��-�#.����ҍf��`f�h~�����X���|R>�.����f.�˴�T@�$z�QRi_�n�oE4��ڋ�u{:���S<���K�bA��,�����h�i0f�d����I���$�2��'u^e�%b�϶@�L��~Cu�E���\`��/��b��*-�?��ʧ������21�\TڵDN��c#5��+�5�"7�~��h��G҆b�|lg�Z=hiK�ɀ�
���/�R:m�̭B��zZ%[ ��a%҄Ӧ�M Y��Xή�t>Ft��6�0բ����K�i>�S~�9 
���/.����\7�~�����:=�t�2Nշ��
�iQG�]�@�����ېm��3�����ph4�)UF�<�/�L��Q
���xpR[�n?8��K��{��)_��^cU9H�\~X2�_�9ǆ�X\�/��b����O�P��Qe�,o�.�:8��)�F�"ET:��+!���&gM[͡����ψ�+��cI�c�?��&Ц|ғHޚY��:~P;����`��$�����)]�����t~%�&|�d$F3.I̛|RuWP��P�'I�8����7~x��&��-�*��_EqwQ�G4��W��A��#2�~�A��}�'��RI��B�V�x���Qj
@u��8_$���,h&|n��w�L������I��-X���з��g���}U�o�R�W���+��#�{��tR)���V��$f扳l�U��6��b�]7�b�IR���g��e��=Q�^J�r���5 �[A!�]<q�Q��Ӎ٥�6 UX�����B�"�I��\�%��b�ˎ5��ͭ��~�(�՝K�/�����Ϥ{o�^N֏�|[LzS����i�r�y�\��DP� P���^v��~!g�Hl�J+��'�\��(z��~ Z��߁�{Gy}��j��^����\sU��-f Gs�װ��?�����nN���R�҃��P�ߪ_Z��Cߩ�8v�#��;&�o��DtS�T�ѱ��)(͔�d��ш1 ��k�P�2��d[������\���$4M����l� �u�5�w�4�*QО;O��'h^�V��0����ua��Pv�����E'��+����D�s惍W`�3tK��ʨ\�l����)���C
M����B�k@�)H�JN�Dld�Q�6�"n<�-i]eGJ{�֯�������W��}d�@Pl�+n!3J���̉�	���;�&�����s҈St='(�{���H�-����~-J���\?s��M��fX��s���^/�8x��Ժ��*-�U��"���^z��<�PA\w]}J�r���o%I�V���X��;G�nC�O`a�m֜5#5�r���`���ʣ��=N���S4�Avz�sF(��'���>�e�{�z���I�u l3��!fwp!�fե��Me;5[�㯕����d(�!����HFn�r�ј=��X�+�zm��Ea�d�hgg2i6�jy�-�=;��BXG��]�s?1@#����d9�gB��
�R�A���`�5��
��b�/���83��U�HR}wF`��x/Fpv�������.��ϫ�G���<��+��r�a�Lk^��]�`��i�l������)�-�b�XS�
����C�G>pӠ�K%yj`�$�s�L�I�l�j:�R����:��>]v����'��!���>"J��W������oФF۔�c�끱�a^h_U�d�)k�[3B�}��[5^��2�m���h���v2�s)���Y��ɩ!��^�w��l���b�k�:X���n�Φ�4i�Џ��v�X$Qar�W�˄�ϲ��C(ڈ�5�I�5Cu�t+�Qb��.�Z�H��l)E��;ys�fİ����>K�k������N^�Fqi�Z�Γ��z��r{Z�5���Bن�J��!\��"�y���އY�M�l����E�"n0��VlǪߑ�A4�3t�5)�o���(���*�$5�[���4����mg�{'-,̦�$$B�a6DF�(�6.*�Qnnk���a����3rH�S��J>��l����nw6��Hbq�7��~#��S(����P�pxȼ|���!�ʲ��L�V�@�f�� �h���{(*Z�v�t��&��s�*����;j�ݤ+i�d� ǁw�8��)��%�d9��ؓ��)p6����N��b��,|e��<�Km��v	o��(��:�o�|VJ���y+�oMM?L���Fdw�%H�8!���sg���g��� �wEn.AW���E�)�i�@�����K��W��ޕ�.Q���H�xq�A��"
�SA��c)�d�f���[��W��29��K�p'Bʌ�U���\H�'�Ql_�*����ݽ9̅v�1�ME^����p����s���J��.!�Uʦ�iB���'LQ|����e�]sK	�ǰ���N��}Y8���d\�ԦMxN��i*�_=���z"�����=+
��g��u��΁jI#c>4���@���*o�G������#�K�5X���︟�,d�[R�?�1��Ɛ������Ō>��ȌS5�=�W�T�~d#���R�����3DF��p�k��Y9 'ci��7��>��y�9�ݯ/���Ħ�����yk7�F[����/݊�P��~@��8��"5����^p��'���2�8E�.�ݾ�W�IxZ��Vd�7�м }��Ǵ���i�t,k���8�[�ԃ��qD�����t(B�̧NaZ�&�c�e���5�L;;���6@�%&��@���?���r�a:be����l3n���3]1���Y�G'�.7��Id���J����-6 <�i�g���;nD��jD���3U�zd���;�5Hr^ְ�"�ىg6_�p��)�x�
�?Y�6���SkCn����1������+@Iz��_J�t�j;b�&B� <L���1��^��-1su�S�������;�z�L8�����|�����p�-T��!A=�X��ݵ����Z5J�.�(�V-7�����H����̲�������TD�n�K�+nk�R��G�׿��f�;!ճ&�x��7��!%}gAy����)g��A���P5��� Vu���%�O���u(�i�� �X�����Y(�%b�^v�2��V��_�M݀����4�~n�-;���>�w��Jp��4e�����I꣘��V�5'�Y�x7����y��x`�X9������޾q��h��O�5��$��R{�;�34M�';�h�V���X���`�F�5A�<T<��.��^�X
pd�
8��=|baIiC(�2u�2����œn}?�ta�9���f�χ�%c�Eu��1m�^�οvn���{Jh|$��-�/p��0[�M����/��{���t�@L�S�K������:��[T!���Rj�*�^2��L��>U��zV?�裡ǋ^�ֱO5�_��߁|&E�$&�{��2g�އ��؊�c�4p{��&�&OAŏ�����X�ۺ����]͉�䣷(�p�SK��v�B�7���2���T6t��ݝ�ĵ��������&ͬ�����M~��/�M�|y9�8I�q�w�L*CM![<�q���G�g�����N�0�����ͷӗ>!v��
��73+���Т�}G
Q����{������A^I��%j �燸[����A����g a"�'���UG�vݞg?�oҜ���$9L_�S��<�W}�9"gQ���6OZz�0������g�싮��&����(�4C�C,�#�Xe��$�׿��~�.-T�嵐�g�sg���I�n�x�S�o ��v=�?'K7Ճͺ�<N>�!�H�w3��9�P��Aբ��f?_�҇l7��{ջ-����ê�
����FcQK[�Sko��iP�E| ��?t�Oy�,V��E�$T��#8��U�v�f�@��gR����M�@>_���b�ܥ�Bz[�2?����ph\���u���	H9�Ű�:�s�?�X?����7��1C)鴥1�fQK7!A$ �XMd�pۓ5s�0:w�A�i1�~ᩒ\�-`�U��!�zhL`��Tw~D��9���PT����o6������h,��)M- =q�L쏏AR�B�S���q)E���I� W���.MC~f�3�
7�@;�� ����̋ȹ�j@�6�
G�����Y��8�j��ef�'$��3+��r8p#Ź�m,�Ɍ���2�G7���� �Z~��6����N�|ĮR:r��dP�@?؉e�E��tR3j�!(3�!ߎ�Q��:��_b�V���fi��+��}��u�ĹL�CA;�|.��nL����F �b��˰ܰ؅,�$ۆ�=�cDV/������_/�;M��zN�x�*��[*�*��7zwS+��r��È&�T���5>:����N��Z>ߍ%�s �T=����]��1��X�khP��"�)�Ni�1JC�3���C�����_�xi�^շ�HD�A9���F��Q&=6��� �l���#0��*U���hC���8nɴb^lw]pD�g�x�� �"���{\�]L.�.����@�ٶ�5:� fĳWP�l��v;0�*Ş7�~dQ�_�_���[bn.�`(.�o�?><�sF3J���i�0�at@d*a��3�9oքـq���>�ig��XS�DK`�u������<�9<Xo�t�"���4ʸ�j2Ym��M&K�<�������z��4�&Y�_�o�Q��YK�R/*�J��&v]���vz�c���ɋ_���N;Q�eᳱ��)�ܰ��4gK��:f_.۬J:B�9 GL�\�ވİ��X�Pz�z{�B�7����q��/��4Rd|��{Ҹ���}B��0P���j���w�\"/e��̆��7R%n������Y.��^��u��u�3�n��?�[�&}��^�C���&���I��ex�)n ���j�}	(#}��4t�����de���I���bTo�RI���ƱW��2#~��Bd�� �֧��8zf1<�z(�Yu��I�/�R��-+{��6;�Xr "A��j3��@w@]m78Y �%��0=�������׍�]���+�bŭo���b:��]#���8>�?�d��������Y{�>��n^Se�V�[�wǡ���� 2T�L>:4+�ܥ��^��)�F�:�5�3̡�M� �HE�H���D��m���]#���O���7BM6oW��������Kt3!�ZS�1=�B�	��r4��z4���$7CC�'mY�<���M�f����A�*�:�����Sb�њ����J�h</�4�p�>�P�7�a��ˌ&98���)p�*�hσ1 �H�;�|1�2e�M�2��}�3'�P������|֞ߕ�a���2)�!79��F7����뺣P�|.��h�Q~�8� V�,n
�^F�HwT�<t!Dz1CY��%��)}��5��X	M	;�&��rj�	�JJ#�ˌ'tU�I�g�FѳlDA�*�k�g5����F�H����'��r+:����r�t�am�+5l�9�\��z[��s�٬,��e/�OS6���dJ��r�Ζ�>{_�V��	\���@=�l���Xf���[_ek�C��p��by^~T��R�ߊ�c��0�zE�&�6�}�+E���ϟ��!�	7��V��C���K���:�_����q�L�Z�Tm���0��](y�Nd��P�����f$�xģ?���������iv���]�3��<��������U��n/��,���C��F��2���*^�+ ,sEQ�I� ��}!/��ѵy��G�˗�L��*/q[�_6�> �q	��*����s�A�O���T������/������T���8�&;� x�ŋ�X=�{aW�E��*�����[��輬dN�^HE;���69���Zv*e���u��7�@���p8Y|Qi�A3V��c��?��D[*&IW!�W��@�&�3��f�K!mp?k�o�Lm�φ-&�)B5���-��'�:�RHo�/L�)�L�Ŭ��V�m��7E�*��4hl�T�����:5k�=תv�5��t�#������у���-!D���%Π�Y���5%����|OP��3 v��X*���e��C\�^[�M/DW'���O������K3���&�� l�/���J��!�n�`��MVLI3��q&�a��	��Z_���{P�9�{-���b\����eI�t�@6�,Gn/��~4���U�Q�C	�vY�2e#�}Ǥ�Bڃ���K���֔�/�zim���V�Jw��&����n!���WfB`��y�SH��eQmfHȪ_�Yx=�=<����*6t/�h^�z�QT(���G���S�/�KG}�\'���\��~q��dv.�JͰK�K%z�M�c�Q���;a\�����҅f�+N��ژ�&�<���x������^�V'���I}�7���Jj�S"N�%.��]���-^0�F��N�.��B���
�-Y���I�|D�Fx��V450$ܐ��5:��	�q�Q)g�*M�娷����J�g�"��T���(�LI��L� F#H]ھu��=��9�@��b�NN��\�����=_���^s �1�*�E@ڞ$��$	�n#�VLMvV�SVb�4�O#���W9
�&Q����G����OT)����$\����b[�+���O�W��U}])e�w�뻓{i0t֩���1�2���){gv9S {*������~l �\���G�aU�����/Ȋb�*(���>�p����E���uw}��Ț���f�s@�(*cx�z��S��f�Օ�"_/}jTj�E�U����
�2�ɯO%����q�#�[3��	�H�H=���c� A�z5m��y�̊�dm�c��	7�R�?2f��".�T�� �v�L>���PIX���
��X���^���*-�´<��$��zA�):JwW`��F +�6��n�{��:�s��7�$$v[��Mwݗ(�F2|2�up+<;��J����^KSG��3E3�;�;	��i��a�ō�U�j�������4m;��߾��Tݫ��	��j}J�N>�l�T��m��E��Y�!4!UR��?d�C�ʨG�0с��Q�>g�xp}�A��yI����C��h��%s�D��3l�pї%��Yh'��}�?��-!��v�Kظ�=3�W�!�[������XJ��!쓨`�ʱ�Y2����`��q�*�۠�� x7V�2N��X?I�fbfϥu��������mW��糟���}�Q�_�{��{�Ҥ�h$��"LQ�,i�;��&Qs���1�d&AI7���:���/��"X���	4������w��������`���#�u�oL7�����O� �?'GΫu�e�9�q���
]*-7B�t˜��h ifCЧ[���̫��O:�~��X�{��FY�O�����
B?m-�B��
�۫3�������C�]>z[��tZ��X��Zݡ�u>u$HM�$�p�G�Հ.�/����i������3�"i���,3KCp�S���K�><K��A�CjK�� ����8��[��n�k.Y�dVg�P��k/�U!��2�ƭ���:���`vE]�Sօ�����f/]��71��HfUi,�b\��Nb�L��*�*�UD�i���4��������c���E�2��(�!�Xp_���X�=�+�~c�W��3L��"6=���s�����s��O0�
P�ʠn�"l�޲��1:.�C����n������%e��À�#ɹ��|�=MW��U���zѭB_	
�;�	J����_P���{�L�����Yqcq�F����ٗ]?�V[Ĭ��Z�}�$��5,|j�w�j؈���Hpg�Ԡn����p^��'t�e5RЉָ�� �:��E(�:I�a�^$�����q>)>0�)t�������ڈ_��+�fdD�p��E8��O՛��mf	xy�M��Y�R{��m�����$���LF�3||�̠/b�U�]�Q"az�j�I�c��<_�b�`*�I�v t� �X
�!�3^@�9��	j�)6M|T۬�h}oJ�)uzm�-X�Q��c�+e3G<Dg�E�㳏���l��l�BZCfB�ӓ��V\0���!�OF�S�v
_�!�Lλq��ǘ���V�E���&zM0W}�xMZ�^eU{�%���"�1�nf�rZ�)/��dM��ђJ5��
��Qh���0�|s��v@�
�JqA��4�h�E�o��=d�.�Ū�?\t��T�
��%3Ţ��0T4�a(oj���y��y�����%EYy�.�u�L����m���IAh��Α"�=uj&��F�[N�ל�c)��ơFͬ)x�QU�~2ȏ����]�D�D��%�����1R�S����|�D<7���QF?-�2��ٵ�N=̃���tk�@�|���9�D]�n�ϲa���\��	�ڊ"ir�.�צ��{�x��0A{��b�K��_�d_Rh�*z��=i��Αl��W�|�A���VČS%`�j�)�z�`�Qe�3�qk�[=Ƙ�ǈ �{�%�&��Sy���6�{!h��i]��BVkXy�z���O_��"gQ�A���j-c���<&��9»�Ü��'H�%;�B�ɏ��7�������W�bnQC����#�4��!D0x��Ӻ
F�Qp�U\E�1�3�P�Õ�m4A���b�kE(��Y	[�)r���7�ہ����J�Oi� Crr��v�/�l����\_�L��=��܇s�ߎ\�;�b�n	U�x�au�h����w�6`Hz%~h���b>���XnN�;�+rv�u��g���d�%1/�j>�O�ud���c'���#̄T[�%cE�6_�7�����+�� �FF�������sE���԰�[Z��q�w�����A9���Ad�@o�ႀ��m�f�1��a�Z+�����ٮ�2�j�}%��+-
6T��C�n����GŚ���zD�w�o���F�˷�Ŵ��_��"���s�~�6�xj ���w�����{�H6���wa:��҈�s�J:�s�E+��W�=j�|�z+a���H��8��Ce�������g�:	�q�BP,�N|i��Փ(|�.�.�+�ʭ:���ψ�ز!,��U�#���e���N�I���{�N���R���V����5���Pb���+�"���Ԯ;'9x�Ʊ��B�%{]���=鬳��	�fsL7�L�3��qh`��kê�=v ֶ�䷽�*1�őR,��>."���=��n�W�@��+��}Ŋ{��OY�R;�6�K}M��
9���Q�&b �� ѕ%��	���z`�;t�@�d���bJkQ)�U0SжM�{2���!�Qej�q��?>��^�%w�aO�i�<��7i$9�K��U��x����t721�X􇩩J8�h~5�Q��J�D4��Apj�C��1!���B>� �W�"їq`�iʒ0~�.���6l����#$�6�D�ә�5Q�CQ@�ڙ�ʛ��]��A`��>$鞖��Ҕ)T�8�݅����d2���6��[�0#�A�:���t(�[wfc!��S����v�����"�6"��U X^s�u�óR���3JSg�EMO�m^�AX����v)�<�H`��/��Kl�V枎�j��0�����C蕾� أ�w  b���:ۈ�#�R9�w���d�lX��g����bl+ �G��`�l
�.^j!"��N��{bK;��T:�Imej��9��O`[`�Oo�Z��^oJ��&:g���*xF��LE�����ͅ!�����ڂ��6��7L�d�}�Z/�[����=󯤰�fV&=��6V���������b���ZgIɈ&�&�+TA)�g�J�:�s��f��#�vjvi�bk\ � -N�LW�=|L} ����ZV��?a�ћ�]l�&Q>�1#�۱j!9��e���
X���"XerI�X�Hu"�O��J���&�OYn|��(�L�4�{��_��F�A�:���h��oC 祾
�}Dͷn�:�S?ZN�%��RĂE����� ��ӯm>�'����n��	�=�nnz)�Z"��d�#Ee�ֶ|s)�S�`j���+�I�~Olsb=X#��A��`E����4s�z�r���M,}�������WYР���μ�*��U-�@dƟ<)�%�^������J�m�d���?RsTr����P�8V��#,�g��s&i�,��۾�����z�m����2/�x{=y��R�8�N�@OvMQ|3ܵ�f�#��8�5Ӭ������uH��7��DT��B��+nL]�PU��6��&����Ю��p*L�2u����!��/��Zse%i�x����P �T�V�q�*��0���2��:#�m�6Ol��A&�b�
�@^e6�wfB�'G���PF� ���Cu�n?��xd��㻞
c��,ֱ��h��؏E2?U�Ot&#�:[��ƞ;(kӈI�f�_�� Et��S�Hl9/�,}��ȚN��A�/g�)���W� L}��r��,��:XSIǸ�guZޜ�GG:������^�3�CɄV0���f=�A����EG��1�,jl(oA�p��˧
��;L��5->��<^�w,AO���Z�d �#7(إ�X�Pc��O�e��=T�x����C��i 7�FX��`���ek�rlI��k$%)��3��T-9�W+;q�70��:7$^����xN)N�N�Ҫ�"T���>�m����"˿�B������ٷ!̽Az���K�"�_�e]M^A{¨�Z
����9�>Vݏ36b�xxN�����}� �s|�GJ�e|(	��C�8Rm�@�jؐ���-�_N�:N�����q��9�OE5𼢰(w���,��G�Y��o(cP��7\�\qC���J	IE���q�FMbq8?��%կO�}�dF
�Ǥ�r!��� �*ٜ����.�Rv�d�ޖ�ߕ��p��-m}/P��A��D�:R��!�:<���Z'r��ZE���z~���$�LPsN�	��3����<u0X+���%��kVi���,+=��}:i9�mpθ�1�*�&�\������TH��՘�\KM�g��2$�,5�1 �x�x	X�N�|���f3;�j�a�\D�FiN ������b�(6N\07��'�!��޾x��[Pem)�	�R�+`Cp�+߾�`:�+�
?3�=�b�,�1!p����Q���:�1�\@�J8�вǧ	�,��}F�O�v���u4z%��º��F��W�EYx̧?ź^�\�rwn�(|)�3V%.�X�IH��ʯ�tv��(-Za7��mo�;Fq;�a?��M`>c�l�!7��&��ŒY�V:㸇����h����}u�6��C����׻�(/A�l���}ӓ+��pY��~� 0�QY;�ۊ�fU)���kr������	ϪBEe5���H���s|��-�:\��=�3�$x ��E�4�cȶ�VU@��R�|�����-��6;H�F�UI��?�=E�S�id6����P����xX�u����T,��wI�q�|=�H��m8�pŕK�z$Em�z���VFf���P\�aa�xr�[;�ԂJH jr8����Z.��vzAY`m���E�.L�-[�C��t���b?�yb޵�W�V�A��w�|}�}K��,�UJ׸�9�-B�xI����r������� +2�v��]z�+�.�kE9�T�%���u��4��������M<z��GF}(��9�+�c��v�����$鴓�)D^�V��W�̅=���s�֦CW��Čz���u3Sa����g���-�}��"L��Jq��k\?W}w:&y����6�V��f��S�f���J��C��{ϸ����(z3�y�ү��a�����:��=�H���#9�kS�Z��4~j		]�Ð>��QAӬU�Ț��V}[Q�[S@�R㜟R��(�*��;��>-�Q�^eRK����:�Fk���@��\��Tcef$�A|¯�c��'�+	�^g���8���1o�G[E�&��e�[�;���Y�k�S�����@�����>Hg�	�p@����g��p٤r�����Dе���`���'�����թ���>��>���H}:�I�3���%��=bd�r�*tũ��YSH���2Gx�� |���lBT�
6���0�c�R�������L���Kjm����G�{��Zۖ��J�h�����RZj��	D#��!!�H����<�5���x͉��J�K�$�Ő-����_�V��|��X��A��}�_�m��C9wA!��w�j�E�|1ŗ_E��2˚������{���ڷu��������z`��~�8�<��y^�#�l�i��:�-!�5^�[d�.��bbn�9JrM��+̴=?<�$1��sN�5vG��7H�k�j�sa��Nf7�#���Ŷ���U���G��� �*�1ϫ�O:���3�����SIPM��2u;ᲃ�/���Gc]=F����o�ewn��0�>vC�l'վ ,ߊ}�:GY�fA�c�T)A>��"�WEv:�~��E�
�z
B
�=� ��6M�������j�5!��NY8چ��X��{9/!�xH��q�T0��|4B�ɛIns�1'w��4¯���$��z�D��"�R=8�����TQ��:�z�*�ROʍ��'�6a��V���oت)�:UV$���%D��3�.���)^�_�UiK�
�!y*��#x�?��Jp��(��p�|AA<xm��)��D倈!���r�S�l��9pn,'��4�K�����}�� &���`,lW��7�0�n�]r�m	!Ϧ�˖��s/�aI��~��|�{���A����̭My1�T�m�{Q��%�-:H�l��&R��10��=������`�"��oG�A��J`@��8�1�[dA��eh�I�/:�]��\p ��v��X8��t���c�Y݇�>gIK�^S���u�i)��ME ��Fs���Prl*����m��b����%_U�7k>������"�x8
e��Հ��ˋ�j��d�-�Gɰ-���� ���UZ^0��y���69��Sy&������݋I���`�=d$.�:��5N����|�A��Gc����]�j{ªq:����)$�㫠S��k�S���э��O>�+8��"M�<��gJ���ng
�ӌ��Y���"G�����CV��{NF�ˏ�;�!�pXP&�������²��� ��n�5���j��N�r�U g�ܮ\\��7�W,��續ЮRH�&}���6 �Ltw�H8E��B�~��$_?�+G���b�n F��U���,?��>�7�ߝ���~�&��ް�!�z��mK�2S�a�b(�}�i#`�R��
6[��}]�� �6	s_��ƴ�����$
�&ى��@�VD�u�qщ�IX�1lY~Ґ���6�UU��p��" ��=5 /́f5R�f��9��s��n�Y[�|fˮs�i����$9�nc�m�P��=��t�O}�dcr/�`��8ɕͫ_֬R�I�C��r>��6�pLv6r���y��W��"3�͕cSj�:\�E�45��cɋ�A �p�Z-�<��+�$~��<�XB|Wf�k�DP��v��C��G�>"6�����u`���ݿ{WP�]�o+�)����dw]}8�b��z{�/��6�j����2U�GҲ�%�`g�bwƢ�j�H:z�왆z���~��V�kڋ�gɊcSThުHa �v�I�-+E����U9wt��|�������Ǔ��~ӗ��#��A��kc���c���S*�Q�]>ϦC4�.���¹�^��T�N<A�ǝ2c',L�S�p����ըkpX��^�x�,&�LPk͋��u�d��А�I�ݐ>�Y�v�.�݅hn�*/ܱsCL�F�S�n���+���� ���V�51�	���s�H2_b1^�N ��_�Uۣ���}��1�4��R���)������S��ߓ����i��������jU��I���e|,��L�R���~�%QTY��t���D���|�8k�о$�KnNb��yM�е�oJ�Jv̙� �`|?dFBJN?(X���&�CGCz���]O0%@)R�����?������{�����0�Gw7��Nj�im7�{�2� n�yzn���4h�Z�ˉ&*�A?�Ћ:9���a#,-hm���)#i��,X(,e�~�ʸ6�����V�b�
'�k�x�m�,��l�/�;�}���RG�FCܜ�>7��v�D�p�^o�j����a�R��o��Za'��|ɗS�^¤�6�
�߳_�A�WF���4ec����\�6�qo%���'×Δc���϶u; ��R��<)=Bo�]Ƅ�{��*�(��l�R^CvWwoyz�G}F󈋿��f���C��0�4��3���F+��3��J�Xo���p�q���;��W���_Eo�Bu\$;�c�.��B�����,��x�hk�I�������o Q�|�^03_�*P��Q+�k�Ɩ����zi+	�����N6�Q�3Qs��и)�͙;J튨�Un$k������*���OW�2B�9<-oE� ��wV�*��R�ą�i���\LZV���Z!�� �T��S/3ӯ��j^K��,���`��ѽz���-���B�G�,�*�箎?r\�G�����\�Cݞ��N;W&����������[7&�f���üQY���"Q�a���t�'6m%���_�Q�Q��F����o�h�օ��iJ= ��w��v�v�4���o�u>��S(���b��#�ܫͫ��y�1Y]@�4Ӈ��Xr�Y��f#�J 6�q�H�湟,�����R���O�(�Hl=�>Y]dq�i��jE͑���WK�s��^���]7���%G rD���l"DX"��Y��t.���0x��l/|6��g���o�l�r�T��h��!��Q��С��$9i�:H���Q���T�{Y�5��dTS���z�l�% �ܥ6[ ��E����q�l�v����NL�-i�B�����J���[N�XX����'�<%������V8#����P�+;�\��}K���:5�=�bT�r�&��چb��m�Lz;��:�&7��e��5{q�¬�8�(��`��@K����`�V+����ʇ5�>��-��gQTx�.��GTmm���ԂH�TЌ�%p���Q��I��E���y���w E��Uh/��N���^��'�}�6�{%��[P:��ۂ�A���C0#*S�	�cy&����fL���%Ǌ�x�rsK�[
��q��0�`�`����C_c���q���,zJ��g��p;zS�S�/u
�q��QG��'�P㡹{�iB�бfh���&�otW;�P.b��X7(m�w�K3�G*SL��u��$Q ;4c:g8��7����Ӭ}W���
��-��V�u/h����;���a����Hy���N�����A%�؊�}^���EJ�h�K��f {6��Ω�"�/!	�����X{��ހ2uu(f����vYi-b���c�\)���Q ({��\���N[�>l��r{�#d���F	�����(� �1�.?@ư�<� �	)�i�/���d�w��L6Zng�.-��{!K����ly�>���`�����%���#��He�W� 1ݑ�\��@� /�kţtLvPI�.k���F�h}�6�1��Bͪ�.�~���`F3g��̋�/}��?���f�z���A�	ܣ%�ś���v\Ah�註~fy�M1Y�Ys��w�}�Զ�DW��!	*�3-w�_�VZ2i�Ƴ�� ǟ��7��~�C���X�-[��"����Y^W7�T�(�zV�ǘ���#�y��JR{O�p,��O��-L��ɨlmfM�H0㘆b@��ft�(+���u��)�Q�Nt�ћ�+�N;K_��].����w�0Mm-+A�kiP����*���K�j�C�]
&r�����E���bT��:{lq�����s��U;{Cq���W��y���3������Iq���q��g��*R�h�ٸͰ��#��e4+>�}���SNh1Ӹ���
���ډ-����K����+%��1)ѡj�Va�LX�� ��х��է��9'�RTh!�Ӕ\E��־O
�)�.�j��]y?<I��-Kp0�YI�j��~�FN�f%L��4}_5ѝ�:�@K!-0� �\~h�dR��e�UW��5�q��rs���8g�j���`�J�k�p���|�{R��f�#�'O�r�.s�����<}2��=��Oxv�]�tw	^�����`��D�zf=��vzxj,m���m�Jř �t����$C�Rkr&����|�Q?���n����z����]�W@��Ml�'�4!�pZ�ؔ�����*��_^@%%v����B���f$D�Á����(2��!������A�82����Sr%�'EID"h��;�I�jfIe@�n����:�j �H�r���7����|�il�8�|��󮼼��%c��<Ȅ�-��z)3��p5���2�q�`�M��dZ�',��au�A�d$J�s���%SVK�D{��g)���B��rM�8a�O�1���6�Q��a\%��W��(�1i��ӱRH������[y/�(KY2��8���Q]��B����"ɍL+� ���-h�x���Uk�+�ƣD���zn�`�ʓ��F��tX��W#��GʢD������_��I��ߤ� �)���c�dY�.������^���u��F?�~�޳s57B���FPz�q$ni%!BW�p�1DcP�eF8J>(z_D��Ev�r�)2���$��%ǡQ^wUit�FjHsAQsO���C��$'ұ�c�9����.P��7����W|	�a�ia~2���!1�!;��ԧ���N��nС$EP}��`%�<��L�Z�[}U�c)�M�ED���iQa`��K�<"0s\�R�\z��5�ȱ N���%\P�o���"p����1\G|ie���0"��G���������l�hcx�,���Y�z1d?�@�ױ��_�3��)&��y�(Эt`�#�ʩ�����ᶗ�5����	ߥNF��'zX	lWy��\�o��)-�	y�W�"K'����� �`�*�� 
�sT[7��e�L�K��U��Z�s�������9���Ճ�砈g�+Ut�%{!��U�-z�ht�B����j���Qmؐ	���5}��({��Ӯ6�<R�R�o�x�6�<���c�d�F����Rq�д5�*�dT�xO���A�0���ñ��]�E�0a�}��a\qʶ~/	k6KI�����/e��vݺ����9� 3U���2`�,g�s`�D˨�X�&��l�?[�}�;�������]�<��Pn���	!.>k��C#z$4:�W�{��Π��K�ĽhO��|p	�'�-\��J�%�-�<oW��
�k�E��zޝf���eN�dl*;$K5=����Y�<���A���Aw� �q�����qS�G��r�h���`�{F����H�[W�Y�U�;��2��j� wbj3�Y�C�+ζ5%�?�k��	"�|�&b5]�+jS9�oo����gG�vXɸ��� \��}��O�h�-te��V��v��R��B%���	�x
���
�!DƧ��h&1�3S��Q{�f��������X?�,�ާ��5��E�.t�7ܒ^hNJψp��j�Y&�h��4W]B���u����$l�bg�}Ω`�E#�0J��\�$���&����+�ڱ��W%��wi&m�h�ʻO�}���/>�[?0F��_CFl��<,W�@�n�V0e�H�0*]Wy�3��X$+_k�@9��ȯ���՗L�<�d�y�:u�KU�f���8�'CP�e}�[t���r�6��jŴ�G�bo5n�:�+�U�E�i�>������q��R�L��� �	�x�X��Y��L{�PNy��!J��"p8��`]%���u|P��CoZWC3xJ�tq�8�y�;�x�'�b?�N���Kк������C���8�N1#�BA#%�����#=A���i��~�@���hwŸ�-��q^T�s<-i���P �xVc�Q!*n��/�)��9U�a��$1�`����ć��T �XC,�%���o�pX�~�ƙ�G��IG�o�L�`K�R.�Y�)�'�Ӵ���v4U��a]C���o#�^����m�'=��6.V�$���nņ����/b�3����,�>~v��1���^xďf��}�������z�k
K����
s��	5Тw��4�mmȔ�{��I�G~jl�RjF#,Ē-u��9]jc�F���l}>bq��ł��.\��� �f*���R
�(�AI�^!B�t"X��|i+l[z��d ���w���l"���j(���#?Pw%B�n�8h���cj��#-�1Hh���M>���"��(	��Oޫ�u��Q����M�>�c�R����p��n�����]��$	~[��.����'~Z�p�D�q�)d���#�o(m�]?��	��U����;�@�:9r������Р�іf�έfj	)N��G��Z�Z^3�_�j�D��H'�`���ާ�g��rѸg���`zjb�q!Y�/+pkbk� '��!KP7 :�&Jۥ��Y҆$��&X�52��F��IZ���d���v�]�
f�֔�Q�QXW��9�;,"y���΁��B�� ���b����Ӽ��,8�rWh4�&�������J:8������r���暔`Hi>�gT�(#�K-@MbI���O������T�E��X\~��t�F1O�M^�3
�L��x��(	B��+#���W9�Һ��k�B��N�r�=��OTF<QG������`�,"��ס���E�O���� 	�٣�WO������:b�)�<�3�\��p-5����]�;EG��7�돃jB Yα�ߣ�h9(���<��G����pj5�ȶ�����
j#ť)�jޘ�QE�)ģZ��pz����7�.���Ц_�3.�Cʂ�G�`q���4#$x��~ ��0��[���tMF�ߕ�#`gyv[�$|h�p�3#�$����JX/"�x�x�����tS������C��8�����c�G������]r8&��;'��{୤&E��l��ί�=�F���`	�$أ���k-݉���_�B#���4�>�5��W�O�.<U�_�,oȬv���rY��?m�\p�� �U��ե�!)�;��O��m;ց�����Z�5� �l�!q�*?.^���D�}�+k��|�^6�5��-=@ak��G8��!�ښ��Vz���f!�Wy����-�$!����Uvw�#�Ґ�FG���V�eݩ�� �Ҁ�t���ۄ� fY��et���#k�	�t:�q�	 F�S���{����k8��}��������:��p�
�f�E%��	`Q\�Q_b/��24�O���kI�?�Ʀ�+��A>��9�of/�s�%<����r*v��7�0��[��Xu���ʏ�c�<,gPY�o{��+�y^_@T}�Yt���z�2� A��X�_������3zd��v_Eoo��5�Jy���QT����NZ����a&�~�͍%��z��O�m$UImI�!����n��o��d4����a�M�vw��� �K�v��e�O�a��7W0��z�?	�f��[�u��T6��wڋ�Ư�(�R������"���d'��]��}���{듗8&����7Tq�5��C`�&2�UX�6�����+�
9��cqZv+>\^ɂ�ND�>��ǅ��h/�'�Lon1ʞ�\)�9RB( ��`��h��_�6]�����v���"֮��Xڪ�p�Y��&�L�C��G��ND=z�ou����-5e����3W�o}��N?���0�y�&D/Ȳ� ~�o��l�}�0',��2�Wg�"I\���m������G@Rl��P�^�ɝWf��^�i�W� k?��\��A�	c	�y`>y�Y��6V��?CV�ג���Gwz�i��
��ӯJWhI�<��:,P��2�{J˅,��ѣu��T2x����Q��b���F��X���2Ƒ��)�Y�t��2�{��/)EIC;����\�=�;V�9�O��eHR3 �Yx�/�^�G�y�c$���F>��tA�ߛ0 G�p[���cN1o�%��M&�6y�R8~y%kW	��䋶}�^�����%���mu�,�<��`���/�V ,U|��x��-��]��'0�>*h�J�pAv����0Ě�*
pa�eKt���_ {�Ė�����/����X����O�Jir��Z�+^5B��4P�Ks�0��&`����:�3H �"�C��`�M
kT����]���"=�I�5a�}HH���f_�?V3�]��b����ǈ��q�����j
V�br�e��#Z�`�x䛿��u�Ĺc ��,A��xV�Y�XV�f��Bm!�׌Y��#"����D�a��@Ê}����Qe�Wٻk�f�L��t..j��5c�8b��lҍL.�N��ֵ��7��{�����in�dT
2F�Zw�����n����s�8&�`eD�����C\� j`:�k�8��S�$-HYVS !��"����Y&�����#J鼷
�pM|
Yϝ)Ʈ~���F��Jk�5iN�T+�q���M҆�7)^��ˑj�\7v4{��kB��
��J�Y�nK��cs�ʡȁ -F�Qv�Ѩ	�+�e-6q;8��"7�G��s�����$6�(�RJOV�A,�"��P^F�0��:���3���ͦT��
�'2��驞�sr	��)�,�4 ����{�V>����+�m�ps�S��Hz"T�M7�rh���}�޿�7�+�;����)��D֣�ばfW�k�v?IW�P���� #F���vB
�`�[��ve�\
��؅�va�1�!��~�($�46�ۛZ�G��oD�ɘ>��O������b��]�v�"�\X��9���ի���lDV_L��L��8��>'�0p�4���ֻB��z ��Ֆ<Zi ��jK�7\�G`��
���$���X��9 Zr�w�6Mԋ�4~������S��2ZB|C�$TO$��W�����9DS���V���:GS߄zdB��{`�H�M��$�kE���\DD�#x\f�66�"c
�R��"%YYQ�O�@L!t �F�j��\��9���H�d��÷�"��;��J!@��^�3g^��5���c	O7�F�/%�n�"��}%*	K��^�SI{)�)u�yqW��ǞJ_�����v�jW��N��]��|Z�ʜ�U�AY��ǀ6��F�ܞ���,	;9�^��l�g�m]�母#|؍�B��8���_����~�^M��eI��9����X��7SE�Sf[�9�PE���7�	h�ή�|�����N4[�zwR��z䷂���rVIpnAhو��5��jP�v^�2�Z�X+�<����ѸY�x���k�#�n���n#����~��=�.��+=k|^]�C	Ѫ�r%��\�pg&]�\s���f�6;={P6�b��c0<���3S0f���Ƞ����_�A�.�s��ڤx7�Zt�A��Hm_��z�����v]hx/dٝ�!DbpN����5�*w!y�L|��{:��m��&`�z�_թ~��)gw���L)6�k�[��$Қ�Ξ�ѱNxY������ָ։$��^�Fi�
��&���,�5"�w�<B��~P?؝<����*�,��֊�Ӳ���;Ɉ�S�]jյ�̂�L�.G�>��B�z�K�#ޕ�x�DD����\���Hm5|YI�Y[��J�T �3�O1�#��~����,�$~�=?�@֤h7�&���=�Ob������|�)�x��k��eGKxт�'; h����雜&	��\�7u����i�j�e����]�#Kh��,_�);��1�3FaXD�3t��ϡ�����+JOrQw�H�*�/��s�y��J0HDg��P��?X�Q9��=�j��FИ��V;X���v��޸��=��k����Ɲ~#�I ��>���#4��7jɣʙ���`�:~�e�͓nV�O^&х��Z�|كJmwJ�Q��ĺCK"�!P���^��X_�y�����@��C��\���g�J�bD8GqZ)��q^��&Crɑ�r4�`d���3���nu�4*I.�iL%��Q�9���:��+�tr�\t&��3Ũ	͏Uq��0�ܣя�D�Zf�,��)�m٦��rP��M������L��b
�:޲EfjV��,���,%� ��k������ޟ�Rz�D��V
��t�!�|�F���yggA3S�h �(�X:rh�,�U��ll�9dK��������6p���G������3���;Qa��'���KnۄS��n��r� ���5��{�	bhs�/�i�$��DN�@֮�ե�>�|�W�P��?]��JZ�Ĕu��LY�%�Z۝2�w$t�6>�����s��Ь�b84L��໽,�jA��N�!Y65��/2��Kdr���~��Yc�U���0{'�1oq�G�����o)B����glo
ֲ#C��'ӯ4UeZ]4X����F�8Z�ņo!�0�Q�a
(I���hY[#Hְu�8�Y0�Cgո���><�Mp�m�f�ǉ�~9�u7��5���Sg��xM���މRdn�7� +u5�����Y[�X����>fU�:ꖩ����vBT}c�a�c�2��xEb�QTk 3v���I�WʶE����ȝ
��L$U��5D�L����*�C��r�p���0f���~�щBRM�1KN�}�G��Ȑ���y�ŴwU�l��;Ϧ��3�,�J߭+�C���Wn;���O�R��W{�+��w�hvǮm���S�>%gzqA���g�E{���
�<I���.����DJ��J:�͌E�E�o-TW��U4�Mi[��X\�?��p˰��/�P��1�=j�چ��2����+iYOZkfN�/�:"�d��D7��k�"j������"~�i"��]1�|_"����#F���v�;"��hr��H�Ʃ#���r�����ք3������	/��c8L� �a� �UH��"�\B��&E�3l����}7�X�uD�\�����?X�0o�B9�2)����E���/���g<EYj�-�Q�lB k_:S��1̖s.&������y��A]|���O_���p`A�$�N3 ���M����ϖ���>nzF�}b��l^n+a��PH��=-�AHX��*+�Z	޼�����J��Ա��vY��\}ɓ�#����������c��	hj��iY]n"B~��7�ę9���R���2p0�#g%�P�8,�SpWZv�It������Gj��u�P)�J�}WO��?r�i�z_�z��N!� �=`���9nf����	b����H6:O���/�ܩ2tN���P��g>*��?}_.	.m�*��7k��-͙s"Ҍ�P"�A��I��S�2Ȥt ��*���e~�j:�itX��ᢗ�$�*���e�ްI')<����@~�ƶ���]������6F�����atV�G�.���@�di��B>]_c2lP�𵝎�/D�#~H�U�(t�V���9�13q�ڲ�V=��E�\���,��F�#�~<-�1�7jZ�D�1�%���M1܈P��Ie�%�f��r{�aR����I5�6�::�����
�pGw�}��
+��@�Ҁ\VR�E*db�R��^u	|w��ڱ���߮������pI|�'�M�����7S ���	��|�qB�|Y˼1������Vc��b��#��Y^��Q��3;M���,/��ݳ���"]$A��>KI:<ƶQ��P��kdބtfe��{y����dL���*�!K4Y��VۂF�ҋ�eSCHU��yo�)���E��Ճ��o�jQ��l�����7(%�xD%��݃O��4%��Z�86�2o�<�I�S��lÎeYm#~�����n಍��1�X���0���m��@�u`��5������6#++�q�D�!�an)W�v�|Þ,Jmb=>=���+�H��ٸ��![���Ԉ�b����kક���ቬ>��"Ҥ���cP���4;�g�7	���g���r�g��GYHZ��gq�'�o����8S�TN�ºZj$�aׂj�̠"k�H�"!6BJЩ+�tZp/�����^�k��u���$�^Nj�i}��#*\��mM	���{�{�
��)�/�E��RjVJ e�>hW���s�R��'T�Me�nP3���g���{Xq}(W(܍�E��C��k�Ւ�t91�g�c��l�,��CJNԛYa�3Τ������K2�ij6-�M\�u�1�ih���^E��g{D�,���_0.��1h���M�<�qͺf�<���y�K4�����.c�+r�qV%���d|� �p�u�IJ��� '�B�I�؞�+w�~�m�Q^�����N�C�ɥ2Y�c*B���`��	Vl����OZiW�(�����7 ˷o d=U��Hb��5 g�^��%�����*/�n�9�f8d=3@Za:�%�+ovq�x�(�n�ªVB!{|��׵t�_��0���DU�%/2�V!��d���;�-�����8K��E'_�ȥ=>~�.xՖ͆|�g|�$>���;�z��<��z�A�=y�dp��kX�u�g��ww�ٻr�66�9�!6�:�Fq0[��L/���;<K�@�Ʋ����!���� �Q9m�ŏ�c�l��?�F�!mq6a1���]]I��?�[�1D��~�f�7���`j�`m�;�5�aK$D';��+�w�[)q���`|Y�t��V�Ow�Q��O��q�5�0a��f;��̜��oZ��.��}����jW�F{]E֝�A�Hl���5��.8��$a���YM���6�����t����b�.;��O�y���%	��㻾`NT��J�g���}*r
)!���&I+F�V��d���1d#�������Y�Br(S�̿�ҥ�ѰS*Y��3�!g}E�ߐ���-m IJcn��C;&�p&����{���-�i��ԘQ���o�.Gw�F�����ޭ��k���AxK�6stGD�V�4��F+�������q�1�xPW�-!N��}��PrSr�l_���^ٝ��.k��^���.���JM��z�4�4�@��⣭�������2H�����cUt������2k`���;V��c�E��K1��~Bt�j�RFAЫ/���'�*�p������Ru4�����1�&|p�XH����/=��X �	y�X�z����gҋG��0ω�;tlxo�+*���R4�����~.��8z��3A���������Q����͹�^@#Es��%l|#*S�u����7�pz��"tbB�~��Ð��f�Ōq�kn���/G;���G��n
BT�dG5���RH��S`��+FS�K�Z���<R��{	e��o�w=���i�_O�o=��4}������X�gcq�H-�D��T�Ri`'�%� ��>U�����$����6gC,��LN��9)wr��y"u���+
�BΠmY��a�����V���Y��&��n��kE0�1w(NO_�y
5�(�⭐H��QAf�y�=�jc�o��JԺv	e=��w �(E)=�h��:A��Ȇ�/o����{�
�x$�Hf�=�n���
�\h����d�t�r�EuG�oq��Q��� ��T�W�{�Ĺkq**�[�/�K<���&5���<P�w��"��E���F�~����
Xxy}��VI���f~c^��1�{h�l^aؒl�EJL�F���@��A����4�4s3�mS<-4����W�_�Ά	I��C�',�|m�9�Y��I�����<3�W`��,�VJQ�u*�E��qĝQ�S7�3�>���#�K(��Ad(2a��4�z�]��۰�el����@� M����<'�hm)]E��v؈N�ı�����u/羻�P����AV�I�d��{��\���#F���4}����B�u�Q�Gk���@<uL�[�>���� ��8�R*<mv��>�f㼋��r���Q�OɇuHX�r��ז�}��à�k\?���� �}��7v�#5�X��O��˛:x\=�����ˢh���R2�.��R�Feg�@dImIn�hW��,[�&�S����t��X���O��˚�֐�V&�b�'{u�.b�Q�V��I�б��h[�8��=3�+�������<�V��%iBպvA�sh���R���ƌ��c֟�.�����3��@v	q2��ٷڂ�~e0En��,�+W�D���G_����5�0��?��EG����XU�ق��%B����*��z��c��P3���P.pxȁ���f6�u�
��Q�A\¾�Ku���J�ubaJ��k�H�@ϼIPf���E(dv$Q
l$)��c��U��ov��5~�&:��Cf��as/��*�g��+�L6��R?��@[�h�ⷔ[��I
b�7k{�X�'����Z)!~�cƑs1��ݪi�X����a�}�M�	s#lW6������</h�N�����<b!%`��E���u��$��M�Z�� �~�Y��k��Z�f"$0���gh|�SW$�@d��̋�,��Or� �N��;�3�=m�w|Rf1㷗�[{j�c+�w!�wӑ��G$
���r�G�I:�(�?7wopoK�Yv���%��	Ԭ�'J�M ��r�%�+�;�V�#%g6�L�ތl�LbJ��	�������SU;�)�P�E�.U����>_}b�vV򴪼��W$�@��	�6B��h��UƑ��ñ@˛�L��"�kڅ�ܭ0V@�S5�nUz9��JYS�֋��eIG&w��onӿU3	��a^R�@�޵W�UnTC�3�t��k�a��!r55��+{3w�����������ʍ+��/�(Im��!�[d��� (2�ѵ"v�������N�PJ�k:���HPY;��FQc�~�,jF�0����� ����^C��
NQyP�v-�lp�&y���Gzr�y=��@�e��Њ")�Z�\��4�^�*CT̻��F��咧��RJx�o.�o5�=�<x��ǀ�ն�,�,Z�{S�.�e/�QR  �݄�!�zO��Y�s��u��M4{�]�`�{=/�����r��Q��B�PN`^(�z.{�h�U�X�i���hP����w�+@K_8���6��X���o��%�T#��\^?E�MY��B0�;�֓������������ax�ԥ���C����#�dj�?�@�J��Й2��-d| pGC���`���&�s��|z�v���%��$�����U�E�?`,�W���
��xd��&��h��V��$^!fD!-�X�����`r�"(|C}��Uw��5�5ߨ{?:��gLD���3��_�N�V�|g�I5�p��R�)1p�5�P�]��g��|x-��V���m�ձ��:k��R��ap�+auձ��+��Ԡ2����Y��w���6}�
7ONx�@-�*/�e����r����A�9T��'پ���p[-r-��O�i����'���2tC?���$��V�����5�����ψT�D{�L8:�0C�e�iE<�1��aX�tq��uQ,'(�|��u�%�����*�#00���ޣ���L���G6��w��ٓ��pU���Q�w�|h6�$du��?ی��9��D�]��﷎��R���b�O��L5��<^��W������RG/�n������ڶ�`ڨ����ǧ�� �r�*#
��Z����ɰLm�Y*u�d���؋��n�-�\Sx��A`�x��Cv��ޞ�M8z�@7 �u���OD%�zor44!���A�Ť��%��Ր���T�%��Z�G�&1;�f�9�ȓ�dGI��*C-�\�ڴC�8�Z���Ȇ1�*�7SN���p�I�P���͎J���?�'�u��b���h^���%H]�(�bW_f�(3�~.��bu��o�X��.̻j����W�V���MLx\,�0u�|�>�\h��Io���t5#R��\T@�is�7�/(�c-+�Q'dγ���ur!�Y(�b���FU�.4�ƥ��W�����v��������t�Y��)�N�ܕ�B����ԁ�B�b������<�1�(>�8I����aok��������%���Q�r���edyk:�^�� J�ꖫ���^hϨ]'���k+�m7dA*��g�jmJ��nm��($���>�t*<]��O��(��lП]����X�EIžF?��NX��W���,�ki�4�������X��^����w���LFP�)�ohm3����
��Z�[��jF�}"%��u ��EMIc	���~���;��+�E,D�[�E�ؽԊ�*�M��
�,���#y;�bE��e␒���EG&�?g�u����p�sI���?���
f�	7�:I�D2�Ƌ�$��c��B����N3�Mw���\��n}cc��2	NI�,���h��Y��l7��E`]H� Ƽ�l�ؕ�v���qQ�r��_�v� �/1=�%��,�>$�]S"�D��ʵ&��<���_� ��NCvW�]v�k��{��b�xo��Va�D�p��CN�����H~,�v]y��U�w�������p�}u�G72��\�]�G����Zdx���e��/wq������xg�:�9R��gU�� W�=���|�龍��j�t
��0̐��*V�ಬ�h�{{e_�:y�]��('.:N���T*P	o�I��c"�|$�#�,�]��yM���*PGF���׵�����I��m�S�1V�v;'�r?�/�=�gMm�9����i4���U9�Saդ�ׁ�����2N$��ĵ�"�&O���DO��h[\����q�o-Y������	���킇1��M��]"X�P��9R�{&W����S	�c��6P ��������{��O=h`�0��U�!�*�avi�$/�ԃ�R6�-��`؇wy���D����;��%^�2��߳Ծ��]���� �=|8�d�����0Q˥�#�q �B�3��qao�\�' �&i=A��*�_��[h~���AM�B=��p��S�e����fE��j��J��Q���"�����4I�ك�]p�K��K��Vt���̀�g�l�C8y|j1�y=������������ ���~>��^���� �	;ZL�~�%f�^I:<�@ʥ[3���UR�Vf�}:�*Q9R0��$�������s<I�&�#��q�>��I�Z�.��h�����i�{�W�ML� a���P;	[�(,
O6���%\���c�X�Zd׀4���& U��~m��H�$���=����&B��;o�Sz�%���Y]5)��2S�q+�u�J��ހx��tB��hf��&��7�I$f��j���HOi΁�r��[FApWW�h{�P�q&�g{����FG&�	88�ed?�W�nu(\���M�ĀS���A�4�l�x��~,>!%)k�2�:�fiP]�Ϋ��:��f2��{���e7����ν=���l�I�6Ú0>M�)e�L���d���h*�㪧����@fg�`�Bp�s��M���ڭ�����u^.� i¤�u�����?R�3�[���cJ7M�����!ɀJ2��YU�$��1����t�v�9'\@���� r�tפF�D}�L)I�#Bp�F8#J�7'k�8��CY��b?��WP5��]n�
�H��Q��"j��!H�m4���?������ :��Rx� [4Ⱥ �����vN���ï<�謱s �wi��x���"���7np��hz����&B�_���&�s�ԕ�I�p��o�!�V��7=�O��V�+��(g3�ۇ)������d���f��R��olv�F�3Ln��r�֯��J>@��)�B�G_
�]�TH��j��֧�[ic��IJ���KkQ}��%�K��S���X��pGu�3����Sݾ�v..zv���<a�K���(�k� ܁�}6��(,�����u�s��?�|��j��I���?��Y&�ҲCd1��W�.�K��e
F�q�/԰�� �d��(s�&�Ū�&��O��1p�e��*�O�?�}���j�C�����>*`{샮΁���3X{��=K��a����܇ߞaN�.w�������0��X	�^62����Cz�C���<�Y�|� H�����(����g4$��"Ps��g������`5�77��������y07 \�ߞ��6�t(ӿ���2�lH��m�=D� �x�z��՚6>�ZIܲX&�� �?�U�.���&�$��A?j~����\�F��cC�8��;Id��e����dd}�D3��^6A��g�a�k�j�3�L^F�򎺁���t�8���d�籌Q��~G��'�֙��"o�R���.B�eLߠ�F�F܄w�imm)���|�bn3�e+}]��}�4ZKa��g0�e<��~������!���an\+����02����D�\��x�:���/t����$`�(����w�>�\XAf̋7��w��Lzl(�(pwy"��ze������ �6�v��7��~���.s����z��	�$O��&�\8�7��N~@r ����Z��/�x�su�e#B.��ۆ�Su��(�!�Q�*�]������ƅ'x�P�� ����H�dxM"�0p���*r�x:%�+%�^j�5�OK��,��0��*�9y�l��Tl?��m���É�o�w�%4i�\hG�x�(n�ko�1��݊V�B�/��o�W�Vi���۩%�99n�r(��T��z1�0���7U��f�o��3�Z�h���J^�=�ʃֶ�:{��	ΨO�#��{0NO%�j Z��4t�ԐR��\?�P�����{)�>��#�Een�:��U���:*�Q�=�O*E@�gt�na������@�H�>�~jt����`����ó�ٰM�`��^����:s�؜�G��|��ad�.D"��9@��U��&����r�r�?	+�Ҏ��i�P������81�:��5k(q%�L�����(��;� �N���U�N�����?�i��+�Qe�*[��l������������J�)�=&�k2���(�:��R��]�d<`��6���w\��H=C�S��s|b�lݦ*m�Nλ�Z���䣡�^7A@���}�`��W����69��Dۡ��WaW������!����4�ŀ>7#�}d
G;\K̘X�=�hб�	�<��>��rY��X�n���9���,�,u��Z��M��b'�B�iֻ�,n��&V����>�:��X�d?e+��=�u��k��� �?r��p^�^9�é1}U�HAf�:��s�(}Z����,[��K��� �%�KӲ��xF-E�`"��@kG�3��?Dg�f�5�r^3�Ѕ�j�M}!v#�*�/����1��m�Yi`;jEn#$���;�Qfl �)+�;|�� ��@ݬ�g�>�(�ERZ�<-�T�H��o�R)�j��%2���'��W�j�฀Z���c���R����u�K}�u���V	���s��3c=�Q��>;s�P��΍�H�l_��>Uc���g�����ж�[q����zx��.ی���9�rE,��g�n(����g�6�Jn"�l����(A$���ӝu�5w��©���o&O�X V��l��͸��gܷ��՜Nsz$���S���;�$�w"��s�>�O�W��)�S�f�v ��p�'L�T�"{�%��%����,W���LF��0ʒ��ՌbΩ�()ZB_�@|��D�&�}���b���>�_�x�yP#E�
�Xe�z�)$H���X�rɜ�8̑v3����A���v{�G}�qb�rvw�?2���F�7�+�x�Dx�(m���=�	��u�s�ū�Lܝpgm0�
l�.0)��g��ܟq��g�܏MA�[[!����Dt�	��Be�y�b=����e1z@#�̬���(4y�Z���k/�E|B`�Ӝ]���d�_�Q�T��7:~���|�F�I�2��.�F3|;*��_�v�exȅJTG�wr�|�Y5R�,��,�mNɋ!��J�<6��>�Q�5�A�ES�]�>�Cl�x3��t؁qa��[P|��XKrW@�;����BB}�%ǧS���/��cH�c�T��	KIQ�~SU�4�E*O�O�}җ3��3��������$����2�s�CL�m*n^��6TJ�le4�P�����X�49�Ħr�@-��3�=R�t?$I�ε�d�p�� \�>w��p=��j��p
n�B0q̯a�z��uənL�=㌢�8�nqy�y)<X�����VS:z}���C#]+hv*�=�\(0�uA%&�-f�<��:R����\�Q�B����Kn���Bn�'�;��mĖ~�g0�S�ֵ�\q�� �[�+p�]����',lP��ͭ_#s椽h�8J��-p�??���w�ɫ/������M��i�B.��h>�T��L�&�hV"��Ƿ��X���n��wu���%/ʭ��o�v)�b���.΢�Va���.���VǨ�mJCJR���P<.(� q!��U��E��T��R�;���4�GW0X��a�[�X ��	a��`5������o�@�I+�F����e��:������?���P�Ve~B_���R���;3a��~p�D`���m=�����|�Qe$�@� Nj���<U?y�u�Ll�%�U��a�q�dx���9�����@f���;�.Ϯ�B�Vv�i��a���w&^4^Y��g�:�����r�f��Ʊ�}���Z�5��bU'.�)7B�"{�mU���D�u�$��C�L����D_�+�^�36f����� ���A� ��ԟ���pʒc�|S(�B$��/��L�H��f<�g$]�۟<� ᣿ڸ	j�h�+
��Z`�ۏ�ߤ�17�h��V���n�d+\�/�g�=n2�9/���>U��$IB�͎��"�2�'G�'��lOP��\&���*�Y�,���	k��˘�����jfo����}�ф��aZ�3b�z�lRMR]l���V+X�*XD�3�6/�)�:�S�U�Ԁg?�_�2���ɯ�=��.0��:]y,��:�so15�w 5H�i��DT�hB���r����4h�#esO���m��Z�E9K�=��_ʆ����l4zj�ez�v�3�Dn������8Z�@����.��J�?IK0D ��:B����S7��  ����S�*E�UN���C���E�6���󀸞����N�zE��ތ��yQ�7�n��n�si;��K:���$�����=|��Ʀ��F�/�����:��G#���7~e3���0�A$�����m��N���p+/�����6����w�9��ӽ�j]�v���,���	}��?&o�r6���>a"��"�5�#,&�ɳ)�4��pv]����R����}�+��T����A?9\(#���a�q�P'����pu�B�zFD#��o����9�b��u�x���f�k�]'�] �db�U>�����D�����RI���a5��pqZx�/�IK�0>�B-Y������6�����X���pL�HYh��h&:�]�snc�R��Nϛ���歂�'�x�֌�S�ۛ��yDLL+�W%�����l��N����,	��4�d6���,Ӛ�������A�>���e��Hm�G�r�c�`��ji��7�2x����#����������ʉ�P��*z��7&= ���($���#�j�. {mْ��*����.���!�Yc:O1�ȹ�A��E�kR	�n���P&FI��Ր��¡.�70,���gL�Dg���XT��i*w��4V6��W�yr�b�i'η��AK0������oTy�J�TE?�}��49�F_Z��e���� c��[o{{�e��D�O�n��i^�����b-ރ\�PO@TS�A(A�Z*�^��Y��VDpW{Nk�H�=�A�� ��"��վ�A����AM���qC��d�$�$�V�J��m� ��7;Z�=�����|_F�6�~�������hLI�gw��K��(�fOڿ��B���������8q:1�M,s��m7�6x�'�v�+�H�����;V�r��|dm�k���P�Zz���u�M�K���:�%5�>y������I��s�7����(:>��K�R;��9�cz�Y{;}����z�h"�5�8,`�����u�?���d\'�O�&W��[FֽѧOI^X��R���d˭Mn���[�����7�Rz���)�t֭�@�̿F��zb ����V��yc�ۈf*�^3s��G����]��_?�3'Քe�F[�kg_w�hY�.L$�=~��V�j�LV�^���\��Ui�p:p���0dg��SH`�@��xuګ|ҕ��h���J?X.g]�ֲ�0ϛG�p��{���_�<����'%����s��\�k�Q�3*�Qz���g��hTL,�n�L@�I��b��\���v�q	:�����p#��P�G���w�u�D�!�5u��R�Esn7Ě���w�τ�=V����|񌻓�o!s�ef���q7-���� �|�ɡ�ӿe�B3���9��frMf�ݐ# �aޟ2�E��1/�'�{�!|�sB�&T
�2�$�����^�ukt��`Ǜx:��.\�t)�Ե���ͯcG��}��� �$�����)9��p�� e⊄sC��9p��5��tF4���k[=~�,V��փ��Z�-��
).ꕼmt����Eg��h�����e&lq/���q�,〹��2�'H ��wm�^�6������t����lY��zb��y͋�>;A���t�oXva����Ht��i�k�����#~>"H�~4�PgC�<����񗸘M�|�8�t�P=>������5G�����dg0��T�4��Y�.o���n7.�5ݧcI���{ez���m���S���2 X��GpNI�S�ƭV�1�s�9Aۅ|gu���@��_��1�Ʈ((��I��ŉM3Z�˲�A_�*�ݢ�g��[����B��܂�(8�$C�:q�˝�CSzS���:T�u���f�[Mz�^)�k��d��T��kp�D�P���Z�ڳ{�� �O�x�*E��_'����a�	&V拁�M�ךb��	�c-���,�&-2A����I��6���-��:,	��E�ڌk_m~Qxr�_~k\��2�%o���t��� �"�9i��E9�T-��;�^S �<;"�$wS;ڼC-�
03lqS�)�pau���G��8���)��M��\�D� ;>@H0��O���e@�W�򺓢;G�'��:��2�;�����ݠ�9# �O���HC�6�+�[A���HL�Y�Be��\��k��}�����A��ֈJ�٤]�O�^�#��������RXbQ)���3w�q=��,�9<B<����^�_v���&��S�F9z$1-G���y)�r���e6m

W�3ᯈ ��U�������.3VR�f7��7���_�3#L�h�l�~����pN~���#�q�=}v|�kCf��	,v���[�,���3ܹk����`��jX���m����JQܹ�w�ʸ�bw�^��+.jvc�]�,8wŧy%��8�罙��7�q?���8Lӽ�ͷ������M^�_�U\"�=�qv<�u�2ݿ}�HQ#�8�S���Gaa!�ʃf�D�0��/��i���A���1�	t$�A�6�f� ӓp���j�/	�Xy����+fx;��̻�����q:O�<FJ��B��my�I�L���*�	�Q�bϾ�K����aƆ����\o&R!��u�41*x��̜V�*��`�~�S�M
�S�*.��X��މm �Zf9���Ӯ��1K���'8�R��,�g���K���R��\7է�uNZA�P��'k�jG/�|7 ����;����5\�ن���D���O`���WG����� jj�(�A@�o�;A��Z���-�}��)q�G�㕱 B_(�f�<9��a��E�*O�`w�֕��[��]�ů��	���&�c"����w�3�/]<�PMٽ�S2�������Z�>S���i7@HV��R	K�Wf�MG�N����r��z-��_���3�5��j7�:UDG�_�I�=��Zp9�t-p��䆀}�ع�I�)?��-g�6)Qx�L�anU����O�VC�};SP���ؚ����Ƥ�2}��������^�ͤk��RWΥ6}��-�>�Ú�6��v��`�!�F��%n��4J���e���рG��(�Z^��vq3�)����i[)%�p�����������jz#	?[�'��q���kF����\(��h�3����-7d:�[���
���@���;h LIv�96=�|]�t] x���<f<�|w��p�W�,�i1�������b	T\�(u�������&�5�/;�y����jV~0��?�\���ݐb���O����U�I�y��>�CU���v?p�j��2�/f�{�(]��%����~�����>= ��O(
��k���f0O��KX��ڳJ�V�a�b�z���т�N��}�2!r�V2Hy��\7t�!�m���K%̷~��ܸ�li��3zƶ��%�$ښ���Qh�a���2C��S	$1Q�+�@��2^^(�U�s��*�\��Y�8}����޲qI<2r�R`g!D�q�I{���%6�������
t"�Z�f�9��0EMח���$�z����S�":t���{��?&9��i;���koCA�W$l�y����U)��2�t���'O���b)�������ڄ�Aܿ��k�Br���Q3�`���Ll|�~��h>����u�/k���-"Rz���k��Y���Wm/,K��)^�Q���-GY�?� /#�3�E֩��:؉�-8/3x���,���!أ!�(�'�����L�i�9o�
@��Q� e��e'~������'��/�f��30%M�s�h2�wWd�xe\�7�Q�c*���7��M��h$� Z-�]�;��6h=�\�� ��/�5��n��u��X��$� ߧ��E%UdG�`V�1�"ݛz_& �An��?B��U�PH9��I��+%ހ|&�&��J�sd`j���z�E��J`����(��T-����p�p~A�[ň�i�f��EZ8<g\���;6c0R�g]�+��C��E�%�Cn}'jlwt�[�̻Q�Vi���İ���Y�oP���j��ة��2��a��j�����e����w�|��r��
��Ω�&�ntFӖ`mg��^�0,e{�U�?IC���{��<c�!C|�v���X��t��ZP� �0O����qB2��	���uŧ+x`ɟ������\"T ���
�}э�s8�+4�_��t����B�wE/k�"Gi��4^�^�b�Tⅎę\�U�>�r��W�B�{Cq��8�{��R��ߔ�>ID�_-P�xX�OO��Զ�,Ј�ݤ�ʐ��� *��W�U̪i��z"5�r̙��x<�R�����2}���?tK^7�.�P��=�6fL�Ĵ-���0���"�EWG�ad���w*�f�G]GLɒ� ZB���D�7�ŝNhZ�k=�$!��!�ű;Re_p::��)��c���K���e�\�{����Q�FP����1g>N���H�5Asq�!��]�*�a&E&yP��������j��ٕ�K�.��u�<_K�� v�!�t}������Y��Ug<����	�l=�q����%�&�� �Qd�wÞ	υӢL5Ƭ���ǒÜ�y���X��c``(F���@�&�����9�6�)�M��;��%G���^�M6X2���]b�	5�C��_��W��+�&�[�~2F����/a0q��w�
��rQ]x��dQ��+t��x]����8��\t��vg8K[�d�	$�>����U�* ���a&O��]��-ׁ<fZ�r\���֙5(x��"�r$@m"W��~q~����e}>�_l\�r���*oQ��*�N^!�6*��2y撧&��O�`�$��p�zm���_.`�����ߗE(nB�##��{g���N�=f8M�@�eq�e�ᆺU�V�"o�&�Z�H���(�QL��SMZ��8 �⽬��b�K�LPp�Y[h�8�I�����3�0� �B�6��-��;"���ֹf�h�2�L��-R��kj���1�R�A���N�ɏ�=js�H"�z�S��$���k݄��E+��i�����,���v�Jr��Ϯ㽢���B�M����I+z����T��Ǭ�J,� �"j��x�8DdF��E���V����7 &j�j�}p\���m̭�V��J��E�$�c��W�כ���ƿ�b]� UA���[�oc�]�3��<�d�\U�A�Ddv�`�3>�J�$�ʍo�dE�v�/$]�<�c�2�j��Q�#MjR�}C=���9r�Z�r��jTEiB���Ie$��ib- ��}�Q�P�G�ϼ�İ,�*�W�@$Es}��x�&]��ڏ:��L��*�u��lR�Eq��������f�z C��?�R���bYυȨ�f%_6�"�a19�3�@!mz,G�6j�Ɲ�0D�h���|�Ľhu��M�6��PU�/�_]��J�e�3����'z{�pS�
U����l�r�@�k�Pub���Si��n����f��e!����<�Υng*�����/�1u�_��+x�dmօtB(�'sY��B�+��=�_�z"�2�Cz}w�/�`��lYK�/-'�]�K:ʋ�}b���ü���Ta����L�lA�TḅR[&��#�g�=��T�Ͻ�1��K����N�����؍��=���b�+�
�$B�= ���g�q�7�G���D{�bS�InN�ID��ݒf��!���������w����(��Q[�.�|l�ӭ����Zx\�����q^x�-Oas�~{�����%���M�+.~��MP�V%\��-�+�
=K�sO��[@2�d@�'#}�2Lɺ#O9�i{��oi���28p<l�H�B1z���F6�ǉHh�3��+��]r ���>f3Dq��6��PnrnQ.3�|e-�����W���_n��X�.��6�m�:N��+�&�.m�<��+R����'�QB��7|�#4�!-���ֱ��U�)>2!v��[	n��C��G�,��a1�|Ө�qv�:�����T�'x���l�G���f���D�_���'���M �a騬9�1Oa8��󿬔�ޙ³X��|�ުX�Nf ʧ�FM�e��<�QUJJ�L7�ά#�+X(��T4��ە�q�F�	���#~(��!��mR�8H@z�0p�Y��sI���VjR���	�TFp'���,D��>�M�y� ��a�o|^'̥~�B��Fܤ��L���&��a�K~7���f"o%WB��DX7/]q�&ʵXk�t#A0(��t��;��4$u3I��#��vzb����r�cp�$L���(�B�Hh���B�v����bXr���t-��fwDGMQxu��̊�![�g�y�`5`���#�z����ܧ
�ڂF��<��o�~u�
 R�Jnw[��ԙ��:��{��hCUhGɲ�0����}��M5vi`	��U�X�@�,��o��-�P����ɇ-�%RMQ"t0~�Ց�)�!�#6��XX�u���U�n&�Ӏ�[u�O�\Bꕶ��1�O��mv�������l2�~�3�L(j�T����d!���r:Zi�,P��E &8�xU;��J��*�"��l��H��|���9�
�n)�����4�ظ聒C_�q�G?z9�C�Aܱٲ㟎�2���sO�{�~s��/��gM\�%��6$:H
f��Y���A�sV������?��@����t\���Y���,�L��Ly��[R{��d�R�&��v�.y��ޚXZ�aM��AwY�T�r�Gh��I�a/j�����3�Giy�J�s?F#�h-��iע�P���A--w�i��	�7Δ� ��$`q[������c5������?�88�>4���:���b@b̹�c-ı/m�-5�WƲ&�;�cy��7`�OJd�jo��}�4C�9�MU�r�jy�4t^�����H��}x��]F�U4����W�f����Y
.-��6�����⣿G�I���&��F'�l���61λ��.������
�F�_�֝c�������2<2����G� �(�n�?6���lR����d�_��C���&��w� Xχ2S<�X��a�H]3���k��g��|>�qw1��y���e�Nؿ,J����܏!���-K�;Fi�~�*}V�:�q�*��,��[�pj�%�]c��MR��>v������'Na�&�U4�6�aޘ�CՁ���p�b�ďf��R�� ��c��_F���$�V�.v�����s'���p�>�K21,ę-�*Л�丽��i�W�8�3Ǵ��F�=�#?i
g"/��3���.Ee$LZeo�	@�����?Yi�-A#ޜ���v��|�G#?�ይ/��Hi^�'� F6�o�I:�,�!����3�gE6�Y��L:�j� 	0��޺̈!�<:R�9(��X��{0�����9y`�a�d�zlxp	����k�W��[$�����n����b�έ����3����/��Cd���}�����P��0���S�x�a� �z��� 	�u��R#��2���(�O�4M��a0�5�����F��JuX��>��uI�G#
Wp�QB��[�Wyl�\-P�/i�H#��[Ҷ��`�+<0�C���\邎�ZS����(��X��|!��=yV}�����=i��I��t��a��׺��m���s%={���
�:�S���,����6�>�B]`��+)�����.�a�r<o�Y�!����T�`�+�����˲
O�Q0;�k������)��G����#���u?���^�4���m�"!�H_4�MF�e��U/з�ί�к>%Ta��Z�ۤV�[?-cz�5D�J ���F�(�^��6�1�ʢ��4No�zЎ�S��(�G�Ω�x�%�8+���9�J��u�4�M�E�z=b�r�{�J�3�%*��'GXO%�gj�9������VS�.��e:�(�����Z?��}m�k�>JM�7���z>̬(�B񩇘��-R�9c�7��OS�_ T���֋���u�"�G���S�ݽi��N�G$�%�а�K��CR�l�3�N�^ԁh���Z'�h
�^��\m���1�+p�%�N����=O�(�vzy���^��*�2sFT:�G!�~��>�G_�k�0b�c� �׼K������j�%��H#O��헠"��,9�[�y�*D`D��5|c=iL	AKi�yL*t�UV�3��>�$�Aq�\��kf��4T,��;���+��ҽ���D�#s�[*��z�X�nb�nu|O���m\K䙠g����&Z�u������D�,�-w�sR=� R�#%��Z�Y��95V�A0��O�6E��.�-��$�5���L=�:���W��΅�V��| ����a�x:��l�q.Y����6�s�OG{}�6�a�jo�����H�f���P'�)bC3�>��Wd��L������0�n`]%�iz�Ԥ4��ĝv��h�y�M@\P�^ l�E*=�l����/wW�ݗ.E�9�,���T�з��̅�v�O�6�Q*s��6��I"]8^8W��A�_V8�o?7�p�9�����]�F�(��UJ�����X!5�[�g�G�;�t��A�L�Z)�<��}h=%Ӄ96I��R�����$9{ɰ�o����;���6��p��v�7��֥/�T7���UAe����6�:��Z����Z���]���5�.9����ug��D��o��$?����ax��i�O~B�v89�:K�P��ޠ�e	5�rҭ+M����4��/L��00������+��̚��\�w��9�n���R�K����Q�w8C���b��M4Dd�wQ�R�f��ZXP�]��f:� 2�m&N(�m���S�)�T�<�<�Kx[�qƼ�/�ke߯|bE!Aꓥ���nO�ʚzY��PP�AaPwB5PҊR�4T#��knA5u�x�Ȓ�J���d	4
�#?m��k��;4�l��(|X{%4��!7/:h�Of�uvӬ����� f�Hmqc��g��{�ȓk���;�b�п�i)/>!rp����{-��*Mm����!��_���2�gkM�
L#��f�H�,B8\��E�{9��Bӳ<c�Ȥ�HA��ۣ&Fl.t=�M���+(�s-��4}-%Z����Zo���'ƿ=5�Y�&�t���X=@&J�c
�%7���u�߻ˑ��fn.�G�h�]tYJ�f�'�Ybpl�A��6�8����rC���6�0��c��+J�=Љ���Sq
S6@w��7��ţ��7f�$��"��4�d�6��O��D��]���VkL���J��+iV�#$z�i�KU�nu
~�=|���,�Q��l��i�s8�a�x�Iz!!j{��]�=�DVfK����Q4���˳��3m���#���)c��z$��)�� ��}ni�-ʖ2\k�-�
]�/2@��<N*$�^EaQ/v�QJ�mT�Oy�ja},��"k֟���ط�H/O�\L��mT�j_X�β0����UHq�Y"���-r7�w��Y�!6 ��9�������P$�@�d@�a��^ ;^0
'�~��o���+��o�϶ �ȫ5���]���Q�|:�4`&Y1G��5������s�+���\���?0�gKL8WU��;�rAC������[�f�6����.'_T��(���*hM˔��>���Ոb-�Q*&~ԗ��a��ʑ���v2�lg4��
�/��F��otՆ�;�][��j�ZѝV��� ����O����޳7O(�lzK�~���y�����p��91�j,�R�k��q��:!�0Z�x靭�Y ��A��bKݿ���Y5���Z�P/
��l��VyS�9�׻T��EbL����c����.�*w�;�Qmt������CA[êx�ɐ߮N����7��FC�Cps'4rL�%��Ff�B�
?۝������x��� &�4�SM��|𽠬۫�< p��7�	�[�.�h�xƿMv�Wأd�&�
`�|Q� b��F%F)�� ��I�i�b�91Ȱ+aKk:��u������������Dp�9�C%D
���~cU���*�J�B���j-/G㘵�dӝ��uhX��w嬙ڑ�I��:�zg�lz�J�r�7j��?R��*�
G�S�f0�N'�9j!�#�^�$N����ozwu�N�.:�K�߫L��AQ:���ޜ���3�mN�Ϳ�s]��X������b�$S�
�UA( 3���\`��g�h������z����:{-�gj�v���D�l��S&P|ԗ}��~e�p�Գ�9�t�c��=G�O��I��|�؇}Ui�
�˸/��!�	k&Cp��O�D�\�*���s�M�y����:e�����H;b7���M���dӌ#�M�����:M�P��J�NE-|�W��n��/5fD���=$j��Q���Dr�@���)��+h�2����7��&؎,�E�*�IB蟇��p���~=�����[�X�nDc��(-����سΝ=yh�-��}ׇ&� �mØ:`�v�ZC��5ɴ���V"��������aH�̻�dw[�#��/��}��k*(%�Ki�����E-��6���ğ����ۗ%�|	A7޵S�3�;�{�=�|��ӣwo��:���SL:N}L��4�g4n?W5�Lj�Sm�6؝߹�
��ٕ�?�9տآ-�1���Y)\�b�Ӗ{ ,&��<!�b���Q��$������ܘ�-�xQxf��ۂ���'��L�th���(��[�;�ň� [�u߻�M�rƝ��?��r���'�H9ۭ��Y�d�� 1�=J�{E�I`����UB�2�k��0M6��|�|��e���	���M�Ty�-�K2�kl�X��y/���:a�C�y!�&�r�ns��⌽e�� �����!;��`k�/q���Ḙ���Y�n�"~�\��sG<�&�WR��<*� 
�?X��>�t�r�L�,�Q�)l���"7���2���H=���)��!=mO��������Q?�d�[r}��I����gVL��j�Y���2�:^�7���o4 D��f1Pj��>ޚ�_�W���e
�U�#�.��L)����E��k@z��Et���A�7.�(���ӗ�M�1<�J@^`-ܩ��Kyp8B�F��:�AE���Vc����UlЗ�h�l��3E�)���R���PY�I(S�'�+⛐��I�Yk"Ʒ��f��L%����/@rV�2�S��<�^M�XBq\ �=�I�b���R����
a�O�wX=0�=:���(�r�FJ��}�tnYL'W�d)��|\YW�bWW�E!e��1�e�/Vpܚ1�vxw$E;���|\־�Us�"i��#�(�:��m��N�e���j�BU�HO���+2�a�<-]n;�IM'�Ж��}�������1a:g�{.d�k��ʠ��>A�Ci�	z冃���t�@۫&��m�vv73�܄	�<��P�Z��Ml|��M�rDjG
�'�yš�8m�B[n�#��Z+r�V���C�xJ'�|<f!�?�
���U	����� �S�4�I�m@R�*qd8�/X�t��'�8-��7r��X���zb�e��f�ζ�M�3���Mb��:`$�ғ��1Rw|ʍ��yjo�p��pm#%T�9�f$g�ul����Z�ӎЂ(e�/�ؼ�Zf��%�c�Q�6`��� Z�ƲG� �b$Z�v�-���_�Ĉ�%�	�����&''����aa��������#���Y'x�h����`�{�B���^�ς5����?  �pA���+�	6^))p�P*�g�fߨ�uM�9��u\��q��B����t����������C��|)�s�&!L�6��5W��cڴ������&�a��_W>/ �W�蚭Pt�fS��J P�v#�5^B
,����^R���ɳ�U�^�#�������L�*e`��ʜ���Rk�Td�	H�������mۡ].^��IpC�sԡ�{$��� �)�W+r�Q�ͼ���~8���nz�&�?�{���Zmm����s�P
b^�M>��ގN�E��>� [����Y�i®:��7��驈cn�]�(�*﬽2����-I0��4��
�cI�hc-�T�#+�K�������?���?��c�gI�9�6���C��;��o�]5�Vh�!���&U)g�Nt"�r?�B��@�*:N9�iEv�N �=�����K�I8XICl7��[,�V�����X�LJcb�`��0�zn}b��D?��-LoBo��e>l %G}�j���1T2�� Y�K���\�bk褝%�V5����Тy|�HV(|���A.�k�u��N��ɵћ�txW��1a��b@Z��������D���&kVY���[:L�G\����	�O�Xy�C��-s��cߥ�4�74��V�KVkB����MB�E1�%�~����nL���]�c���3'�N��Zệ��̩q�����Q	k	ÅTX�0��=0i��1��K�e�4�D穒��o߆$a?��׫�w�}-M����&�+9�ϓ2��Z]QK	iǴšipz����E���ꋫ�D���R�~ń(��+ٮ^�vf�����Ͽ ����W�׸�*	:ė�i8��+G.��hM.������ 	�<[�mn�i��%�|��	��E�0�bW+-�N��h�0�k` 8��q�.Ћ%��#y���9Y��WA�g\8���	mщ����l�-���Tz�(ׅҙ��H���;?�!��P�@�<��»�9�m�|��w�/:�qr�!��|��q4�ŻH�j@ʋƖ�_�e��L�GYt �љ�� +N��$��\2������?ˣs/X������݂�.l� �-�?�G��ȫ����U�����C���0��O��j��o�+�[�;�m��T�?Ik���%�!U�F^�`Lc?�^������
T� �C��%R;6����$j����E�ݿWo�%�\3܃|_-���&���ҹ3�]?",9z?��|pj��CH��H�R漁BO��LʱA߾_�KD?l���d�k\@'�>�k�%�a��3��3��P<- �SC�L��69�c��U���km`.��ƈ��$b�-���S�&c��I�f�@��&����$�0��_�ȩm��1��V�t;�kS-�el�\�l�1��|�7���6�l=�z���6�y+�Y>�a-:-�p�\PWH�MX�t�J�<σh%?���{<!z��!����x���A����b��)�Y�;W�^��fi��a��`�D~AN�:}m&�5��@�2�:G��
{7��I�&�Q�]��Y*.�zƨ� ��%��E[�&G̡��n�~R
*�B�l=�K��_�F�!��Bel��_ ������l�#@�맸,�gu�n��6z��0�"�E1���BTܒ�������ϡ��;a"�Ƭv�o>p�M�"d;�x�[@�Q�q�l۴d$�:�AAQ`��$r�x��y�2�fZ�Do�|Ƽ�@��<%� ��8��@��C�?@z,(���˫=Ba�<�����y���y��&Y�B{r�d;����*?��c_X�wM��/�@��
�kaܠ>9ȼ���e6����sܑW�K���..)|�$%��$�����GH7[bܕ�-o����ד�3h�v���ҏ��]d�T1C9�����;����r����Y��~��0&U$z�](>���]��)g=<Y�!���R�Q_��
j0��p�aQɸC��"�Y�-TE򮿌W��[?37�h.�`_⎵��_^�T�j}0��p3a�G9Z��'���#�4�3��_fF.lI:.ȵ9fr��W�T��Y{�S�.�[��c�[�����!����T�50���m������JN��e��-��4�o�9\����Y�=�U*� ����4��H�����۝@�Lw=-��E٦�R[���]�L��*b2��R�4VVHT�uM.�o���d���L�=I�OM��l�n���)�+��2�s���q�E[��7�j4���R�5��xL�������\���>�M��h BNr?�1$� ��>�+F������z6�{��QWβ�O�v�:�����U}����$��c���4��� r~�<mV|�~>d��o/a�5������On�� ��,�WK*��_��8ޕ	�,�&���.��<� �R�x@?��s7����J��2i���i��WϜ&j�
�x6��<v�=,|K	e�k�d��y�K��,�V��V�!OJ��/�4�byBI�h��y!�/�h��)9��������A�J��c�){ý��S��w�GY*D��\C�"�f��JZ�D�\� N���4�D���ˋ
tX|.����>D�(A!����n��}���eФ��Zq:� tI.[R�X��7C��Hٹ����r�|}ր�IJ�2�Np�l��0�rR�1p�+	�N��6�XZ��g�O�7��x1=ў2�%B��z������.��.��gVJ	���
�u�.' ��ı;̞?Л�P@��$Fv��߈�#ݖt(o��QzL'������ںZb��~"
�����`���[GtBd�(&��Y�0��a��	 $c�iJ���
�bH�E�z�%_�6WF�h#�~����+<�"�b�{&|�h�.�s%��ѫ"
�#����y�u��b����ׅK�>n��儴뚺^_����ڨ��U�|f�r�-5h%�Q^_c�V�6��L}+
�w��9�`H��Z?���p1���w��H3s���W�h����~�K3|�V/xD�Ի�I3ĸe��CJ\�QKa�~&oH��'�'Ͷ���<���I���Zv����Z�֢e�Z�^����E�nwCT~X+�o���F<��	��@��k�_-�˗K�ô��� QE���Ȑb#e�i���2Z~v;:ҝ>Ơ g'��u�C�,$�g�l�'�z����1|�JJ���[����d�-�5t���ЌsL��o�E|�r�U��F}����J�������a7�˯ǟ���0�:J�3�O}� �ܡ!c���K����&��f�{#��$O�R%��;m@[
 {���)q�������ҧ�/L�
>@�䡱����#����Z�O����Z��Hf+�Y���*Jݐ��'^{�6H��xdBp�w��R���ߠ	!X!����+���x��@m�XK4�B��~fZJ�IH�_�;��9�y3Idj+�9���\��Z�v���={j�y��,rf��y��;����j2�'����A��nJ��~<W�"�'�z2x>�z6��-P*
�:�5�-�w���J�����0�:�Ҹ5�����N ��&���j��I��N
����!�q4�q0�{)�P~��৓lM�,	��S,h��+�Bi��D����f�av�E�թ�^�$_�,�T��$�_�r�'�(���ƕ�M�Q�����6��ʇ�f
�|~�]���'�rmӘl�=�;�v�R!��~�_c�Ex:����'�V �%+��Ų�N�b�fQ�\Awd�<�kn�\y=p��������Lx�I����l����ln�ML}�/�.���IU[�4��g�c^�p�[	�S�j�l�0�6�*
��n5*��M���h��x1%u��ẋ�R������T����C�D�,_p j�X�?����{ͷ[Ϛ�W���V�U�7��� Z�����}x�D��-tP�m>������w��9i�4X�u����%�5dU�"��}w�a����A��V��E��u�����p;7Y�pYԂ=,���]�=�mjf����� ������&�bI�U�����]�GFDa.��wKÜ癹̳h�化N��GH�8�b,��?F��<����ل��.?�}>�������̋fؐ��0��wfz��+��$}s.����[��"�;�)�	˕1�Cm�h�}��G5��8���R�(Q ����b���;�#f4VM r�y��)J|���Ofr^
�2��t>J��dͱ��|��ՌF8�?`iֿ�n̴�3}F�g����p�
J͜��0d���Mӈ*�L�nT"Q��ʡK��$�MV���/�B�D05��W�O[��퍢N�����">�^I0J���k��erն�J��4Գ�|\���t-�����D���wO��������y@��0#�'&U����"���a�*����|g���i�0�L��T�T4?�.)�
)���د\��+�Lh�TW�Q�˖ɰF#���h���x5��(9L���.%q�� �q�
�1�%vy�u��wm�wW���5(��^l>��j)+B��p��B�
��r7d���0�p���4��5;`k��L�R'#ܯ�Y�t3pU��v��PV͔=y�׽����C���F~����e"h[z�G6���*tG�~R�t��fU%����s��~��%GO���+NPL����w࿪������e}��ۅ���24ˈ��]d=�����>���j�k(-@%{��m����_�s��_�,�s ��u���B=��O�ר���|�n��yy�~�����F��m�Q�A�������<y4�X(��6x-�V�ul�x+}��6@��;e��9 ���R�=�����&�;�S�oS�-�ǎ>����eYH8pc� �9��*�K/�5-�
:�[q?{8i���=�%�(7�i�(ė{hK�Ŀ���%5Mg��I�����r�8L�r�$h��<��o��LC1�`�M@�o��j5y��X��I����'����MX�=�7߸�}�4w_��2m��!�VSc�s�q\c����`� {�R7}]�N&�B��,+|�F�a�ϲ�g��S������f�̕ �)5HME5�� J^���'�p��h���@�y��f���;��z�^�OY���NƬB�ߣ���S��
J�zP����9R ��)��y�9�cRV����/A���E�y�lfw9O��0_��%�
B��OD���d�i���買�BR��b@d��:i�6�O|_-4u�Y��o-��n�#�͛^��j|��K���ME��9ٻ�j>��F��N�PY9=ú���]Yb�y�:zz0T?�tve�Ou��LV�$��Wm��H�@%k��E`E�}���~�9Ǭ�ŵ����n���u'��N�N�t����u�~����7�dm���� ����3j��u���3����s��� ���LE��.�^9�����.6��NG����=}8�v��Ϡ�Y�]HZ��QU����IVg���O����ƍ�{����Kx�b���j��q�9l�������8�J�� ̹|���h�x7�%�O�DH���*��X�[�tu��ϡ!�7�B�' �.EcO�v�E���S�*�Ek�d�Y4��t�wƇ0(��s��f��~t�n�a��ۑ���[���Pm���o�~1����P�'~�C˙v�@WJ��x�ahJ{3��ּ��Ն��7�"�f� A'aT�ރ��'i z�G0G���Q�)2���کܐ��9h<�GC? )�m�ڀ{ݐx$��1ja�>]�<$�L1�a�:�"�荱Y��I��?�'�X�ޑ��#w�����:z�����#�' >
éN�a��y�(�]
�9)��b9�� �נ�,������"����5�PE�U�/*ȇyqaH5��qKF�{�׉�f0p�i�Qo�?�^/�ˁ�x4Q=�q���m-8��1w�z�H"���A	-A�]�Ò3��F	c���{�i���O�de���t���J�aa+�>#WT��GG�J�z��.[W@�t���#T��#����'%�幌p⒑b�����.�� �|JI*�Y$\���sJyԆ���W=Mo����:��<��?ęB��N�s�Ob�v��U�|y�F����y�ʯ���vM�Hob�n��|Ђ}�P_�v~O���<�l�J��iO�u��1��>\�����P��-�ן�Ч.�u�Q�!��+0������g�����89��1w�~��3RB�Ô�al[��4�17��1���#���f>�Pgnc{1��?Ql��Y��b�6�#zQ �B6�k�l�:B��^�;i�I3U���t��]�ÆuY�ʦ/�s`��O�
���t�G����i�V�Űd!��(��^�(�dl!%j�HT���*�/ۇ9S�$散��d �]����D��5T������P�����"�%Ny�=��P�`��#�E���A>�V�;��B��ğ� ��B�j�RlL��b����~��2��=9?���"d	��&�X�VK:dc �9�#%e��kZ��Ê�p����s����y��ӳ�ț>���L�f���̓�ۤ}u~@�;���x֊ԕƅ��ȂbO�������?���9a�;r�$�������7��Zʋ~�_@����{*o ���w.U��af��������x�I�hZ�JJ�<[�{���iS	j��L��=��RQL$G�2b�[ZU�	��R<��<�Q=��74�r��7S���W���*x���A1aĂǧ]�ڏ��
�la�OQ�.ӮJc��!�34J�)Fc���>X��dx��(�OT`9|6-�&7�4�nu��9%�+�1Z@ī^�}���RȎS�`��S��y҂*�w�{�>]z��B��_�m�v���[�޲���dS��Z�ÈgA¶C�Èw�ƿ���Ã���:j�-�D(����pN���E��8e��ύ�S,���>����5(�!���!��6/�$:7�2��$�Xp��T�����=`����]; ������^\:"8mSڎ�1�@=l��@b��ț�օ��)�N�=�)솅G@`�bd�1H�+�;�c�Ϻ0�e�c\9�<{{$̷x���d^V�10�yi���>I4)�^���.���T���[�r�1�嫓W9�6�f��"ۛ�O�d�E���li���	�Q����9���d^�^����fu�w8���D�(1�sǚ�}�NzO�ź��������y�\�x	���;��LV����<]<@Њ�Վ
�1{'{�HM��O���)�
��vө\ �V��B�]��J������O����kU^�7�d��3��SސWbw>P~���|��<��N�f���F�z��I�o�\
�t�9�9C����H�t��a�{��Y-�ץ~�|���!J)OFJiH4�|�7a_��P�����Wo�p��������(�B�ȮؾC���ˍ����W5��5�2���)ڄ21� ������'��Y�S�����9̽w\�l})z���_i� \@)��I����t�"�G�����c�>�0��*�|���W��o"N���fMq��IE�Z"ES��ؒ�`ٷ�ƸaAr�Ϭ0��:�^�W��d6����SN�X
�vZkA2���dސ�{��bB���2*L�oT�A2�Dwt�K*G}Ȝ�(���J��v�خ���#Hq�'�=MQҭ�3a��d�n��	���UV
��6Y�[_��ٺ��c������"pG��M���sY.�a~��O(�,k�LNB��揵U�GG��s��*Rc�͡v�F�#)@#��(U�z�Mݎ�(%���h�+6�ڧD�sD���=5PCZ��ç�h�q�ބ
�N���((���l����Q�G\0�����v�U0Т�>�b���25O6��rx�M�z��b��WT�J��bb%T��\Y��b4":`�u��د�fÊ���zgQ?��X�o�g���jO�v;u�,�#C3��}e~��!�X�9 ��8���5%UfDF:5�pQ���/È�o9�����j��T�L�_)i�pg�~�C�+���,��
��6i&��+�����^���$�S����L�	3���q�,��A	���}�S����:ԁ�\���F�SGE:�F#"��݅0`�̥Ƕ߯�<'-Zb�K��}��� ��u���Yym��T2�w�>�{K*G8�$.L?�I�׊L��0+<ߔ�4?AK�VkE��0tb��:�����cVF@�sz��b���v7�Cu\��i�
B�J���:_ܰ'�{��Y̗�ґ;)#���A�Ԃ���x�{sѥ#�7�UMAY�s�e7�J��,ّ�fs��8�cÂ"�bJW�/t+3���$���Y�������������C�ϝdv_�^������8r��W�<�%$���S���'���4���k�����%�{�Pk��Ȗ���iL����Q�A�8�L�Z��������l�HS�I��N�/8���������<�����B�5��Ȑ{�t��?!kZ9��j=X�:P-MIZ�le�O���=�@*-��g�{�S*a�g�� 3��)^�������
f'�ֈ�[�M}�V���&�$���\3� ��o�4���1 \g��4]����R�]J��{C)xz�U%������j5��Ʀ���7��S�R�s�Y�'O�ˁ괕��_����L݉��ǟS��w��/E���N>EE%�{������gf���(��y��T�S��=�D;{���[���,�鞹�;�ˠl�f��1�^����읡���fԶ�64��L�e�3�'�1oi�/�~A���F��LM99d-����;��"�lsi���M�ع_�7�?ē�-lFˡJ�����ND+��uІˣ�am�}*���Q�m�!\lc�lg	����9Ϸ�־CV)	�=iq���w=q��2����{���kDEebE�
�~�ڞ�i[����:e����u�y-����mw��b����^�7^���[KװwR�3��:�|�C'����m룪�%�?	�&�"�o>�t�E��^�`E\��Y4P�$`k鈪Yeo��ӥ�Z�������*����ɶn��+u�>(s����|�x�I
����{�����_fc�G����{��~Ij}�"N��s迦���We��`�Y�U3��?�D�=_^h( �%��6����%,����/�*��i���s��-I��\���uُ���m��S���"����~�_�нB��\8���p���j�ߐ{�q@�� �l��Գ	l��tH+�^o�|��ˋq�,�4)ea-f�9<�뮿�O�7t��Ӫ]dzZa��C>�X��s&рf�!�0Xn��?_X�Q�9t�Mqxm#���jP�t[�b|�	�lg��U43��o4�Φ��#�!X�%��C��:	�o�D��+[���s��͌�9�m�M��>�.��i2�yɠ�վ@`�:�2u��(�:xl|7��y�ݩ-y�"�/�N*�#�۳Ⱦ�Kgͬ�<@|6�g�%��o�$��vl�!&��Q�q���jy0�NG�K���Tw,�v��y�yc_c�+�!��6'�	ѻ�T-NK,Juq��w��j�kz��{���A˷�
m�F+�[�%�,�v,�ѕ�]��9,��ӈ�औ�I�]���k F�<^I����L��h�	akQ�I��X�0]���%岱]e5�XqՀ�Q�Ϯ�����g-T)����������> Qߞ8j,���g)��� Ⲕ�D�jSV��V�W��ѱFF:�:u�����|�z�Yra��Uk����|!�$�
�Rr�It)�"����v����H�E�E>��nd ��UG4���/5�A�ҙ��U���t|x��:���)z��_[���ὺȵ��.�$��tImW S�6��z���
T?^�*��PG	G����]�/����"�3m�C�:���|0�� ��� ����`�[�Q�U,Vy�n\ui��BX�3�_���X%�L8�8&]����1ۂ'���0��] ���<�8���@Cx#$cr y����$�6��Ml�y�2s�,m�ۼ������t�w�D(��Au\���s��M�'��{��"s_R�ׁ�%L��s��,�Q�Q�V{��{�ߕ8k����e�_����bɬ��[�zO_\��qu��n3\��v��XQ4�ûI��B+��p�?^\����+g����^'M�߬6s?���nc�fOD="�a�t%���ޝ��=�ɌIT!^��U�%A��Mv�z�I�v9@t��Kԏ���`� �:��4T�=���g��zP�|���C�k'G�ڙ#�S��X��]<��;a�p�~�S����g�m4��Ve�.�Lp����=t�!F��1-�˛���a_U�B�_���~�:�P;�e.��5̅V3C	�!���w����g�o0j<�߈��@眻hHِ�-?Z�+v�D�'i5q�5��N@ H9��X@ �Cǂ�r7�w�T&%!�Z��Ja]B��$h���v�9kñe'��-���[!3�y�*r�)��F�R��a�5�.瞻8T��|rmR�V��+���m�ZB�;��-�h���g����A[�v�
�ֹ2� )%� <_fP�w���B�D��Z��M��k%C�O''����I�]Җ�F�6�{��e9
Ԉ?Ak�6�S��G�~���uX��ןl7t'��<�8=j�*z�$��p(�4.ueD����]�g),&�D���Ay�؆\t�e�r7c��}q��'��׃��Q�o��|�d���x����������/��J��(��������n�G_3U@B�a���a/��s)mW�x3�x?T�mV�(��j8;�%��#a�[)@VBS/���Ω�KNE�A.�b_6��pB=F4�D�N|���bcS��-"���I��=Y��n=�׸�u��\o��V:Y|�I��&�a�ET��X�%���E����+���!_x��6	/�P��~����6�@㔄'���)4�RF6㓈���2�|��?��$G���QR��֮�DA(:c�mz��L��N��`���m	7�Tw������(eĀW���"Kѧ{j�T�Y<b�����e�Q݌%~�N�\Y-��G���l�G�u&�rM�Y"w���B1�������D+n�M$�������M��"r�,���7BՃ�H�HTL O����?0����Xx{��P����ZP2rw�/���3�2z�45�c��� c�_��m�q(��K8��/��Y�,���_�+^�6>_�W'��풦&�*i4u�Y�+�b�(��S�2$�Dy�ֳ�:h��2��t/�km~�Z
�J�	��"\��1�?��q���RKW=��3�ck�����]t$S=ob����~��i�,���-V��^��ng#�rF>�X�	tA�:�֝ ��8�q��ϣŬ�����i��C6a:��7G���_��̝�k�&;���xSM��%�D,�෷�:#g�B�Ͱ�#q��f�CW��A"M�TIg��E���	2�zL�O���3s/'�NP����^eӌ�u�zÍ�'a�ە2�.R�!�b�U늚��St�8�}�<@_.�6F���G��Ը_
W,3��tq��qdvC'��q���v�8�]o�C%"[��o�)isW�p$�Z��&��oɟԌ�Ү�j�����������	��H!h�����ԒW\xUh�[���s��K�jT�F�	�ˤ��.}Es�E�'�ہTDB�k�>�Ukg�|��uE���Z�R���n) +�t�m�H��n�P�T��6w#�-*ݩր�,M/�SÓ�� dj�ډh�2*n��W+es��	8m�ק�d.l��SQ7��f�0�ǄH��Ԫ�?��{���t��9ת�pµ/�~�&���X�%Vy��Ӹ�@ ��+5#��B���zx�/� �9fi۾�e�������3�^,4>U�5q��[_�I؊M�w�,?f�VQ� L]�c��a�x��ؕ��}�e�h&�D��E[�z���xg<�K��MM[����V�i��t#��_�障�"XҔDB�Q)4"k�b��WvCϦq�3�nq��3�}9.]��d➥!^�@@��b��w����߂k�3FX�&J�5�w��6���Qæ;3�=�q��_S�3�d[�����6�>�\��o�k,>��f���yT7"f���^�����һ��A��@��ͣPςfG���HP�֛R���L1hV]8�t���'�4s�8yn���&H�����Rt ���l���j*h�N��4�	g�hug$��l�"�_C����q_2=uw��l1	�t�7�Q8�}뿒^��Ci��HD8X�,I��v2���Ã���R���d�)�x@�*%�K�~D�u�� ��Q񑲕� �͖4�Fb�ޭ1Iְ��Q�&��2I�/���?�S�,���A�V����U�)<ć~�Ăb�$Z�/��A�Ӛ#� J����r�ˬ�=V��1�ه6-}[�����C�[wv�y�@��v6�f<�I�����-M�4ke�M�%>�&]xd��xd�Ca����{����5����M�Ir��66΂A�h�����ݿQX�9�	�z�&���c�8��'�т��0��u�Q���������M��f�ԝ$�,�Z���U��� �1X��&6�2r5�m�gW�0���'�E� �s�1�Fb9��Y�~���_��?��]�F(poF����6B�Nـ乁I��n޸S�:~	Z.|�=&�΀�b�Ϗ�йͣ+�=�����������˷#tM7!��F�PE G����0Q���7�ZG����r?��C��q҆�:�dy�c�*��f�pY>}Y��XTn,�=B<�ck��	K��͓I�L�}v ĭ�/�=�B�f�U�,,qZ�|�jL�^6Ү7�a����cFҍV{e���C�>�N@���m{��+��D١�g�e�eL�x��-���)�gh-�;�S]��'}���㭦�����1�{�(���#_�\ZG$Ʉ~�W+(�i���F����a�%_�jx��1`umc�M���Q��K�������c��:�����{o���xJ��V�=�̧+t�5%HOi��X�"���-�~����z֯��:.�CL�H�n�����9�����1(<�5�=&�(�ْep �9M�������zE<��-~�w�l!��-������WO�R�,��~j�����^뺭 `�7=N��ǡ�.�M��t�������#{B��&��L�$:�&iH��/{h����Wx����(Puv��M�/��~��ds���]&�q�?�R� >��_}kk���~��d-�J�OU�&��	���G�>E$�}j�G����yB����7,� �`�����Sb-���{�U�b)�����?	������@���h�ļ.���X��4
��ÿu�֌��	�]��؏��+�&Z+W���j[��}��X��H�]���E#揯�������J#N�o�����T�K���ūs��P��,$�O�������ڑ�����)X�X:����{=^�[y�&��dr�f�tZ��kȪ�d�E��+�B��]_D��CS���w��;�k���~ k���u� &8�EbU�O���cm��N�<���Hy��RAhD�����y�C܈�훝 �+�Pu3�u��{�f?=�~�K��hl3t�H��R�ڟ����@���n�@b��~;���/3�Z�WB��{H?;���������������I(	�L,o7�����
WQ��"���@+ե$q@� ����mY-��o��X�F;�ϵ�Ʋ]a���V���/t�d���� W|C9�1����0��rx`&.� J��A9���!LYI����*�R��q-
��<��t������Vq�d5����_�#
[
�I�J���M{��yf�sV�#�͢�W,R���bK�hE�>c� !�"/$t��؍T �
x"
��s��h����VT@�Z�^K�H��W�=4'����M8	j�"�D��g�q_�!���x��?%0Ǽ��Y�)H�|�{��֙�d:����t�G�y��a�l�(�qDIb��m�9���S��=伺c�ǩ���-:$$�d6�G�3D6���%^�*�h���TY��������o�����:�������` (ҁw3 =֕Ǐ�q�
ads����-z%���R�*_��0Z�:�2`#:t	 ���D��̀1��L`u�*�-�����W�>+����mR�%y'� ��)L�sm�X>qLr	���<����O���T>��0p�M ����dp��+��EV啅ИQ ��'��Qg�18�x�=}-�۝���Q��Ȏ������"�V�C���P� @�Y�g�B��_�廷5�f�<�
�^�����0���ȍU��f����nV��Y��䗐�B��x%��33^U��r����VR\ld����4��ot��s3%ke~�����C����U���<;�Z��SRQ������;��L�Z�D�!��+��Q:+��(@B,+�HM�,_�9���Moڣ�Kܩ�k󬬙ұ�1��XNs���q�>U8�Cd
��YU�.i��
P�2��V�F�97��� �!����6�3�YB���D�~�e�sDgR��ڔ=������H��]+�HT�V��F�L цHլ��3|��f����kF,�2 `B>.�hN�	%݊��n��tK���'&�:'í�c����&��/��#��}�8$D�r�BƲ���V`p[ +RAT��Y^��Krnn(�fN��Acrm�*�()�k �I��ԙ4tP�85��O��O�es�-��E��� f3=�<)���L��8k�O����^<_֋�l14�z�w���@�a��a�'f������|9�U���N��mN�i'} ��33?0x�7�[z��5w*�Ʌg�"I�fi�	��F��E������̩A�TlF��:p��������K��5zs��gC��Ǟ�������w�J��9������?wz�J��X��L�V:�L���L�y�jc��L��~�&]��} �b�p�5����O���5�JY�f���ش�v�o!��e5�0Y�<�0��
���k�F�$�S���� ��-�Na�M��d<L�:;��3"U�~�Ud��P�����(�� ��#���Y�_ilZ�]ɣI:p�rX<r��-����3��ѮȀ�L��=M*��8L�=�|�JnKe����lJhvBo�$x�E��1��[������%�Z(��D����cX���yG�!�Ie毱�0�����<��\�-���a�K���en�W^��\ۏ�"��[�i�Ea�7��fvM �E�-�K����& �Oq�b\��M�.ͫ�۞�L ��5�ѐ)��J-�G$��2�B��b��ƣ1q������R�����fâ���]@��� ��0V�T�io��G��mH&��$R�;��H$���5A�D��A�/�_���~>S��e��m�~��vý���otj�;�]R~�f9���s2��f����mu\Qi�銓��;v�3*%t"9qy�����g��2�#�7\�3H<ڻ�{8Z#n`(_�������8�=Z�+nh+=�����^m��;�ݗ�V�)���-l�E\��'b�O����
��k���Xʿ|ac0�1�����%{Y�⏫�4)���a#��:B�*�~r�C4+In�(��'�b��~.����Y��5����>���
�*�B�'�2�;W~�:��Z؟�D����[y�G��P-��ٞ;gq�(��E+ح��ى�p���Q~?`mf��#ҙ�O���2o�]:#
��H��c�@�a#]������J2��iR �7��c��fe寔��%$=�xa4�t��]Q����R=�J��y�?,S�޴*%�`#*:����jGM��H�/q�:-*�y��9`-���]�yV���x�t��Q�EZ�4�������R��:�jj_���&���`��[�"�@�5!�$k�W5»���)���_��Ôc�9-��-�dS��!���W�Qd��I����D�D�:��y�W�m�s���H4�,A��d� ��'�����Ɏ{��0No�����֐[�JKJ��b�Qj�)�P��WQ�}r�40��q"9�bH�:�)PL������ۓ[���{�����5�Pu�hW�] �N�\�:�P�M����HJ�=�����1nA
*�)��}��͸v�INJ�WB�4���C;iN��PI�Q-���_��bD�Vwΰ��~�j$g��^gx0%%�\�EciP�>s��r��c�;Hǉ C�0`�5ƟEZg��\�_���#��'�h��F���;���l�����s$���!�?��JV�3�-ּp$"���+��J=�#����z�Bm�lw���d5�eW�!WN� ��IP1���:e|����v�1��{u�V-���	�)�<4#�Οa�q4����n��w�/C�@&��lH���߄���!M9'>q�7(���\���Y��'M�;n|�LA����G�^�^�;��2���xb�
d*�5!�V��gו�$qB>{�w-.�pA�
��
�)��V�[W�k��f5L�P�<�
�W؆�~ė>����%��@�%�:H���'�T�I�W�g�A�}�ެAC�K��]��5��ߧT��6�Q���Uh����{G�A����S��=ʻ�߯��#V8T��J^qƢ�_8��0����pg�i�\\tǿM��D�z}�l��t�G�>��uL1��;�M� �$�Xπ7D� ��2�h��UtS����I.L����Ἑ�n��@��0\�ҏ���Ю ơ@�ԭ+N�Zk����~���`J�8Gj�s�Q���e��ץܷ?%o�ql���
ܬcu��}�e4P]�\�U�f��]�fD�d���[����_X��Q����z�0������O-���^�x��4n�U�܋���V ��\�do/3X?&�P��L�k�M}����u@�:0��Wg�g�C�Aw��ϊ�a�T0#��=����	�a�&��ZiWb�.E�q�#\BN/O�
��JUL�i��XԞy^Hf7,v�AXк�l7� �)����
��דa��'/ �e3�Qw���c��s��3�#ũ�a6�@e���
{qH
����EpZ�tx��N�Y�I��}���y�+R�ޡ=��}�g���RYQ�y�
t�z�d_*��Z���`Z�nL���H�)|���5:�wd��)��u��w��A4��A�>�U�$�;���k��!�(Hs	`#Ԣ$@��Ry��`#�P�[)��|-����.2J���Aȧ`��I	oݱ�&R��v'�Wz�?g���=�a;M�=<�Z���1#_߇�)�$-�ެ�~��\���f��*�6���>>O����vs���J����0����:����6l��"Y�<�e �zI�=�E�o��|�t��q[�o�H�%�D��t��b��S�fXqn�F��T*
� �9�����1M�0p��PY�.���"���p�ﳸ��CUX ��..�7=Q�9C���U�~�
���|�70vW�?Q�5�3+�i�"�7��]�����J���G�5G�Y�I�B�m�
:� �Ћ��'4k����{����-3mVW۲�@pbT��	I��p�~ʑ\!���0���J��C�h���7	m�=����n��vK���7d��M�A�W���/�F�p$��	Y��/p����M��\Y7�4!@����\�ď@ֈ&��r�x�Y��W�'B�B���R݃��ϛ$~WXw{�1��e>_`��6�)ԭ���(A��s!t�x�q��V��E��R�/d��s��*KE-S��)d�O�ft>Slٺ*2��N����8�z�5K���uXHl_��B��ԯEo�WS�QB(���d�8�j�w�lц�%�Yf��#&�TU������z&���z�"��x���HC�ʳe����4�U�d�w]aT�gfyMM=)煕�����qS�SYk�s��	�ׅ���٨��0�e4�T4��� {�Fb��*s.�U،����0�L��9��,9{*ҋ��!a8Rɢ�s��$��H�9~;޿�	/�(�.���NĦ���o�Qef_������CM$d��uPka����S#��L�UN<�B���?UK����>ѭ`JKH�8t0�ba��Q�<q�b�{`�6H�eI�+[b�끨:�z��y���W\ͼ/`>ڥfP$�g�_�R�Q�*�@õ���R���ˏ��x����`�r�E�5V,�k�'c?4F �d���BWK�'$�,�-���df;�;����w��6���-���b]�w���?)ˠ�Bj:}i�D������1��P��'<,��f��K�;�������}n���¾v��ԦnSE���6'�HK�����*YݠG 9%�00k��ś�L'}qr,En�o}}�S4���k �2J�̒��{C��K!U��
�LP,8䷀e���Wf�H�M�I�Q���W�i/Cޙbѡ� 1Q,.�g�~����:�N��>��#N>��^�E;=��JX� u3-������"}�`�Ԅ���M��ސ%����ыw��WpA��C'vf�6ր.7��	��(�k�^U��<��i�ʕ�H�g�DMHQ��Z�%	�h>k���m���������RדX��k�Pa�钎z)7�<+�\�o��w�ӹ�`�h)�>B*b��k�����Ю�%ߝ\H�fZ�Y�����~S_Y}+zq��&i�&�ZMU 3K��ȽMZ��۩�a�H�(q�뗰�{�9\��{�u�w�J��{�$i�ȷ���&�Q�� �E=��@����0	e��~in$D����go!��.��N�E�.�Pd�kSK��e:h(�k^U�т�p�C,��������3k�?t�ȫKU&��A�d�@t�>�NJ����u�>0Z�Ng��ga�^VP_���eT]�>e��-)䢊���SM��)i��)��>*S5~�]�O]��Q\;��EZ��j��}��ҋtӃU���W^܂�d�C�3¡�Y���8���VRa�E���Q�r2�A��P���w^����8Dx�~���P^�H{�V�E��䔴?'�
<�O�8��<��ps�|ìqwg%�����]n
1yo���� ����p$���^ D'�ASp��|s1�Ǡ�Ds���M	�p����oں8ױ�� "��l�-Tܢ��X�Is7-���
�Ӄwv�y�gޗ0y7X�o��E0gp3~*#������.��P�[yj ��l�����F����T��5r�Cًu�e����
aGt�tX�XP��N�m�2�|�»��V��6�g �Nh5��襹�B���]���Rpθ@��KhIR6�|�� l�����iaL��7�)�>�˷#\+��
�����&����B���DU�|i�=���~�n��lDr�ժ���Y#�jW`KH�ש���*�/nCH8���-�g=�#$���&T�=��^8�O��䞌�%R���_)W�}��at��}�k���z��7�`p�t�}�&���ln�A��}�q�-�L����X�d�2����9��}L��~�%���@��HD���j8��fD��M��=��Ԅe��c��vUz�VE�e�Sd��|k=��E�ף�g�*Z��d҂a�oC���qY��4�g���Pn����x٧��5�̵�Ā&��a;\o������E� +��@�G�@h]8N�nŤk���f�wOa�����Yd)�b T�+��9p�K74�g���Q����Ӳ�^�1�`)2Rr�1ϱ��� ���^j� u�dP������G@�F�F@Mt��LRf���>9���^�	?��Q ��z^4_��l�}��b�p�V��y[j��q��[�����������k�����Ϟ��Ҏ)h�g���, .�R��r�/�Siĳ�A�-��k�H3���ŭcZ��\W��V������.���\n�[U��I	>iR��V���!C"\�}!<]��ĩ,���-G�uV�$5�;y����gD#�,�mi�/#V����%=��[gJ��]O�f�$�`�~[o���U1���Z��M�ȃo�z�dm�����	����`����%�I
�L�*���=�T>��I���;�o)/���|�ܱ�)�2�nd�ݝ���X�K�~c�vg|(�::'_���`Wjǒ˪ �B�ii�Ե�tN��	g������N��Yn��?����m(J�Y{�b��Y�Ώ�P�$��ĉ����ᛪ��z��sMd�ީP�9���\T{%���G�"���,|3��/{80�D�Εkk���` /�"]��_�uP;�Y3kb�W5�Qn�J��F�*q�������w�L-t�������E�dZ�:-����T�\�Gȃ�LSG��L��HL�ۍ$�	#4Dع��1�*�<��A���;Ƕ�q)�o���oMG }VA!��rN�p��?�<���%�_Q�B1�X�E����s�y��%�ާ��N��v�E�ٰ�D{ �sMJ��OO�0��_���ŵu����Q�����Mr��2�h-���銃�57�r��Z��o�޾ ����i_���42.�Hr#C�d�j~2�v�y�x�e��������4��a��@�
7�`�V��5�D�^�#SQ2>c��x�,��7�ύ�ꮩ��ˋ�/��(�BX^�B_����x6]����8[_�ˊe��U�f~��$���� �e�FVQqvn�1W]�.�B�۵���ZoO����Ɠy�\�Ŀ�<d
�b%�^� "��f���nA�w�������(8 M�fJA�$��A7�a�]  �}C<T��[��đE���a!_����U�,����B-���(��2s��_�=�%�B����S��5�ɻ�v�PCw�_�=g� �ʛB�k�!iG���l�ơ໗c0S;z�r��sp~Rڤ�b�H��*��xU_GP%����6Wp]�����^�*�!a{Ӛ_[�Gb�}�t�����v�#4S���Y��������Z�?�B� �W]ݪ`�v���Q�̀.�a1�OG�y��P�֝.� ��6��ki�k�C��ٳ�
�f->�ke�0�Z�-:�^�p0�8�o#��c�1�ʉn�ҺI�n4�'���G����4���#KK���xr�"QW����m��&��	��l#��M���<�Y�uA���K�7�%��Z�Y`�
a�MśNO<����D�R��M�Z��퇂o��+��Q��d�1t��&̀�"lNM?�]kZ(fp�����g��+����F_MV��q�X��֕��Xs��;�ED�Z�VۨE�[��?1�]>e��~�5:?�ULiX�>f>%n)�����yr�5����w����>���U��:���a��]޵�	�R[�VBE_��m�i�Rs~U��Қ���!�EbM��DyQ|.�͌I\�ޝ|9������I��n��y@I�����Yew�%�1D���aG3����Vi)ܚ����`M&��}�7fщ'�Z4�0<��Ӯ=�	lC[�y#�9��e�.��ړ�P��(j�a�/��V�X3���`K!����>���>��jTNr8Tܘ/R�mS�Y�t����y8��zI�XZ��!��j������;�S�E�
D�~Qj�GȲ�i���[�J|���B���	�Ϩ]���U(%'۩V�F]��\��cU����iq~&�U 7�Qe1ё����X?x���nɺ�1D� E ���i����
w���+�;"�1�&���H"tL���/�A1-��֞����.C�y}���-��j|*Xz�c���XP�%�4	u�7��<������T&,\#�].l�a��#	�mDfn�ra�4Gb`p�'����<�M�ȓ�H��t�����*=徢�P_�P��Fn^Y~R>���Ӳ�{����W��L4�ķWLЩ��/���E�z���B6�6]R��&�~��s7�a�& �i��-�l�v��!��
R������y�N�p���r1�M��B{/��X�)����Rǖ��J�'
*�:d�M����睋w^S*k6z&�e{��*]�ih�@>���Vsз��;Ǒ�����&��m	[�1��ʃ�3~����ך�f�5�����z��}����2(Z��X�%.jI���YaB�rl�e�M�E����9A�/~ҫ=t�wāz�c_g�mP|�����Mih���߃,�ôXHՕK?F��U@2����c�{���@q]�U�1s��ׅ!�9��i#z{�.wG�'�TVQyiB�iI�(��c-����A�^|��^�o������%�7r+$^r"����9wR�:�r�o�����Vvw���*�X�M~Q������"�R�,ٮnF��	a�W���Η�B+C�h
���-s�oo*�Wߘ?�uStg�_�������,���-�B�<I�+J��"���,��I������+��mh�w��l]��w@�V��MuHWB���̂��*1�6w��"��pKj�{݊,Cyh<ZAh���J�+o;��Ӎ��?bSG��cY��ko��OV<Mc��<��x��i�V:s:�ݷcuLQA��;K�AB�<R'��]0!mH>�d�G#�f>t5	��k�"9��ُ��L*�}Q2^y���7��\�/�l��S[h��r���aE�ݟ
�L��J���\���'����X����O��j�nM�}w�ޤ�`|woF�&^g�cl2�[�]!�k0�ղ�����la�\x��$���f�2(�ƶc<�ET���Q��
܏�Cn��Wui>Z��&��W:6z��3��Ru�y�@|v��+gZ+�Z���$���]y��x��Y��N4�D�B͂�q��@W���f1��]�/���N�t��ӈc��,z�1��;��>����,�׼tV-n1���}�WUAF�@�|c��[�0в`؟��|�U����x�D�U6,!���iסn�| n�d��S��䆐��y	g<h=�'�\�?D��>�(�0>�[�R�D�+l҃ؓc�OD`k��DcS8J*��7E7���+7��'k��)�&3s�k{�������f} W&v��\�.�;�P�j���.ͥn��բ֮�S��J7���M>a� �b����+E0��f�H��%�$6��V�:����1P�|���}N�p���,�pW��k��>������hCލ��@qQL�_45�#3��z�*�K����`hJ�i����3����*�|2'��
���scBL+m5�ҌlH�Z��yGĘ|�k�ˬD���8�$����H�/�؉M�j1t>t�ڿw���p�D��DH�O7��IH)���D.X{Pc�����'�?	�3�u���zL΀��?;�1�+0�����)��E�8����$%??�b�5��)�8˕�z�h5د@���*m>t<�l��>p�s掃��7��MzȀ"�\R�"'���A�i�E-�X������l��z����f��b��.ΪS�8@l�Adw~E�:�5��
���ƞ�j��DX���*��.{�wVcY���Ǐn,8�l>J9Pr3�brI.��"�`��/�ΰ�c{�/�/VQ�K�& �s#l.��w�8:�8�4ş�J��z�B�Z"��b�"��b�pI�j��s'�5���/%�,��|69碠I���8���zZ�G�Z�o�M"����?�}��JT-�d@cEd�[�Y�(a�
!NSU�iѧn;�w�#B.�RWex:��f�a�y�� S\_������
KU��>�����@�\��s� �َeSd!Qh7�F�dU'���W�>7�\��P���5���ڻ=�mR�-�۴�"��BJ���4�p#{��8I�h���(���r�P;Ӧ�>C��r��uAj�	�<���6�?@����	��t5�kc�ƹ�,z'�:�?�$I��K_x�Z\�bl(�bzd��e�7��RvA���l7"Q- '-�._Ӵ�Y/��o*��Q����.��9]��a.���8����OB,s_b~��򊢷�f�P�)]̞Ll\+3���NUjJ�B�s����맵�~��XI<�g�S�S.�/-45�>�
q��Ӳ��?)Ŕ�Ѝ����?�۵������9�*G��rqaW���~NeC�)ے�&Uv�@R���4�����O�����|���c����r
�lL:���j�/e�p�{%�J������� e	�4GU�&��ĭ��.}ʹ�V<WH�J�ʎ3��p%�c!m��&�����AP�_Cmi�L
���z���a�/_:�Dl-�t,�	T����>�Ȟ!���:�>�빼r'<�f�uT=��D�����M�S��A0�t�j�l���P##��6���p���0�uì�DH���\�[����Όr��ƻ�� �gh��N4+�]�}���ы[uieA}��)�b�\4J���4�b�����\D�Q:h`o��_<�+�:�,�!׆@Q+�G?�l�-�<��ד��M�Os�}?\P�nń�Z���I�i�FKx�O&_f�
Yݍ��2n�Q\���ߤϦJ��5,�v�u6�|�F�s䃊�z�^^{So��$pJ�ی���/��.TB��&��9G��,_��RӀ,s�b��DX�UPX6�|�s��<O�1?�h����l�)Ȟ��
���z�2���󣁴@�
9�?�{�y�/{Syт��~��Q�(dZ_�C�v��O���Z�.̧N���������B�U���(ц��O:�9잿�Zɿ�:#g����mʽ�+u�d4���Ř:7��W�>G{`���C$t�̿�B�z��尔�D��N��|%%�k�I����Fv@��r^���

�v�7�RJ�QR	~����G%��O���e�'�`ǔ
*��P>��'0璳�O���,�N};
�h*Ȇ��x�c-���\�A������W�Ԕ�;GB��/�F�]������ �^�������}֓�DJ�#�)�Ug��}���z��� �
.h��p� j��T
�pd7hWM�YT��s�h,���):��-}Q����f&C�p׆hO97�y�n��bz~�7��J�W��j��C���3d���5���N��Y��y��b�{�Z|� W��^��tגNg�n�Qe�?�����f�aX��|�z�G�^B��:��Щ>|����R�iUyp�ayz���S?	����U`�ևC
�a�Ư¸�F喕N�M�M����g6|����9�zR��j]�1��M29Q�n�A��Z�K�L*�P����@_p�uЭv��V��Vc�s{�~��:W����O�@LN�6��P�Ȝ�B��Z��Ԛn8y��$8��E���<��6Z�QN8w &2��}�Cb�q?P#�Ќ��-"�d��
z]7��%I�$r�#ibm+ꜵ9If�"�@L���I�6���^`0�����y�vfa���j�!�L|�$ڂ�K�De?��K�Gs���ද����;�������')QC�j�-	P�i٪$�]�.@q庿�^���J$9s$M<�FЙ�h��WmRu�1�R�kgE`N�n/+�`VP,M�IC\�L�"qwQ�)?�?�ǓE9D:4Y����L/�!��y	��L��/>�=���+���mm�|���s��t�Ƥ`���b���B.��"&)��� 5�zW�8�s���F)����.��Ƃ��U�f�
�h�2V�����9؇�PᐉUO�7�Րs���s�=�rP\�Ks��b����V��2��c�!�Ժ�9?m~bq�g�:�~�*���;O)-w>����nQ� R�VƟ���!.�p�T��Ɗ��+�Lv��-���!X���g�A���L�3��p�=���8�jFGm�6ei�	��66�%�p�2�&H��V�G_�����������a5 ek��|���eq۳��`-琣���p^��-�b�c���?��R�h`M�Ç^�M�X�݌����X]M�y��|�m�_�NN��� e�8�V=H0s��:y2<{�CsE1������f�j3�
��H�έ�]?���O�=i�����g�.���80����I��ѱ���	�L�	*�P�Ϡ��=v�n2O�Oߎ�nW��]]'�|�����;PK~
����W�"�%�R��(6�MY��*`X&���u��$���Xs��%�\ϨӚ1$���@72U�����IQ�������~[n7�|B�i�ut{�����S��e���.F�H��1z|�R�P�*롫�;CE��߀�8	��T�����vB�N�5�"��q�D�"�ֻ6����NoH��;�2��?iT�u.��M��-��j	���r�'�J�÷<��S��G.�����|���ʨ^m��~�NG!t�sb�M���r�-9��r�/wY����hU�?��/��x����B�!��m���_jl�؍kT��4�+!�9ғ5�{mؚG��*Ryڱ�������O�#{���1��;�'�@&יϓ��I��Ty�:�o���+N���hD��#���_
�Ztk7I��)	�������jQG�5�����7C �茚�GI�!"@���e�bX2;��L!_��x�����*�GfPz'ލ	E��j(��j-���ihL�(���;��B���I���s��p����csCb�5le䨽�vmA���u������T��2Oȯ ^|��ςC�/�IE�p9R��TU��U5���]�b~>SI��y_u�nq�~���|7��xy��D������nBHװf����a"&�]8{��r$fV~�c�����UX=>�� x��'���8��ԙ�V���a�6v;&�l�Q7��z�z"+h��*��6j��/C�3O� ����p�I�
��7� ��/����'�O(��T���0N�y��F@|��O�Q�ˑLAy�w	'�d4��7n��P��� ��� �|y�!��#M���9a����Y��+�2:<9(6
�O�>w�cZ�׋j���g�(ӥA�.�W�a$U�<��p@j���+�������9��	�~Hه$Y�.S��m	:��b�4�*�]�~Xy���²������&��G����9�1�MRVǚd9�J�.ش�O���Y3
1��h��u���8*޹�C�ʛ��ei��*�_p�֍\1��ukm�D�������tj�9�d�:ɾ���i��<�3.�n�
FeȚ���&w���
'�f�zN��l:j�^�@GF��Y�G	�8	�2Q��1SA����e��7�mv���U;�T��<�����^sE��i+a�B��L���B�-��Ȏ���<|
jCh����B��Ի��r���'(��)R��:�젆^��B|����G;�x�.T��ߩ]��Ō��̵[+*ت�[�Je��,`��W7�x����]s�nE�b0�ŕ�����M��i���D���{;t0�흑N�0�AL��M�7-�����5I;	.�G|�G��Vd!�ȒKg�U5Ղ�����]g1�G��Ƥ���d:^&e������eoO��.S�f?����5
���RdQ�� ���З���Z����}�^�U#�W���&�$8(P���d�u����m��Y�g.�~,AS_O��B��{�n��'%����mtH�O�����M̈��,�<��N�J���@A�yĲzK[�� 	4�ج���!VK�6飑��k����w�iȠ�'Hv�/<:�r���mgW��A#��Z6/�P����|�9��ϝ]��EM�u�ݕ��n�j"2jfְ����ȱ��:���n��o�/ e����c���ѕliWU�_p��TD>�ql� *t�a��-9l(�,kC#����Cn�Y����*���a���ƾq�S,��N���̋�7):JM��G�cn�\�Z����\�߻�8���#�.�O��_o�+�����S�Ao�A����h��{s��I4)V��N�e}��G���j�Z�1Y@ٍ�\�1����M���#~�˙�y�2�Q؋f4B<�}����̢��n��i�Gň�?8Q�^S:�=T�U[��ܕ��!�3��M.SQ�8���p�Y�Q�Ki�~P�(�b�v�<F�:�/?��� �v)-z~[�K�L�<�2})����H�-��{%{I�1�!l���816q� <�H��M�6�@�!�-��Y
�c|{Lc] �����6�t�,�8`,���α�h�8ǹ��A�yD���xrIp��՚���9F�p�~����@"���zrٺq&�Du�|�����\��4u�cI�m�"2y�˲s"�<����`�*Ӄ� U��N����~jD�|V����̈}&ӭ��l�I��7䆺��@��Y�q���'z���0�U���!
Z��
�/L*u���:'��8�w٩B��LJ/Ã{��&�H	�=,�7+���4su#�<���@���Mu#U��+>�@��)as����q����ܣEni�;f����&d����HA�(��I�
�h��ҭ��x���V/Э,��(�L���{ug：F������V�?c�zd�jx�ޓpz�����`㗛/�H�#㕩G���d��.��N$��to50M��g~��ʝ�K��"�KwĊ��Z�u*mY[=����Zڧ۸���"A���MC�t��k8�`�C��-���q4���U���Z��������Ҝ�K
{�){0��L�e��-Ú��d�����" S���M�ػYlr�m�s��V�᫷|�l�W׸��q@0����W�P�5�T��fOf����Hǧn��,79G�������RȽ����co{)��=�mT0e$^����6e�4M���� j��BJ{8�u}��!��j~�zH��.�~n��&�{�xv��Sڂ*O�>�}b>ĵ)�|:�@�y�k�o�{lS!��PށJ�Υenx��Xu���^�=�z�����J%�����ni�[��C	���Z��Ģ���SI�2뽩��-Fs�J�*%���t!��{�����4�#7��/��Ar(��WW2�p����ʿ���!�n=oc�:�yH 	��Vʻ.�Hy>Jt�"���l ��Ȭ��ʇ�O/��m�.�֛݄�kJ��u`��G��<�h�k!����4�1��� �0ܦ�ҍO�Pa��������ZŔ���m�j���o�1��q*������3PX�h?�O�u��C�r�]�	���
}aD�S�&�/;ְ�|��JI�QrH&�pOeV��vwL������[��*��O�1�3\�8p9�O�'9�}�!��f+H�k%���*�r�>92�ɁН*1�D�����1R+��rX�-�6i��C���>�ؾ#'o�oʯNӸ����*�K��o�]����U`��d$��:�Ȯ��=���͆<dX��e�����֑@�~�茇�6׾�\��?�5S�t��l�OTnd)�-�bz00Q�q���5�A��3���d8V�������Ē���!g�,M$2������������hϗ�$Կ1�-J�T����Ը�i
�����a@�?�૵Z<���_�D���3�X;UIw�fb�4��m�'8]�#��<��²,�؍�~�qr��Đ(΀��ޱw`��/��m�.Ӧ��Qྯ��ln�V�p�[���ԩ�x2���ru{�"W��4[�Ʈ�^v5�������ǳ��������0:!J�Z]���͗
RpI�#������G�}����U��j	��^�Z$�)��r�-��n��w@���<|�LR>�
����Jj]��L�ۋ��tV]/rّ�{'�-ߛU�so
c����ޜ�2���Us�����JMbf�R"��n�w�i2r�X|XAqY|d�/��� �6S�r-giC�ֳpuQ}�-�d%*�x=/^�Ƈ��1�O����^�c�<���9w;��"�'R^+\YbKN*8Bڈ!����˱�ΞsB�����W��.��5o���3r�?�X��*?��lɬ����?��5K��.�ap)=OB�lZ���M^ֳ�V��\��}v}"��<	'�R#�c]ت�X=W���\]� ʨm�v~G.�KyZ)�K18���)�����=���^Z'�GMĸ	�wI39��`��ߴ���f�ϴ� .3uh_vb��!6�g����&6�b�� ��yVQe�z�{6;T����DN��6�/����� X����5�A�`yMieO�(%z&́����q��XL���i��ݝ$�Ͱ�!"��T��{�R,0f�7�aG�Tw$���w�r�垣Mwܒj���}f��&�M\�L��'���8q�`��~+~Q5"��r��p�z���{�9,������tyf�L��D�p�G�q�u ����� Q�����Up�C�.?�N>��@f�ʷ�F5U��a���=���&6�.��5�$����GO�n4�ម�9N9=_�>��N��z���;�b�KH��Rb7l�.��������q�v�eJf�Z������<ũ٤��b�*l����#^'�P飨��O�p+�?a�v���u=z�C�7�a �d6τ�(	w�r?
tK�mB�y��h.�������Wb��E����Q�������u��iG
�xvGJ�<�Tߤ��$�&��ǁ!arLFm �d/��i������p!��h���KWf�z��XJ�'�`h�	Q$�^$�5q��J��s�-����9�,L�×�o�"U������Q�B��W��_{ƭ���h�G�8&('<b*�'���=�]��Rn��M��t��E�_���R�*�>#�xǪ�r#сM�,�f#�-�@��*�%��h���h�c�� ��in3�k����W=���Wӓ�\���C&�w�V��L�vc<��*��H��SB&�`<_c�����hؐS'�_�G����>uC�%[[��}ر'�籆q]��`��{l|��_��EA�����4��i��\�9"F_OB�'W�'��&�A������?N`�.��` ����xK�zG��@O�w�,G议��Y�J�k_ʃ����dlr}g�фl_�	�2v�a��W�2��Q�	�J�,�L��f��<r#D����g��Mem�F+R�?9�dO�#玒H�s��o��xW���r�nE�|
*���TK	���s����� `������V�yړ�	\���~}�G�J�U���GG}G��k��?Ⱦ.��E r�?v��s��HQ������O@�~�'8Xf�-�ڂ�"�A��Isq�[yS�?Q�C)���`����R?�R0G� Ҡ�
�A"��1��V�`���gU8����[�`��v��BeZ�:�#�:�(�?���M`��QOĎ	�������Y�ҸI���[��?b�^��޹/?a�>��G���;z)�Ti�Ӎ��}Q��&�R��E9�M
��)b�;����D1�%�w���r�&�4�c�y|�Q�T��
+�"ښ��;g0�\�����vsǹ/��f/�L͆�v�V�>�q���G�0CGx��1-��Lb� N]��_�C�^���ʱP���3wF������WO#�b�,���WE2�)�B9eF��ڽ��,v�Ӗ�vا�&#C,�]ѿ6'��^�_�DFx~��-?S�Z��a.��X���?~��m��;(��|��J!V��ϧF�xݝaH��5�%+�����3R%1��tJ�.n:�1�,�#���PZN(_!M��K��aEh-%��^����-ǉ9�L� 8�b�c����d�|x4=��y���HV3/Y�u.4���CӺR�����e���SSy�*p�g�>�L_l�UR���PhʌK7�KӔ,ϩ_��1�h
�{pY��U�"�Y�\m6{���6�����j"����|C�G��TUDa�y������<5���
��[9���!��Is��R[B�VC��p�#A�%"��)GrDċ.6�**�7���$�d~	����@LP�����fi�YodD�H�B�2	�d�(!1��z�>za���K7��	�0nk�{�&�M��N���+#Dy�۲Y���d��>���=l�s�����4MK�B"'S���G�ҳ`�d��k���س�r�d�ず�����1'���l��̧袉1�`"sU�ɘ�I�$N��on����y�JS诪���f�?���n��oa��	R�O0��E��c��
*�F��hL{C�n8겳2��Sb]���e9�B�b���h�m=��0���HJ�a�cdj�鴆�FA��5tJP�8k)���`�N4}�yf0�*Iy����O�nke��Y6�z��"G6-�Uk4+��:%zdшI-Nz~�[���_�w�1��I����_z:�;�W���Ò��x�
5�W��D�f���{�{?
2�W�5������]��R�?�\�ud�r�^�)��$������c�?�S?��c�α�,Hh��bW�{BI�mQ R	up�	�c�#��B�O�FH�{��-VF6/*bgz1��ECϘ�s�^�Km�de�����9�/ lO"��cJ-K���P;)7��!�O*��P+\0~��]��������bA�7��Ȣ�{��7�^��Ә�މ�3�2�1zs���r�4R�_���@"�C�����D�pq��t^�WK({�`�YEj�ژ�9¥�Cz2t��)�����7��l�c���N+C��1�ʗ �`�B��(Ա���2�A�����F]k��ʾ���Lv�įv��t�B�0����dT�_)<Ё�����#��ɺ`����r�Ɵ?i���_0 {�@Z9h��榋�(y�u����TY���<��}��(��J[p)Б�
k{i�r�wS@_�q|Z�h9i�K^g"�H��j6|�3x�N{D Bz5^�&�w���Z(<���[��x��֯�,`�t��5�m_/�I�������RR�!�>d@�{K�R��gI�Ij�7L�J2[�8B��JW��{P<�r?��b�=J/�T���h�/Y
*N�1L�`IAB�:�e��M��(�N�J�ı�]E�R�CbEy���ιo؎�6~9���?9)�9� �)�)��j�����p�<N0=sUg{F��4z֥��k��{N8����K3u���0����ׄF"ND����%j�����@��.�����ų��ui�mBZo��cT���t�&�4[��ǲ�uک--�E_-�G�:N��?���0�t�.ck3�.l���-5�Yw	0���zX����pK<E�� S)��C���0_��i�v�\5��zq�������y[�`"��מ�R��H�BFYKW������9 �/ϴ�@��1���'�9��1b\���i>J�S 
��� �ðhF��eN���;��g��e�z��M%6�+���~� ����?�	���Sfj�,��:d�~,�K�Ҧ�m����i��tEv��Y��P�I������NrM�������5݋�AwΰE�pܣ��HH��m�5�L,lj,ؒu�?ڂ;7I6w��0�V��Q�|��i��e}����TE3�Sg�l<��=VԛR쏍�a~��^8<��������_�|���{a���J��Ԙ�qq�дu`��ww��mɢp#b�Vh��, [��Ł�r-+�O�&������{�=�˘19�? �#Ze�3����}\�V��AX�=�9�8�����[3.��,⍥È��a��Xf��i�[���C���EL��T{,��Bf�-\���9Q,����(�.0yp;���\k~b�Q5����w���`U��������f��Lm�"ڜG��Y[����������wX���NzC�L��O\M�e�>E��-��(���.(��E�J������Dje�u�$I������>qV�p/(�Tf��>�G_��/ׯ=*P8����)�J	]�L9�Ú!+ 5ꭔ�HO�_hHx�K�	��DK�����v����݃�=|���M �.V�����j1Y4�3��R�p��{���������$P��"VEBuz�a�{F
FD;H��Ϗ��f�����؛)�ty��>Y�R��\�f�#�L���l��ꂵ�4��)���>(�A,����Ɨ��gъ�nK͊n�:�?��d�'�^�Z�@A�s
��Y�8>-J�G�0�:M[MbID�v�����߭�kW����B���f� ���o�z��v��D�m��߫��Ϳ�T8[s�D|�_Fl�.�B^*�[�N���t�r����\��S`��c�箻�`�m�H^�����Ɯ�˥���y�n��_����Kl�p��m#�o�;��>4%�VEZ]����KPCCr`�_OY��!c���'|��zK�
YC]�i18
l��h�9��0 D�K��cP��u�$����v�L���u-�ȷ�Dȏ��E�i��P��*�̙������1@�cYL��|#OB!d�ϵ��z�}JƘ���̀�lS�4e�t��m��enF����C�D���J�SM-�g��BG��Vϑ�RK6�ρ4�b^S�F��_Bf����\����&����2Yӭ��X��g�v���R2(�_e8���ءd�eP� ���_b�;����ֿ/�a�Я��a�F�}*e/�[���}�.��f�<��!������b����?l&������)HҔ#��e���\�H�1-�v�)��W�@*j$���+�Z	���n��ג���PÞD�\����E��*�qxɀ���No��I)���/�����K��b�>R��G�?�5~���NP����g�C\�W������ǰ����^KWè'��bNC!a���@�`��Gݳ��M���e�,2E���e�����}�k�nM�eGC�\ֹ��/|�@���A<�m�L�a��-�L��֗X�N
�P|@+mXֵC��"�i�y��8t))�9�9-�:��cܙ��_���c��lG@	�w��!h�6,Y�(��Xf�D�I]B
%�A�!�42���q%���^�[P��Jm�!�'�ٹ���9XC[��^wWm��QS �Q�����4EgF_E��6��:����>�UP��g�s��>A���r݇M��A5�5X�x��Ԧ��KX��J�[���U��%oå7J(�Q��U�ϾU�	��ϙ3���g 9�]�*8q ���.G�W
TJN.����I�kh��*s�8�]id��Vd�K~�>���Dy�h�"^�A������'$�Ł�.�ŅG�t�RQƁ�54�w$��]��߼��4�t�p�M��$r���:�f����'�U�֥>����/R��#������y&qb�߈�.��E�l�z���a�Uf@�s>��R��Cs����y^H�Ⱦ��NED�sp�)[�q�B�צ��$��,ف�zA3�%�f���F85�c�;���y(���~,�8��"���##�,XqY�>��[���ɨ�: ?oٱ�����V��t����ґ�7���ռ�*!wɇ�3��<J�:$�ɡl %ߢ,���ڰJt��+����uf�\��O�o����O����Q�|���!�P{�M�`.D�9C[)��DV��P*+ͅ�����V�_�[F.Z����4U�g���A�"�/���ȁu�Cl���Q�Scm@}��3���(`�FZ�
�Fi���x����. ���9s&�F~��uP9?{�=Ǆ�+#8����xD2���x`��r�c�J��U��'�z���Wb��..���x����T���d�/��z8M��B��U_��ťWѕ�����B�P��b' �r�D^�mV�u9��z>c�l})ɟ-��C1��8B���a������ˀ�7�N!J�O���3o�#��.��o��Pc�������2S&n��SK9N����A%ヹ��z��L2��+�}x�$��ɻ�P��t`��dрﳢU�v��(�����~P�h5���Mj�#N��Q��?����G$&� ��� ��������ڌ�wvM�SD�K �|��=oX�
~J���-.�OL�g��w�?�[@�W�0���Jȁ���%y���q;�A6	.�ɕ\�#�ZE (U�`n|L,f������z���;��@k��D�.�G�� �J���A� m��˨��W|��2�^կ�@jO@��giELZ-��Z���5Eho]�����&q�Wà�� N�6��5S�Ē\H6���^�ϟ@�xU��$[VC.�
fS��(�����=�i�@�n6V\ΐؾ�|o&k�(����?nV�{3T��Nl/jXdw��'D&��"#�í&�8��x�!��>�֗�/iyIgBQ[ɨ`�]�	s:Ɂ�|x˖_���!�Ra'�j�.����v�����)�
�����U|�6DX�K�
��u��BV�(2�LEl;�򕡉(BC��=�-��������.f74���+���(�'iwo��L@��ԣ��y�c�\�g{W�".�u�SB�oA'k��PMk�YPs]jy��y�@9.�۬��!� r^������\�e٤K�vB���fA6	�w�:�Y^�� W.k�n8�H�oz[�ōʗa(�'\qO��נ��$��׎jM�)���%�2�2����L��;R�*ϱyn�e4��\�q�e�q�u[jp�ʩ�z���ԽF�J��N���5����͎����1��-W	4�F&p,WA�����*J�M�e��� ��U���Ab�O1�n[�E�8�x��A�5~��s%*��T�2R��®	3�K�t�O�q�qiu$�;��kd���n�a�N}�h(�m�j��%\�ird�o�ҩ�ȪY�÷�YҴL�/��tTUF��H�Y�i�i�\�0;��Ϫ�����3���wa�;#�ǈ�N&Re�it@y�smGa-�m�֍58et���U�5"�|��BR w���P�^9Uj�ks�e��L��ŏ��[�î/��	D7���pHWqi	�Yf�ݰ����S�-ǯ�O�z
�o�"���e>����Q��n���_w����8���C~���{ۯ�g��=C��{�1��~����$F�Wv��2��	"x� R:y��h� ��q�Kԝ��j<S�׺ࠍ�Z'�����g�:��u�(�m%��@Nh��� �a�3�F"�<�Ȃ���<ۥ�T�j�R󳮊N�Iщ5[Y�����Z�ry�g�� �1l�tB2�6��n��<�E/IR/�3�g�x��a���y���W71-�Ո@�����%DmS�k=1+k���� ESf�7�q b�&2����DfI�����H P�r�,3]� �����E�`�6�s[ziF�:��Y5]��"�4'-X�����+-�3E�h\�q�sIa��[غ�Š)�X�N�g9�_}k�AJ^��t�5��C%$���[/�CGa�����#t7��^�E��/f�1����"��Z�u�z�Z�cWp�D��Kї+��nYܘe����9
'��?�[5	�\{W�e�a06��o@��О(@�Q�aT����߃���հ/�U�����&2c��h]=�yB�k	�:��D�~��Q|`fR{xwǣ�\b�;=e��X��&�!�J;�)L���
������v$@��~ո�&���U�����
��g9dN�&��*FjL�<a�哻N�=�O�ad|��,�Fo��hW�{R˂�?���v$��gػ1�Ѭ: f'�[�����֫o)�\.�a��g������N2�	��+/Վf�GOWV��X�&�I�^��ue��i���,x��ʀo��pQ���KQ�����I"�jou���'���E� �o㷄�#� {'���۳2�)�5��گh*��y��n�h�ޖ�C��WϬ��VG�����(Ɍ�Jη�Z1<v+(����q�3��C��]i���c#[�A�D62>u
L�L�C�������a?�C�s�qHYvCX�q 9��bK�Vܫ��<����:_�}��$ܮ���N�Ν3v|F�����(������:��ī9�="�>���*of�G�<�h�~}q��4�F�Q�����9�{�������@z1�b��$y�`�Tcc�0ă�>%�w5�x�t���|W��)hp�����OA^&ח�8Dt����l2IK�݆K���9/`��轵8~�p��r�|�9{ܲԀj�����$�9I��9b����D{L���B�+��������Ĭ�	����O��`?؉�����κ�Y�dI�ҩ��Z�F����� ��+\hC�%�%r�1�ܙVE�=�tYݧ��N���.mq����k���G�zE1�'���Rq��r48��y+�AY���ڵF��;4����+dE"olZ�YR|��4��u�=�+>D��Y���,lN�x�sDuV�[:��j`���ؘ���LD�b�N�2#�tnډ�w�8Ў1��p:�jP�pPd
�5�{�y��u�`,gG�{�u<�C��<W��_��óA߱C@�g��T$ �"��7�&,�m2�kd���fY� A�ܣ�H=�/��e��jN���ҊH��	V喍�L������p��Ab�����߬�3rv}ťk	�$�᷃��"�%a[r��b��ywFB�m�r�	�`_��<l0ۏ 7�~tπ��A��F�{r����LJK�]��E�����8[g1-��ou�_�?`Z��L ��=�bǖǽ4@bق�c�	E%F�&��*��l�����3��^�NF/5qBh�Ք5ps����,P	����q�+� j�S�'k���~�V����׶w���%>!�m��@���[C�����l��m�sɣ���W��7@�>��w�_A#����g�|�N2�Φ�	9O� �Jl���M�>+����AZ�,�F�^W��n��s�|;��_j9�*�qv�C�Æ�ӊ�~����6���0��2Cí��B�V�"��ċ�s�5pܮc ڶ�T�<
|=%���Һ5�����BYu��/,y�U��@3�bu�ܝ��[L����D���+.I�{P:ca<�� ����+|�3c����ɑ�$ݩ6W������3�-4���L��T��d忰�}FfQ^F쭐�����jHOڕe�������a��Fg���nR�^S��A?)�Ĥ6b�/~i��Cdl�P`�f���l�����f��`�k˛H o]J|`=�n�� ��3�<�:���m�G歒H�h_7�i$vr�u=ｻ�з<j��_+$� Ɔ�^� �׎n�4pT�f���N��w� F�Qz���8�4����������ooYȯ��C�2��a��A��~�/6��R�#ע��8#ļGǫ�N��QvYǍ-! X�%�S^铵[P��K[k����3�:��o��<�'y ��{OV�e�q��s�n7�|��?��]���s��7�������Α�����"ԉ�>F��m<_�9��ߵ.G� ��/[�ɀ��?��s�v�8�L��eДԸ�9���$�r+��Y��ǗIUk��,;xŷ��@LN�H�[Ke7o��ԑ<-����,��R��(
`�_q;�d>�~�ǅ���YMH��}�LI� ���}�iwV�O��U��=��/]�Nǆ���|?�	G�J~�/[�H,�тP~Cg�4d�^"T�-#��T}�o��=��Z(���J�.�jq�Qㆌ�B�5�i)2cf�it��X^��2Yx�|/�I�@�����J��n�?ێ����Zxa����"������޶���D��ab3�i���X
��ݹތ�u`oGH-3!$��<>H7ո1)P�>7�_ 0=��~SnY�l�ޯ�mb��"G��V�m���w�����t�8���^5+��ܗ���`�;�y-Z��Y��E�� �n������Z�c.j-k�K����![
^�7�2�.(ߧ�9������gV~w�����N@��1���i���d�����A2;0K
����P�z�]�����l������t��x��0J�&�z��b����]\�jɰ��k�R�����ݐ�dc�F9	>���b��D\7a���}���u�,�ފ��W��SUX�'l�~� O�:�Aw�Ϗ�p�|�U�e8�I�i bhI��-�8�"�SA���Oʾ��V��Kw+�5����5������HniB�69s!}$ܕXg�[5n0�;*I���a#�j%���H�_��R(w��k�o����J~s��g���5�h8��g��c���J�?��IՏf��塼V���n"s'8�a�&�T�u��VԢ��I�a\�1gH�Y�Х#9��a]�y"�/�;m���N�d����
�!�v����w,A�TwA�(�%D.\�T�E�<5�Ѕ�:R����Dc���B���y2�N��+��1��l�f�u8��=K\�b���Z����"��u��|a:*�Ke_����:׃�x��f�ctR		RB�������۹�`��2�`i���42�5?{� ��27j��2�s������L���ً���Z������v�݄YY���L(צSvH�/h˗�o$�')4�[%�ʒ�8up���抯��SlG�8�e[0.I�4ū��f��R�/[�-i��2�aB25op��a-��(e��3��#�i� �"a$A���O�-uĒ�r�#$$���N�8'���)8���m���d_Gs���k�<�u�,6w�`'�P /�Ħ�+�p���Yps	{RD�m��Xr���p���T���F���"� �|��n&�+�c�[��G��W�@]�`=�=IV�ޠ�]��]�z�6�V�ܠ?$�2����!���Ar�6H�}*�p�:5_`��b�92�5O�z4�[����ӫ��44+u��&J-�������T��U�bÀ2�09�+	}�:nD�����A���u#���D�0�{�; 	N�@����{L�,�Пψ(�+#��W+=Cb���ρ�HŸ�^��2���ddG��qi���7PtE�qv�S��ܐ���v���ʓa�t-�Ťc �S'<P`��9����H��b�ZĪ����/�r,R���)�`�~N��k	+�����DŸ������]�L$
Flk"�U�����Ӓ���B�Wz�I(m/� C�3J��Umh3�'w��5.�2q�����MX�LP�\vEE�i�I�[Hf6�XK'���ߠ�B�@���i�6[����;�h`l�:�8��d�A��ƫV_%��R7 ڀ�_��u��!Ym�Dg��k��RF �S�S�?d(� +���&G;� pݔ�@BF���d�ǣ����[�5��0�Z���нK"�5�з��vt���u��H`����74������Ԩ7����A�ˍ�|�����ƨb�v}ƉBJK8MjRڗ��}�'[-�r��S��:R�����=�6(���X�8]9��n��8u�mǑ,7�*y bLC��o�[�����"ȳ!�t�ز�z���ԅ�Q+��1G�,��5#�7����N ���"�=l��A�^�J{�DQ���lͼN��EA�;Z#R�s�q*�f�����g 5�t��H|�� �(�[?gb�_v8t⍨9i�����6����G���4����w���b��mG�FG^��u��i�ݍ)	Z�B�ڒ���=5}6���'�r��)C��]�Ƽ^=� wŝu��-�\6k�i����isi� [�J�Ņif�ԖC��LQ�Bxm��1��oNA614rY�4�g3϶^��5#��p���ͩ�u�K/1�v�����=W&�r�Ƀ<oP>��/B���PP�����F����Bێm4�".,-�TC溰��" ��mO��i��фY�.$$��1�\O�xJ&P�x�Sj���P(��N*�3����:�zm�J��=�E�t0�ȧ~��Ηj�"m�X���E��>�9�d�M��M�����V�C���ll6��+�[���O�(�â+'@����Oe����$*1BF��p���%V�uO��
����w���3�7,?��	cZh�@�r>YL�ֲڬ��ST�[�mB�D�$?�z]�~��19��@sxGqP%p)�U�>�Hw-<&��,L�`��V�͎'��
�"Xo.�Tu��B�8ӫ'�����u8�a�I(�g������*J�h׮��c��էr�ڱ�8��	����Br�Md;�ԋsD��L�r)���o]�OZ��6�$��^�`U��FWC*m���$z�c�s�M���(��+�.Չ���c�ˑ?�N�7��$B�(E�g"~�8�uL�ʅ�o�D�Ȋ���>�� �����5:�tp��cF���amB���w �����j���o�é����K?� LIv��d��Q*��#F䞩�ѓT,��utD�P�z�vŞ����1���޵�`okh:���O���۳�)�#L��d���+�ƛ*�	#�| yי(~�"������H`�U�0��y̦H�(��l	A�B�_	�V�e+M���GAH%��sBdq�y����� ��`��/�/�(��iv;wH��k'�x-��1�C;�W��O�6�Ɇ\�ænV�[V��m��X#Ȟ�35}]U.����r[yG��%�[���y��9���wG0�T���G����	�7�2���� 2+���j�#��FD����u%E��PD!.�����O?�����3� {�_�@�Y��'�i�΄��a��ܲˁq����4��g�������^0�禷��۝I7��H�N�y6GX�W!��ɝ���˂L�qc�o��B

�J ��p��N�iO��NW��*�@�B��y�P�h%�s�=F0_�o�� �R突?u/Ň���,���ĕt9����Ԩ̟?���13��'���%^�]����p��G��/���I��I���,]���}��.�y�`��n�Z��.���|<�s��d�'�y�|^��9W}�Xc9Nd2|B��Z~�G�+�o~;&1���fM�R?/]�*�%bԷ����8�C9��G�07"ɡɧ��6���l�U6��{��oY������aN���b��G.n rFyF�Be�ݿ�1�;~@r�/����l�fނ��m��,{����@*��k�Cs�Y�����y�k��T�^�x"��k�����@���r$e��={B��k��K캋�nǵ�~���FEiE�,)غ�]y�r�2��]���: ֠��
Rm��}��`��^�F3���C,_�������\��26OʁC��{Р�{\k�B�q���4���t�]`�GS[�+Q�AH����S ��֒�/f�Ҽ��ʡF
��侨UCK)��������%�d����:���=�/�/�.��y[�0�������nw�BKؔ��"�W�������u
HM�f������$���ޓ�UO��!�{B�+&М!/|�l�-)׉���x��|BQ[,������Q���_��Q0�Z{x�c��4@�w/� )I�H�c��y�,�#Y� ��b�G?l���¹� ��M���S�M�Ps��3�8�η�;+	��:u@�	
:�z�m}g���3\a�>������`4��ƫ2w@�"I��Nm*�6��x�^Y�*�m�v_4��o�İ��u���#N��G'<@�â���TO��,U�鏇�h3����δ�'q�v�ǎc-�)5�mm0^�43a)��B�H��a���KvbƲ���[��tl�I+�"��z�K�á|�%&ݚЦE���������C���>g��c��G�/o)B�Qq[��r���V�����$G)h�5���`��ꈧN�|ޔK>Aꐖ����5���?<���ryz�ߨ� �2���.��0d���I�i������1������$�
�5��^�1���^#-Pj=7����r�S�ς���{��|//��)w[�lY��e9��(���Ԉ���n�Jh�n��Q?`�o��*0�F��
��wqҩ�j�p>ћ�h�
��:ڨ���5h��=���q��l�T4�-R�䗛J̱_�u麹%�6:�T;p�:{�#
6o���e�v�6bK�ky2W:֔��9O#A�3�~g������}S�[���(U���1�RD0Ym#�I1���]���:{�a�Z�`6ͼ�U�H�#Z|���d,�Ү�Ҕ��ϼ�	����%&�V'�EV:�{{~�|�B��Ёp<��Vx\�zQ�~H�o�c�m�Vcҽ�)������]�,V�0��Y	� ��Z~_��\��YD{�l����u?�f+���jW	k���%��$/��Ҹ�,�ܜ��'����'��=	�"��f����C	��W�k�u ��D���ˁd-��T )�����O�߆#bݲ=�W�ѥ�Qh�M��-$�c����;ƺr�9|r�C;�ܯP���� E�r�x6�{0v��L/Qxz!T��抔#���¦�k�-�|����q/�F�D���bP �#�6�Z}�w��Z�C�=h�܁�EMQ�\���CY�WVԋ�\�����鎓g�uT�7sd�-bE(�_�ev~�*tȴ��rI3����<Z�Բe�9�s�ʇ�%$+pD��e�#M{+���lT��8���V�g�R3��:�/L�&M�Z�^��`��_�tc/-ROC2a�Τ>kLG��y���Q[�sC��m�-S�T�w�^�]�[�U�&��L�8�+�_��Sf�3,"�Y��G�<�G��^Т�֭I� ��#��V�C�0S
�������W�Ai[I܂���@�PN�Q�pz�/��jA�r��ao
����Rÿ�6���#�ޟn�$�v&�M}�蹶R�e���W�\�&���k^/�?z��/;T� �$��X�����>	�Le�țP�;p��轧RꨒU{N��J�xm�f��"{s��K_?�p�e(Ov*��0i1������F�j�Ђ��j~���C����#&��c�0q�E%	��7���-sa��]���DŢ)'Y=4�?��|Y��� �r�odYtk3���{F��jXG�i���%0J�c��<G�p��Z�3���:�7#� ۼ��R��Ƒ��h�¨�.��~����*{��Մ0�Q�"SQM=[��D���̬� ��y���ę��-��[�nDx��f·�ƥvNPv�v�|:��T�Hދ8NP�ʹ	���	~�rà���ZL>�~�t��YZTP�^I2.��F�Ft?$yUt՛���A� ��hk��G1g�{�ԙA�,�[
ܥh*�h�4
���l)����3a@R`U��P`�{y�"9a��duq�%�����S6�Kf��Vd:fҠ[���n���b���r�p���d!�s��?�tG��
�tmi�_�u
$�HF�ۏ@@	���3/#�:��4`د.�;|mq�^�������y���w+ZN�ZW��\����*�̪(�R���ˌ�2h:��P�+f*"#|[�	�_��x��[i~�ø5�_���r�i�[`27J�k~�ٟ�E��E�s�D�׈�z܋鳧��{=�A��X$˒L�Z�Ø{q�.���>�Xs�:��F���=��������ft>��d]h��ч��~�_	��������r���MS\1��$���)����W��`E���R赙Ū3XM�g��m�t�n+�'��3���v*36%l�~CW�9���<�V�持��ء`����het����t�D���GZ�Ju�L9%�ؽ{:c��b��ցR�:i��2�@�I�8�� �6V�!�m�yU3�����ǎ�����6�����7?�ė'��Ỵ�21Գ��RQ��|%3�t�#�}p�0�0m�� #RI�j���w9̿�ю��T2�O���E�#0š�1<��j0S�K��)�%ꙫJ
�`F(/$]��e|v�q��J��R�jq^hoĄ����%?O�]y�+�1}ݚ��L�t����ap���N�V���{�Q0�|M�:�'�,�����"����z(�+�;/��/1��~K���G����J�q5qF#�O �P._�)'ġ�d�(<���W��`��a��Kh���H� �Z�6�q�[���F�Kc�ပ�':v��
,3RS�]���=�<��rbC$]�
BZ�W�n�c����ˢ�{�VH��z�}����Z�W�@u��3�rg'�t6�:���]����P�z���twӝI袬Ϝ��Q�ͣ]a�!�0�<�Ю��H�L���2p�@�l�Ѡ���-�	<�d̾_���{�4��;'���}rCg�d��:�����~>�����3\KZC�ܛUres��Ky?��xz�R�9�aZ0&BÑ҄����'�n�ilg�s�Xˊ����啹B�������T�{
X����Yhc��5!�.�Y���p ���M�0y%�h���@�>�*��Kp3N��M��ȃX�������� 5���a�T4<���60A�9�U!K��!�m��ɰi>,YU��<:����^O`*9���
H�P��� ]O(�-O�S)_�zx�g��ͤD��5�7o��8fe,�|�W�sS�X~��e�^��H7vIJ�h���0�)u��+��0j�M�5[��1�@LI�5��H��Y��>�$o�Cef�Ay��85��)7����/IDuS�#wJ�x��I����c� u��_�Y�nd�(\���4���dE9脻pdѫvB�ʏ���is+����\s�[-��>K���`��b^��J9ͽm&As#n6Q������i�6`�k*d���ih�ґ�Ԩ���M�W�k�~%�݁�)�O&���ȯ5F��+����&wk7.*k�sg�'4��]�c�k�~ͬ�E�->��;[8]��ڿ��-b#����c`��s��|#�U5��Rqrc[	�M����G1k���M�*hT�c�*�j�	�ė�Sfh7��pc|���jwS���c�X�2�ci
#J~����ux�e��_��1n+�� V�A"C�O}�bqP�T���i�ʉ���ΐ�����%%��8U�H����£2,�^��,�@�o�Rw��n�gÃpCm�=�w��s�#�Jn �.�ȣ���u����}���A�� ��c����Z�q�b�E��{+6���1���2��>/�xA�:ef��z$��������Xģe��?�b�ˇ���$��v$y��9 ��-�:4��[5��V�:��;
P'ҕ'�e~� t=t�b@2�6��8D��F�EL�6wt�Z�Ζ-׻�9�J���^���{ل��&u�u�e�u~��$>��T���š\���P�j�S�@��r�=�BОs�2�Sy'*C��n	���y3�ɸ������ΔI�WTl�~�<�$9�Bx�Z�-y��cl"rU��'}l|L��:o��e@7��8XpҺ؇3Zd��I(?��ý���2�a�U�hwz���Y����F>���U?W���E�~�U5�|��ʰW�>�T"�����DRT|sh4_�M�f�+Z��53CQ0g�PJ]{����L�&.��NF�`�Uj)r�	�ul�x]@�`Uf��`��wM��a��I?�"d��Gڜ_��������y2���:�"$?^�i�S9<�[?G�$4�a|�?�a-��~��03���)8�j.�XC��E�!��xpx�N�-�5DO~���~����*/`t����j�4�����a �L��@^�1�*OU�H�rR�����̺��]���&��b�/�aҕ�}\V誂�ʷ�]��2�*r�4F�d;�W�zϜ)"�:t�s9Ļw�o��9��M��trS��1�SJ"�/:�%����J�@�X4����������T���]q���̯PЂ�pI���W`B6�gnN��z�C��j<Y�̞q􆔿iL(����W�Q��*�+(;���K/F����V-�w�:1�IO[�j��z,E������Ⱅw��%ZW���ⲚfZ��PD�IJ3��H�}=��@/Y�@��GȾ2���~i��dT�F7kR��S۱���2�c�e���<�N�����Ixgɤ��A��.��.�{2�n�`ӹ}�|�L]���IV�����a��E&ռm���� �P��㥷p��?*����#�4B�jfG�}��1�d��'��Ï�s{��cQ�9���ϔ{7@�L�qE��ЏG]����tS�b�C14wR���<g��7C<�Mm�Z�^)i��N���k��%?�º]Y�5�Ճ7�(�F����9`kJ��-Z1�'*�hBt<�ޖ�ӱ�xA򽘪+X!\�Dק�G���'=1w 	�[˻1 ��Gӽ'sւ{ϙ�-��k�q��-�S��Cz�OO��)=̀�';��x����1�Q��%�s���h)�i�8��F��} X0Sd�M�2)p�M��}��ϽZkU"�B��>�[����ARvū,%�\�ǈo~E����\���3>��a�a��cr�����@�����t9f�w8���@}�`_[zo�����"�PKߩFK����b�*��l{ʬ����E�Y�T�
Rm�+��[��勁'Us�J�a�}���'��(���*~��|�7W�U`Qm
�?_^�{)n�Lw�����ͧ�Z�Z����X�tO��z?[-5.��a��z��~�	0t�f=�r��O��u�U�]�2XLf���?NB�L4�gM0�/<�6WB�ѥ����4F �a=�F��/�` ��˕+c�������{�aS���08���B���� 9E�x����9u�$,{�j��mO�'y�za$^Ğ͟N�K <�������gԽ&7���*C�d[ٲF�HA~�i�{�{�e�ʊEB���]��7�Ul��U_�_��#U�F��Q`}�ªNv����M�в6f��)J��;v��!WE?�)��15h�FbZF0������̘��/ըC�m�����<����x��^D'���m�	o�핎k�5ї�Tbc�n�w�1���4p�(�4`��;d&�:���G��P���8	#�@�hJx�ոA�
��^`Fj��b��[,:$f��l�iY�?�^�xL��~5�cH�S;<�=[ϓ޽�e���ˎLK�2�	*�4(�U�'J��W z��a���Un/�.jYq��^�_)�Pt<iG��
{���f�*y��a`7��?씟Ki��0ֵ�3Z��V(��^ 2x���M�E}�Շ�2�E���Iĕ�`y�l�I]v�P/���~�S���28ҩ��k��C���;Hr�W����ץǒ�+�H4$�|��M�Ξ!��a*ˍP[�n�X$0���R�r�k���g�>��_����MQ59�Q�o`�&�6ƬN�ԣ�6
sF;��XX�������Hg��k��m���F{}M�8���#���v��Af�	Q��6}��T�O��a����}���<��~xiq|�IQ�c�%=�|��N��� @�j6��j~�f����a�h�H��b������c7�s�ˏ�Z@� �/H'�(%�6���!�@�[�#4�����H�zF{�����$������7\�ݐ�K����=���V��)Wǃ��Ҽ�&��MP��x��M݃D!�-�kJ�s7�~N�E%��
N�]����D.M�!_jJ�+�mr��I� �u�GC���p��H��i�*t����1���X�}�\�+�����wl����?�͠�����W`f���o��O���dR$-�f^���3��h�sR=<�*T������F���<r����`����z���
O�x*���+S�R�ު�;N��,�gR�^9D0h[&8fBµ��g"�5� Y��wӏz����A�l�&d}�콎������]�H~1Tw�a1=,o,��z����#�E�f�d?�bj}��i�o-a	Q�K1���O1��|�t�6��lM
����3�瑒��2Tdڶ��'<���k��Z�\��ɐ��I*+nvK-�����i�&fX2�=|'�^5�ӡ�A�/��_	���-[{.)�K�gg���Y5�x��
�\�(lnT���[�������+���
3�x`�iC��ܻ�a�� ֥f��I�4#�"k沥&L�)	���/?K���d|�O�\�,�U"����$�o؉�mR����`��`[�����~`&l+�Ͻe5�
�	����=�Pv�կ}ѐL~d�g.��7�jl����إ*�,�ep�L�C8a���\���2�#��������P��^�U�~�4�Y&��EfSr���eB.]
E��e�j!�o:� �E21�|+}��YQ�Tc�M*�c�r%�>����d���3�ZЧ:�:.�v�{�X�_�1����Fr5Dĥ����Q����*�m��s��1��PE�i�w��h��z;�(�|dm�m��SX>��Ì3�t݉9"�g�(k^I�R��d�aCb�/�Td��g6�KS�����K�i���*��"E!gy����T���
:Ի�֫�K�v�B[�
 Wt�-�}OfS�xB��Hz��]W���gN��_��)��R*.�*�<�4�/�q+��qv�ǉ���"Ѿ�o�!C�J<��eO����%5�30ӰS%I�6����3�t�ShB�W����L�gQ��D��!�Z��,N y� �sBZ�9N;ơ+gEe*2�G�`�P�k8`˰p����U�4����m��P�
�BCz�W���L:�Sc��2�I��W刴ꧤ�u�<~����x�Y�a��^s����t�TG��=��?P�����3.H�O�T��|A�k���u�g���ն�L4Yܶ�{S��B������� �C�������6�,I����a��<[#���&��(fg�.�+7���C�ɍ�j�LQT����-b�PQJ���̗�����;�ܻ�ς�5�w<g/Sf�CSI��Ƅĉ�tl�$��w�ȉ�.ـ$-ʚT�������+��Z7=��}�9U�Nf�!�Y�����8]����g8x�i���T�BW1`�w@*�����w�P�Ea�F��[��r��+鑂e�����5����P�+ڥewa�_�ݵ�Gf��t�ս _h��N�8�(s =����q�
���\&5�YH�gsl6s�� ��'���:ff�5-V�,����!:&e�
n�h��*
��x������b��Z��Ŗr�"c/0�����*��Q�\�J�.��2��c�N�r[R�=#B��,�ɺ��Ӌ�f�Z�Z��ط�4]^$��\	ݥ���4Z@�~�P.VۛF�V�+B��y��5��f���O�\R_�V�xSG6E1eͣ���v�_.QY��c�7tƃ+�K�`���������R>k�,��1�|�$渾Ye�dÏH�2e	�P|���cS�	��?/O�r��߿��&���~ �i�K4h�Ji'��ޢ��5��0��k[���u�u�|���j���wk�~�(��4����g6�r����e:��
�����s5R�-�� 9F}��Ie����\"��bn�c���( ���a`�"����;h��T����ͪ���uP�ݎ�A���<;]��^�o��^&���0�J�ĭ�Q~d=�Q6�=�O��\	�����n�!n��w��*j�Lъ��m��1�&�\����U���B;�}���[T5��`uZ�Y>J������0��+�li~��+�u#�h'Sg��X�!�Y>B]wϡ���$�B��= y�������XWgTƒ<='���$���_)��H#�ū�j&%�x�P�H=O��FyǱ.o �8�c�����͹7�ѩ�:�D����AbH|�%y}D���
�^	=m����ݞ�<@�H�uj�'�K?O�ZE4��t�+Өg�sU��h�-�+I�R��[�ܰ?}����nS!����V����3��OF?;V���.+��]�'��q`��6q��n��^��Ą!����pі+�A���U��x�pMC�E�Zr�Ӎ/��#m]p�Ѐ_K�Ր.��0�
���O��r=��_G����g�8��8×��[Ͻ"�F��4���Ŷ���Y!�쇗��M˥|��BQ��quI#� eG�Y��7"���ݴ��0a��1��ER�U�9�	4���7Rau넰w���������>>��l�[�_����B�h�+�a��I���w�?��jĢ���cF"�yf�T]L.e,Ki�<hp�*�ۣ�x�����- 2<|@��Q�v� j4SU���/V4�k����( �m?88đ:܃\�l�����L�o� �v������3�����6ƅ�V�H�bOV��$�����S$�J�pq�m��I��+)�A5'�v}	(",��o&F�0m0�������$�Q�h ��t�i ��@Ɋ֑�d���E�+��.�Q	-A/`L	���t���X���jґ����6B2�l���?�D�t�\��i�'ȤD�G��C�����7�PcT#�)�c'����m�X�����O�֛A���(���:�Q�3�6s���] ���]�C
�-�QP!�A~F�L��9���F��,$����������˚ݺ��,�)�b&���*��
,�zIN�Yp�mv���eNT�U�>���k&V��QF�Μ~6���7�7Q��hc����D[�.G^!�#�4(�
L^]�]���q��Ab�u��Ӧ�'c b��~����m���6�ZACI��5>5��z�`�`�F�	��i^|!�����HqO�Q�#]	`l^�`�.-=ǡ�Rj����AƠ	��;���.8>�7�(xCM��P������Ճ���0���(A�lH���Z�@�����Q`G��}�����FG�v����I���^�����f�������	��uڇ����\��B~qx���`�X��4(=_	.S�0�C^#ܸ>X��.��1L��}2�2���cu٦4�ve�B>�D�?"
�y�d�.�� ���(5�����Iz����T���ng
���ى��7�ek]z����$]h
���OR�k��
<�����vH-�*�Q0��Rt�E�OWkUV^��������}�V�w����w��q%B@��Sb�/~S�̓}g��R �����GA:dz���HcC�!ʾ�~��P�X"��A�p��&*�c;�>Zn�c��a�EK�8Mx &Y�ڱ�"��~ķ��Jʔ�d�I�栃���5�s�͍|�d������,�@����\�3F�����ԓz$�F��F�\�<C',R؈JM������;]l�G#���v[s!}�@�D�c��<��@�����B�����m0�,�k���!gr�ǫ��E��p���u��_�"������.��+-�+\��亄n���]�A�1�e5���ȏ ��ઍ6��E^ �
2d� ��{��Y��]�qâ_��!��c�.o�B��rL�1t)b��x����Bb"w�=]�s�؇���O�f	w̕���'��~����\��L,�K�v��c���T���q/ͯ�\IJ�*hUL�/hK��ʠ!�j7�"�%�\yyracb[3�����6'�U����Rw��*�����c��o�d|���,BlĒ��Q�e��+>����9�,��0��:vM906\&�;���t���hW2����g��b�r������X�;uN1���QAz!��Bai`Ia`JM�b�6�7he�s�taW�9�F�Fq�ރ�B��yi�s�N�'O�p(�܍��@=m���*V���d%�.���RNTv�b�r�x�d��WY��

�P�䎾c#Tp#�!6x�S �oR�*�n�<Ї�� �J>1�h��'ӑ3�3�P�&=���5S()�4t�w�K�Ɣ&�H~ɼ֏BP'?������ly Lp�]��W����\�,7�I�^���m�\ܮ9S_z�ډg�"�F@�ݝ����#+��m���lI�1����&H­(�f�2��κ�AD�#=��94!Lւ)�S��-S9퓢d��7�*�EG�e./�;��q��y��|�%{ì)��`�43�6�-\8O(�r^5J�y�+�=���+=\")IJCܤZ0[ åM)Vv.�ToI�/,1���m������K8��.����[H����Ք��o4�m�?m��I��W�2���ou	����6!1&�֡I��(�����$��f���w�\��3�K��}�{�S��Ic��Ǝx�@O�"Z�}��o�W�*w �Zq��t�`���d���J]��d"Au7�فVZk �vCHX5␉�|�~���U����?> i_l�O���v�����\���:��)�Z�PT���Y���,�t� 3����j�X���	R�i�D���Q�Ԁ̬8�iw�,f9�����
 �^>��|��N���S��E�CoA$�>PD_#�z����V� �:x韔��O2�X�\�wih��a�jb��'����:�n!���w}�5o���D<m�4	�{n���5ޟ
\;�T�s��������L.��k���.�M���0G�.������U4�b0m՘��/���tђk$��ߢ���5�?�������v�a��u�%k��^��t�8=#��|ރ�Crؼ	�t;��T���4~��#�h��A��R	nt����}�(��Xt:����m��:�y��M��t��;�7��֋�<���z�g��G�v�6��s��w[���_+�GǺ�?X��:w�i��uޅsf]2��Ӄ�:Ѩ+'�]r�-�mV���ݑ$3�M��}D+ZSrֲ�B}�C��~�Ѓ�_~Y1zp]Q�3,�^�8g�r��0aTݛ�<���i'�O�����V���~S�N��J��?hm� N	<����=��J|J����u(�6&��8����ؼ��8�dLߕ�j�ӮV�Q�Ր�/D�Y�`sSC�)�R����#��ۥZ�;n��C;X��RC��?���_9GB��K$XM�W���8;_$�n���c�t��6�|Y�v��[?t��������?v��\�,���p5��=��u#��я3��A��_G�3rm|�m�u��TO`��x�<�����a;�Q&8\A���f�D3�!<5��gٻS����~��w&��qBcs�+;����]�b�ŊD](�>�c�!E @/$X�Ys���[�Oµ�����v�Q4����v��;̐�;8yH@�LDJ���"43\��[S)�0�p�/���mK�$��m�+�D�	�����5����}[jI-~���e�Q�0���@��;��E��de�1q75�==p�溼��5:�+8N�D�i4f�zB޾��W����t�bp���0�T��YQ�Q��F�iX����y0H���P/;'���9V�>�q�r#���?�~�!���q�������1�~�4��6e/ä��{ ?��f���
&���Ī����lȳ�����h�a������{p�L�X�vt�5A��Ј~Ԣ:�0b˦? z�T\�֒u�)-��� �Q0���ķ�^��@�����e�����=�;�4��x[�TE����v�blㆫ������<=a���$���:���Xgh�h�Z��H���}ְ)>��N�a���KZgc����=rfh�s�.�F�h�K���+��LǊ>t��{������tq�G�P�u�j�%x4�g�𛾪]�#ڮ�Į�\��[}��tӖ@���ő�������.R%�?�8N�m�R�MU�D��2�g�j� ��5|����p�;��Ѝ�GW�f��{\�0���C�d�X����-$��*i%�J�C�N���hB��'�@w��:fP���s#/}Ǫ,5��#O�z�.��D��,������7D��Ý�A���vP��9���x۸�����˚� ���]Ah�ǩ(�/��?��3��ё
�����R�>*ow˔fhmB�{#V�[�����P��1���H���'�	���h01��쳶��*�ک�x�/�_�*n`�9+�!Es`I���y_u�1ĖEj�~��N��r=�;�dJ��?=���9	v{�r��[C�r\�Q��l���[��ޖ��5�n
-`�&����P��-�S+�(�i�[�HV2 ��%vЀCu��w�����!��7љ6a��J���#����͛y�6I,*�F$zڵ��7\y�찭b]׈��ƱsI�i;,��i�*�z���T�����1�Z�'~O��쏓�p)-�˩�C}�o��^���<��Ji�����}��7�;��TvZ`��,������a�'U�����*8)�:� �! c�>� ��nԽ�67c�m��^���bP9:���O�U�8]�g����%�Lt����U��W�|�@&�!�6�>�ǀM��u�/d��R��p��!���]�3���W�|.A�mV>����W�Î�<ms+=�}�N�E���y�3�^�\�̓�靸Pŉՠ&��P���O^=�*��"��h	��
�J!�w��\HrF�:G���6Ʀԭ]?#]���G�,�^ ��+�3�>�_K�{I���)ZHeO��fs����L��-��Y�
�Bq8f`�x���r�g4l��
E�^I,�:m��Q��&�G��4ըά��5D�R!���9c�v�K�T�'B��t/�
�=<,n G�p��r��ӱ���~N�׉�!�������p|�2i�/鐖֜	�R���j����HsD�=��P�g�(}0eK��5���C�U{�Ln���� �UD~�S�<��QuVM��+��/ɤ� ��-wݮ_|p\k����;t�bHw����ק�CP6�%1�	�C w�ᷟv�V����$��@!����*!}��UEG���Xb;���.o۸iN�*�c�������k5RҁY`��l��3�B�Ø%*C߆֎�p�ʝ�k[lF��X���,n���hO�����v�`��IpΗ���#Cxa��:�����V5��m-�Z���ii�S��#)����n7�H���g�=��V�H��0�_�!�����Dx6>�(�����s��d���Y������4.eL:�6m���L�����::M# aBOV�i����i&�5�a�M��k��39�k�:�-���`-6��r 9�6JH���ȕ|
�n���|д���4�$!Jȡ���-J�%��|�AnG���r>N��ݬ1���/PA��`�����h0
9�'��� �������ƛ�%��P��5��(l���lJ� ?�$�{�cf�JW���"��d�X�����a��bƵ%R�ˌ�d��R1˘dCY��{�~v�Ti��F6;��b?ԥ(�����K��8m^�V̱?7��<l��#r��f^p��nh��C\�$�\^�.���_��h@�����'��}'�#�eB���kI ��"�5��2�3�y$y���
�=$��,|�3k,�sײ����	)��"�5Md�3II���3�~X� |M�?�kی}���-I*EZ�T./�ʘ�N=U��ozlE�${��	��j/�\Է��a�����SI@`�e������l�8� &wpF�3���'�K�D!����iUaz�V��[�Ֆ��V�q��L\��^6��qݖ_��K�w�8ީj4}��<p�K7����^bV�"��֭-L��~�C�=�~���zV�ݼ�
>bma��G���� �k�x�G�H�ᒄw:a���o�a3mJ�NZ����E�m��n��vW��r�@�%Z��������|�`�:k�m���:��z(���v'�����E�;�q�;����/Ă>��- >)����$��s��*�Cǀ���)�跒��K��tZ���j���3�`l�%
����O������}Y���s�jq������f����X���onջW/U#`��h*
,F|���qo�X��'TW�@D��@BF�؉*y|�����_�?�p��"/����@�.N8��@T �X� *�����V�m$��4g�򇐴����a��>����	Xy����+��k)-�X��q��sx�jOM�< ����$3�,��?x�yEsdƤ����F��:�XYt;���nۺ�Uu?��`>C�ﶬ�Hg0rj�(���A�e���@���P�R�M�յV?�r���[5�F:���=6���l�5K�� �>�{�wl����!x_[R�vIʻ��V��_-�n�6
ϜI�u��q�:��Hp�
�%W�Q����Kz��u_����<�n�͒�~LI��6�˙N��Na����H�/�V����z�g�V^��qc\���9W��:��2G���b0�$�&�PS�'�j���T�E͟�	]�V�0Sb�X	y�=>۞4���u�c���� !�O0LU���������G�e�e[��3��ƀ�Pr6>�:��������V�������hg��X�����t�_�S*,Ȕ��H�/o2+��|v��wQ�V�Y0�K�U���z!���_z�w�ð2�23��n�x�1�+�����k��^t�>։b!_���{]��a�����y�-߇:H�'y����3ge�7<�ɲ�苚��8�I �|���E2��-&í8��E������SxWɺ6�|_c'�|¹eOv��_�ѻ@~��ͺ��L�eK �'u�v�9�!y��<��k��t���q,S� ��O%q�0���B�W��fe���LoV׏69��f��*����d�q�l�/M y��u�>��N!IH�Ĝ�`)溡s�����9T�P��[l��E�j�������k����Y7$��u_��Wr$��4�˝M�	o#
2H(D)hAx�ͥ��uG�s
��������X�5�{�ۘ�t�/�z׎^�\G��\7x�?�*�����c���	��.j��WψɁ>����%�z������x�I�L�~��8s���b��f�H�k�	���������IU��8����1u�,�7��
�џ�]��Rks�O��h5�lL��}s�З[��k��N�7I��J8�.y�r�b��;��뜝�w3�VnTv��HZ�l�5���ie �3 �G�'r�Y�N|��56��������K10�o¯|��1���t�he�\�gK�ZG�lbh����k���:92<��I�ݼM:/%��O�V���ǠVۭ���'��x�Oo�ٔ(0����Ӯ(����<HG�W���ۍ��8�5']����m���T�=��K�؇�g�tO�^W�c�۽l �`
�_�˚��#��1f���IڣP]�8�O�G�eN������3��P�l��+*�gl�۔'&�n� &d���ykUc��ޝu�S�k�c���GsnI U�>`c�/��&�3DA����m}��A�W��7�`��m�����H8����6&Aʚ�iKl�<H#��g�<��g����&�o�_f�R�M7��|0c�n�*��?'�v(��<*�O�X=8���	Z��_��+M]�zb�s.y��ȼ��81
R�:�H���r6�)��PV�O�ZUc��m&4�ҳ1}WPK�����j��ö�J|��}�G���>yۮ�15?f�=�#oi�6u�?,,J���L�=��~q��
����=�b�{�v�t�m���41ɨ&���%Dx������W[��a,'#�����y�2=�p��G!��(�S��j��q/VfX��\5���mj����1�O[D� ���
dعw�$��c_�7��H!>�
��x�:��� �\r�rу^�<��z>�|>b� |W"/�/1@'�S�mse�����FJ~�l�r����	\tav��� )�V%�|�� z�Y�zg��O[���������i�NiSء�+���Our	_���K� R��E<V�p14�t��@��g�^��U�L��$�������w�5�{���6�]�Sl��.Ȫ�����*�Ϟ����S8*J�P��WS\o����<a��pHY�;������%�����{V�5��-��Ue��f�6w��'�7���ƍ����ێP� ]?���Ͳ����FJn�iܗ�q Ǉ���e:�в�c��J�{\�9:��^
���2�
���Ÿ� mkN��D@t���zk�z�lÎx���
ȭǤǮBn�����'�*2�j;&F����S"W��$$7��:��fRz�h��슃�۹��mtL�n�vԅ��v�:���u���Q��H�x5@B�wگm����)���ґ��j�o����[6�7���#"q5�3�H|}�Ѯ����3��XJ���~�I*ȡ�s�����凔ߡ���RQ�q��o�hs�D�U���`�5p�V����v7��/A�Է �FfxBd��=+"_;���1���Xc_'':}�k���j���%���+!6r8��j�^�D`�&	�v�K$�C�l��u��u�]:�P�J��i�r�DN�КĵToL�V]5l.>W[d;yW����u��gb�"�(�_~��#���	�}LA�_�]|����9P_+6O��c�Cu��'�m��O������YŨ����$Z<N����%1p{���SR)�j�ZJ��C��g�I��A�	�]���7����P:�Yn$/z=��}���{�%׿:m_%���ށI���m�U���`��+�_��Ϗ�D�ɖ嬦���4�x!v��٧�&��x(oy{Ud(��fvUT���s�0i�����D7o�pӲ�����ZQ��+�;�T��M�6FX��j��ǆ_*_�
�Ն0!�~�+J��R�^0��g	���4�<c7��a%�Q�*pꁕ���C����_�՚Z0P	K������s��/�EP��ز绵#����ᗁ;�4��$bI��Q�����&>��&M�>�Ν,�/�J\��9��t#��^Y �~���5��&6C��5R�dO
͗�{�4{pD�X�V/v�O?%F!�4q�mE^�r�Ɨ��[*�uY��)�@J��u$t�f;�z��4
�Z����F(�yp�b5`f�gL�Գ&�F��y���^�&.��v	��k�˼G��-�(�6��>����e��꽬ᵏ�3(��~�շ�p�2�Mؼ��0�T؅��Z�v�~�c�^&�tvsі�3Y�#���-�y�Ik%��nS���=gb-�U��M:Won~�ގ �ձ�,_d��T���.t-�O�Nj�H�b���5�F˖m�OQq ������{��zɀ�������;pW*��K\�����w.�VY��*�{�p�[�$� B�,Zm��kx`&�p��z��ғQ�˹�̥/��ǋun��Ƙ	T<�j?+��F>���Ed�㷬�0"=ǩ%�	W�#&��V��A�'0p��oL���#QiV�� �:�H�ҖW�2��</I��d�5�)sr���'Qf�^%��4 1�H���_H2�*�b�G�ip�m���w�hYx��{��'EfY�lvdnjR͸T��lhA�0��S���U^��P���ԎD:]�:XN���뗘�?�K<�s��M�-�gw������'@2��p1�&b~���(r�>�c����O�+iwY
����,�h��PW��(�1b'�jP1%\��E�������(+\`?�'��h��i@ӅH���f���̢�L�t�����>�-�4��<�bc�%0 A�b,l^j�ٸ~׵�d�y�3PTȆ�!��tZ>���PN�ý���D��K�\=v�z��8��������T�l`�������G׼3�y�˺�"�E��f�.�b�����������ǯ�ԥZ��&{�G�|�n�F�K�������D}�˹ �ƃ��'7G��v
~��;򷲪��[j}N�Cz��(_�O������[��kg<��{�����ﮥ�潹
����l�������ě�e�=�ځ����*\�%��1%xV]z(�	�[���ѧj��.�r9.�Y�u��30��Y՘t��d�� ��2Ϋ����[�m�8�Qs�o�;:5H���҄�@YOx�s
�)]���ͺ�Ύ��z2Y�ɱZ꼻����g�uv�.�#�~#B��͸��ܵ����@ �[	��-��U�\�#y
c~TDQ�&�81j��k����e�%O(ˉ ����ҩ��M�����a2Ff� �\�ih����$��&d�M@D��(�Z)��PL���eE�-L�b�k�U���G�Ņ��.0��$��("�ot3�zL�E�2��"m}-��_EKA�?�<�-a����I�a|gE�gPP�d�l�����8~�U����m�}��p}�e.�F��n�����d-fjb���,�.Ѻ��'��~#����&\����;�]�v~����f��%��0��㕇1/��#[����'�c��3�z�='��Dh�n#FG����o���m����;��hI�۲#>T�z��������c�f��\�_`8��FL��<�?���e�Ch_���7f��#]1A��l�FӘ@W;�k�^@)`a�Ē��W��$<�������w;����a[Uq�q	F*3����|T�H�)y�߭K�k� au	���Q�1ӬmV���kp6��_8��#9Vy��|�J8N������ՐĞ��-��g1��,n���=� j*r�D현ˮ��e?1P��Ѷ�ȃj y-D����@,{��.܉6GN�O_�o^�Fh1�s�;voO~ת$R��MF�~��B׬�5���Tz���!�~-욗�_�Π��А
���a����=$e�/Y62@�T��i�Gq#E�M�����e$���<.����Z�Ve�-�'7��]��A�W\Z����� �Wk�A�uQ�خ�ĒXD�(HW��PQGtF�;r�}A��/��u�d�F��}h�����>ş��
��ӁP��㌘���V؛tg/�@�*��#�$��K�cz��|;���^��y�/Ɗ
�> �rd'�'�
��Ř	���1	�PB���*�l�Y�.��8����%,eW�~��ʯ�?�HA�LC̅yh�a������ktW]����7E����v2��G�qW�Z],��pl�O���7k��|���pS��Ѓe�����|�7��q���2�80x��K�[���?֌_�dT��ꇿ�[�|j���{PDKˡ �L!�@�
����Ȫ�#
��p�?������d
�e�>�ࢯ�Y��''�kPz��� 9V����!���lގ|W���Xvh���t\ZC�/v����L��X���0�A��Ù�2��5M/�3��xy����#���^<���.���5���b�{ ������U1���q�����
Ѣ;�]�2���������Ԓlq�L��C���qv�7��7o�X]�Iq�IDq�����%���D�͞�xʜ�u�������w���'|�rl��r/B$Ľ��G�]=���,�V@׶������\�s+/p��� �S��z�T��`C~�"7x�V��N�ē�H�s|�L�u-��_O����c�JώW��p־� ���{�����pg��Z@�z����Db;Y@�!l�?�7P>G�	��&��Vd�	z$�a�[����vd�q=��XN&���B�-t_�[�m�Й\%B�t�	ԃo��m�=�zʰ���Qǥ	�v1��j�֬�Hb�<R*�ϛ��ۘd/=M:�,�U�		!���kq��vV�BK2��{.��lO����D��X��fin�A�A��6S�`�v�`|����"��(�\���(��y,��(Ɉ5�VJ|��3�]�%�z��ǈ��>�Qg1�D��i|�|�eű�.`�)T[)�%J�fT=�X�˩�(F|�^ϓ�s��c/�̫��'�Ƞm��(.g�]�9CˀCDY]��I��b��:�M�p5Iw���(k��TVˊ(�˻u}D��p{���ZJE�;�J�|�y��P��^�Սq=�zEr��
">���(ke��(㴛�pU�Y �:�l]�q���-��욠�Z�d�Gk\:4���ix�5����XhJz��>+e9���m���V5'�l�yh�`��#��ݲ!��&�۠��s����#F�D�c��b��F8����d̃JG��3[ ��ɸ�"�3����0�-�(�x�ߝ$��x�U5����>���Q���/���T.��N��S�O����d��g���B���] �#`z)�u"����Mu5p8��1���'���:�x� 7f'�$����@�=�ݾC t��CB�K]0��m��z������Xε���с����s�����bxЙ�~���6�N*|N�@u���K�Fȱ6|I�� S9u	֮
��
���mӃ����3{�2E�}X�٫`�X���P>�Z�&&���� ç��	5�K�r#�T}��$��;3B*�t����~ w�!
�{�Dk:쁽� ^�e"�˘^��Y��i1^j%x�"$1��PP��شu��-	�Ɋ�>gwl�-�.���RY���戞��"�
���X���G��~�C �PDO��ľ~pT͒���y�����<T+��	�%nrǦ8�O~h���K_�ޅ��-�H��u��g�EĒ��λѧ �Q]�I�>1N�9��0� �3����8�+"bX�"���n��EKlN
~&�):�V�k��E��iJP�p'��n��i-N���eq�ڨ�٬�m3�͇KU��H;20�ڈ���NT��Oa�{�B^��H�a��'���`�˄�*����vRԯΣ�q��KP�5���Z�4Ը<'���h�X�W�W2��HB���roa�@��>�f@q���.��N�ߢ��S+��K�1(�zG�K֙�jO���<L$y���KRNY_�v���|t��[E&Цʀ<'"���D��5RZ�;�� �aߤ�+�JNT+�,�"��p�x,R�,D�8��u�������]��`�+�{H�
�iU (�`���wY۶O�x����ןA���S�F<�he"5;��.4X�f�*E~�K\�rjƸ=���g?qN�R�.pK��,*]ch�r��"�o�(��������+��<�>7�ˏ-a,(��)X4_i��%N
��40F���xÑ\]-i /�K�YvVr7��Bj��-q�{�X���.�ǲ8f �'�sh����F$]���*ұ��92xe�Mo')����V��3?0^=�oPVR:�X^*�]��+`�w��tj��s�-�`���;��j^�M�W~��Y�"�|i�F�*�H�W���a�[\���`ި�$��w
Z1�Z� ����B^���.K������������q�|�;�vwU���QF�~�C*��^����`�7�B�>!���h��b��IN����ۆE�1k>/�7��??&Jh�TG9��M��ڊ�gq�����&yĲ%��i�/�8m
(c�Jx(��xG�S��@���^��"�o{�҄Ax��X*�9[w��a�!�^�@��E	��4�."L@n!S�l�N3��5x yk}�c6���C8�����(�@~U��8�U��E��D�3���(�pV�<ۼ�u}�H�I)��4jea�E /���<7R��݃Iv��6PE��k�]���Af:g��T^���Ak�^ك6Gy��� ��J�Ė{���~/�:�v�L$��c�۟%��n���6Óh�  �R���{ţ�?���k:��`�`�j�& ���u�NØJ����0�H��9. Z�ɝD:�Ղ��ڶw�Y�کI�����{�S�������8��-J��q�X91ͼ�b2��̅
7��;�y- W���P�rAxU������Us�J��C�x(_��#	�v�>Ȩ~��Рǅ;�5�O� �����.�h�}��ZD�<$�X�8�<��0�XO*Ŭ�&<����#�������m 2d�&aQ�����ҳG��A�-��2,3�Bf�Fb[!����{Z�\��̩ۧ⢴�����%�K$�W���?�U���[�i]"bp8�K�éㅺA��r���H�v	K�r�3+ܒ����r����	L �o�e#t>���m^�1<e0%��#�[fC�p�O
aVڰ����"��'��S��sff�-����N���B����b�������u��alI�:���ۨ|
�Uʤf�e0V�n�fD3�Fǣ5��������6a���q��,D �U�'�AXߺ�[��G��g��{Fw���!��͋�(���Xgj,�m�ud�
�p��	{������Зq,���|����`IR8��O�P ����Ӽ|2�<�Q)*^%+C��gQ1����y���&�o������!I��꽟�3��s�F���K�?���Ȩ��@{)��.%�L���{b��D����B��-��=>���_`��F���eR��zZ5��>���&�#�?�6�S��݌/��h�R�hpl��qӘ|=��9=��rY�M~XO��h4`+��;6��K���3�� �Ӯ��F��Bu���vr�������u=͘�`�U`���d����#�;�Ǧo�L�fi/i#�%l#����t�!�xg�Zq���23g�";W�kZ��H.�	��k�"���5�G$�b �к��(���N|X.�E�6����G��;U���|˶�:<h���l��l���!N�hq�V9��A݋l�.H @�N]�J��^iO��'�����<QT����__����ʹ�(;{�v8��f{`���.��/GO�1���)B�C>�9Y�f�LXЮ�G�b��!��� �*�~�ŕ����f�����zqNý��]�\���<
�xm�1�v%<��y� �b:am0I�Ji�Ɣ�y�{��d\a�+r��ڟ� ��|6φ��i`�L���D��ErA��k����b�OO�)�
���(��hX�;��a��) ���o
�-�sFn��Be���#td���}9�A���������yY��2��Z���4��ƍ�6��(�[ p�<�'^D^�n���}/A�!�E:ܡ�C������tu�[\,i��g��5�oF�$8�Lj�d� ~�#8��ı��?��,��<�� =�-��AuWF�f�s�/���J�L6��xֆT�%uI��c鲏L�p����^�����\i,��U� �����8]�k,�_�1q҄5y�^;`(-Q2É����]0�s$oej�a��}`7�N����*���s�(Z^�!PD��¿�-'��x��i>aA�:b��9���9 ���V���y�	�ՠ���NgU����������L�@Q�bݰ��Gvm!P%��9�3H]pVu
�]oSB�N����Ś��c$,�(l�!g֛�ҧ���\�n���~?��f�2lM_1}!�5�J����9���P��iJ��rK�l�̘�}�󮔼�j��d��Mׄ�ow����V���1�P�W$��#��DV��y�����u~觡Dbn����427�$)�`DZ��e��}T��?Tķd��S��6���U5��F4�W�*�����1ZWŉ���Q��S���旆���[���.ivf�i��2��['L�4���{ȅBQ�g6??����N1+I�B[鸕/���1�qhX"G�:���HjB��=n��Lm.h���71Y�[ɳ�0��L�}$�?;�sF�CR~_l�A������L�@'�/^��l�62	i�~�%��pGQi������X��1T�xؾ�o̭�"p�_���h��v������������w�
���,d���Fe���+U�"���3��|�z-QU�Qucq����l*��u6,9=ȩ3�ɎO�\<�'��D��i=��xnz�����v�T��Ըy�*�/ve�N��W��8���1"��5*4��B�\c��x�Y��(���E!�d*���X�)&1t�T�?PT}C���X��a�h��ģ�z��U�u,�Q�ͣw�x��#5��P9Z���ce�H�DF bLT�/�%,���R�wwR�+�+�7o�7���hf�;��*crֻ��W�8L
�g�g8B�; T1��ݶ���E4�$�q��s����p<���3'/����d��?~�\����/�gl;�g�5��Xʋ��������U��� �B�@��0��&._�d��I����cʝ��6m�:��n:k�)��6�T����;ۉ}��ߪPi�g	���1.�hY�E�4\5&�ү���A��� �����ެ��� f��_�tc�X�L��$�Zј3K��`+զ~<gpŘ�s�D���B%�	�\��E[j���yV�;�-����ո!���;H�رM\�Z�`��oT�oU��w�A�����5g6��ψ�U;}���Xl)�W�'���U�1 ���?��6�%f^���ZA�����I�=V��o�ɪ(�W=��ŶNs�+6�?��?B�9�%�(5�Ya� �QW�����k�˃Ia��;"7y|��),;�����׊@e6n�d�������T��n4�`pM���Ou9O�I?���A/��m��}�Ī1D�dng��U"���4�om�)��M��P�j�z�����>�ھ�0R8k>�gSc{��'����*�>������0���~9���1#��v��,& ism�����|[��^���)g�,���8�*x?�<�*�r�b�㤚����6��{<��� �m�{��c��=s�a��u���F�Es�clwF�	�4f\DP�5X�<�<��k����o���Խ���;�	�d�{r�!�̉T�N�����W�4�I�����Ru�S����\+?"����#<�\���W���	K	�̾�Cn���Wª_H{r*�ȝq@�D}3}'��q�8��l5�>���g]T�?N�k��i �vnU�����;��$�`=�y�.֒�H��j��R�\�!*#Jx1������8!�������u�潑�$4ܗ�t�
g�$���)�?&G����+Lu#��İh��?��S/!��[��u�j��w�ӎ���0ʅI��x�(�/+:�WV�9$�S;�&M���S��o�����NvC�F8�+�N�w���>����l�Af�15�8���6�؞�9�{��5������uL���~;]^;��/Z��[��+H�5�S�,��=F+X���n����� �(��#�e����[jn�|����<��6��l��D��vlu������>����!7m��D�&�-TђU�W0]�g�P��3��S>G�'m��t~�G����):�aIð'��_<���6�����Aӭ�2�ȏ(��ˍ��;�Rh�� `l������#�>mC��p�i�a��]*���f�	�֛q�Zf�����O�jSd��!1��к&d6�����Ā]F�#��g�����
#�L�~�ǿ��aqX�����%��2|%�.Lc�^�f�(Ìɚ����5���'O8��.Ǿg�	��,1��g�[��}�uY�<A;_Ql�5��:ʿ���$vd�g�yq�4A?�:JԔ����B���we�7��!}q϶���d�l���+O�Nh^Bt�O�+� +������` ����{y۱=��v����0�6��?f��������W���SeqH�%����/V��m�
�ۢ�5�$��[H�����
�.[;۷��`C]�֨��������7�*�MUB"�:yXo���f6�"zO��3ĸo��Ϭ�/����w�TH�)�d���wՓ�7��=hC3�I�썅7��ɤ�1x@@�%��pr�]k� ��o���Ҭ��!�1��6����4��z��ֻ�^:/�FD��
i��&�avׯ�a�jj�$��>z�'C����yudjCFo���M�}�#^��
�1{ߌ�RBRt�G�����4��M�Ak
4���w��g���j���W���$�V�qC*mV��وX����F4y�XgH������2���X����](L�'2 �X���Nf��㙎{����뚞�6��g�
M^�1?��OR���5aq� ����1����2#���xP(K�a�:�ߓ�����V���U�iSR)�Z�G�s,2>��a���}�Z�E5�ڎ���.%|Z!�G�`�%,~�N"fF����G�h������;nf&I�qzj`<�b��zY�9.�U��:�e�cq���`���~�O�H�N���(~nf��K�����L}�~_�fu�B�1������@��UTZ\<�*^��,ީ�à�2�j�q��pt��=�'ߤ#��E?�sE4�QRbc��G�����i_sV��JCv��{�p�;$�&!sg4|L��L���n����m�}�0��ILo�bJ�EF��Q�$���j�ļ�����/�C�jbQ`N���Y/*��Y����nv6ӄ�ch��N@�RNf��og�ڭw�.�bE�F��Z��YZ*'3�"b����FiD�8����� _T8��{o\Ć!S�k~e*�v��'�?i�f�tr�&H����m��R���n(�
]�߃�n�B��(�)�,xV�Ǉ�]}n �=�g�|zf���Ө�w����� ��p �C��:
�.}����U��%1��Mǿ����/�5}>L����P8>D�����'���(A��V�T��T+̡'��h���;�3/$���Q���/�6\���1���ePbnD7�ۗ�($�@���m��b�����N�;w�bd����((�8;���ۦπ�f�q��8_&3o���ED��d������w��NF�1�2�	�U.����p�3���p�v��c{�3��Zw�x\W^���#*�K��9:���H�up��=>A��1�ø5K�LF�����?\�ռG�\~&8�������Ps�2ʎ�64j�pX��db�pB���q�����͵�{#�G�p��_')������H��qI'R�����]�u`2�t�n:�f�E���������B�C���֐)!�r���j���t �s�u�p��q��s���)����������%k���A��QZZ\�3�}Գ�"ii�|yl���C_iCy�Y��� �#���P
|�e�z�
�����V��b�8���%W�e��i�.����� �˪ ��fbZqۂp���8���h=��$�Q�b{���L`��Sƹs6��`�+:�EE��J=P)≼:'���ߖY��;�W���e&h�)�D���J&_�W��|�+{��*?T{�Ci�Im�G�����c�������v:��7������+�X�l�~,����[z��`��>�t$���g@ ��0����*�%R�>_�@@3�x��W���U	=q�H�z��]�3ԝ�cE�$��`K�	��I�!ף�SMֽ�v7�;��ˎ�o�j�[(E�Q�l�w���#��+�Yl��s�(!%��P������{��X��2L{'ʛ�l}\��-q=��}���٘j��Q�-�@�b��9��_���h��m��s����:*��I(J�g���������E|���H�J�������"llM��04p���L�^�r�\%sx��H����L]1/�R�ck,#��.�Rp���?k������P|�~A� 	����2y�*y���w)�Γ7a��i~���>��Wv^\�&_\bR���cj�>�s��1v݄�w����W�.+�����!=�Ca�ﱣ�O��q��f<��M$�G�eM`�bj\�65�{G�!||���p�� K��)Zǆ�6Ȓ-xD8��:��8AнnWR�?�h�_��ڈ���[�����t�3,�}O'��j:�G������2��f�6zW���0��:76oA$5�w�-e�q�P˯:�7�MIޤ��6�D!�� ����L�#u�%�3n�L9ED�w%[���7��t$�-մ�^�`e��xMNB�6���*p{�4��BMy� ��	X��RZF���&.�e�YZ\=A��4��R&�*��*���~Ĩ�D�FZ����L�	I�L�؋Y��J�3��P�#hr=C?L���*�pZ�Ǿ6O-^�`��Zo0�>XB����#Вu�J ���|��~�F�3v�D�ߙj�}���P\�v�j(�L<n���k	n���@���H���\��\e8�>e�~�/��5�_�j���7���`!`2\�+s�R�;΀�Ge"!����~�Klx����uQ�G�I��Pq���j�����!۴��Pq?��&��S0l����i���&�"�6�|�Z�kԮ�H�&CY� Uda���Օb���B[�ʐP����XA�i���=�B�����
�^\����74�L���,����)<6�_� �ו���䳾�I:L-v.��#�jic�Hd���{��:���2u��D79�B�PR��#����@TS�	�l��G��.-5�������~XJ�{�R
"��ܺϗ�c�W�-����M��-�l?�ş��Q�'S�J1���b�ؤ��n#�Jh�F�Q1�ܧ�guub��G9L�X�J2���$�G�<N��d�a`�Pϕ�����o���Um�Y�h��\�<Y�B8���d2�ۺ',����g�����󋁥���Ԥ��>Џ�a��o8�)$+�����9�w����� � G�;8�Ԝ��b�b����K�j��½-�}85�&A��8�t�>7����r�^��S�Pn��0�L�T������~���:G�o��e�U����6E��=�S��1�x�����G�-��k�/H���n���]2r���:^Zq�i�m��Ի�.Y�������
�LX���������vd���l`�x=�â���3�\TB"��
�q-�M�ьaUn��o�m��O�ƀlb/�����56c".'ua(�v��q��Q�'ǩm�I��(3�z+P�y׮ci��Sh�z��u`ε�i�R-����*��~�F]CU3`�,���槙$w&��B)<�t���<Y�q���W�R�ʆ㐍����'�¹z�X�.��κ�Ư���uD
[�NH]@�s�h��j������[���t�4��x�2��~X�]��0j#��"�*Y�b�����U[�f	�Uv.C�>�F�X��׭!�'RO{zґ�1��/i�Z�v�p��P)����%���5'd_�?b��_�ߵ���p�fM|�����V�8r8_	t~���w���;C=���0��wBh�*:���ut>��ۓV34E��xK���Y�F0�W��ƞ��I���)5�����Lh#�ȫSvl��`<(��иu�r
d_� �p���ܹ5�W{
�@s4�56��ʴ]�`�hڨ�����W�aQ������������S����
+���0�'�B��[����j3����Ӏ�n��k��we�d<����ċ�����O��As3���?�!�N>N��,���=��ZI{�����g���������S��F!��l4��#�u#*�_l�3��ZLnJ�p�0y�4��1�e��K!�i�j��9h#ؓ���U'���[I�9�D����Ө(fᑌpA�aH<kP}ى��l�UU���kUFF�r8�f�!˗2�MH�����@	��趼S�+T�es"fP/RZztÀ�����+��*��(Sن�h\���3�7p�P7�2���X�N�w�5�G�%��^=G�+�"*��m�y��R��u�6�k�D´�E�x�>���dps@|H�0�;���**�0�I��a
�Y���ⱷ��rL�ҡ.sME�됺_�O�l� ����ه旅dZ�6��M��}+�ꋉ߫0��ڈ�~�C���>��T����e'v'c&y����LmeG�c���	��d���""ɜ9�A�{� �m;��!k~+=\;�E>
�?��$jLN�����4l�٪X�FJ0O��(��g�!����'IO��鹷�:�)�K������H/�i[���s:D��^W�W�;@-������o2� 9�!��$�ʁ�����ķ�����@��3SA8/mU�$����w�t��7�h�u��֢���P��3J��>Y�`!I�ʳ�zZJ~!�����
.����&Qz��"D����蚟K���J�xB\9ɗ��D]�Ǭ�tEq:�r��G�������IVb�����Ax�{KaW�p�ٯۻ똺���ƈ��(���g���Є� BN�w@��m�DW�L<�S����9ɫ�޾��L箐-$����\�� ���\�*k�nLӵ�$O,ves����pA#
MYwM=�������h����!AvlI�?�<mR\��Yڧ��ʏ"�#LϿ�Ȅe�-�W{5��$�:�@['-��E:���Nd��Z�Bgݸݰ`  �˼��S�<�P��Е�0���;�R��e�-�1Q61�4�~!��̄�On�v�Y�אf����2$�sYpПv�#��A�� Q��Gz�
D����]Ng 9j��J�	�� �~9���P����"*=�J���!���ߍ���%<�HڞC���ɽ�fM{�8"X�T��5B��T58�a"{�O�����[�ϋ4�ӈ� u����yj��!LU�#,�΁�L�V�t�g��(��?�՛z��-����"��?�4Q7�$�b��mf�f�M~����au7��C屖�+%v� �L�'���lK�����r�TGe� ~ȉ2`oֈ����(6������EEf��%y��`��C�:�y���c��eh=�<ú�P|���16����ԟF|̚�h�7J���!]%�X��O�(-а��8m��d���k���k�F���ԍU��( h�KJ_\*�d�Iw8mH�g��6<����۠��ס�3\1%�b�X��iSB�V,��|$�m7�۸݅[ |1k�NfG�~��Äͦ�~!<�AL�i�W�Օ��@5�K��9�auZ��&�wc���b�
�ijW䥼���2��/�����/�'��ˡ��v�(����0/B�l�<=��-���	|r��Kg��4(�6�ѷ/�4�|��@��D�a��p����m+���Y����D�:���^c����~9���~?���7�`U5�th��[E-k	�]�D����'m'�'N�DK�Y�&�^L1�*Z��Rِ�5܆1橭U`���^�"�H��H�b�V<5�.;R�>��fۢ� �VʀbKf��/��1dlH0nB� ���i ��)����b��8_\��sS)�N��]�*f�co��-&��7!���)a��:9g������r�f�׾�F�����g�3O
�]��Z\���7����Ќ�h�ڸ�h����-& ?	ejG�W�:>�jFS_��d�n؆��TIe@o�^a�������l�.�dGD��7,8-��X ��3�&����[n����"
�J=�|{�Ԧ�:3��Q��qmR��àb#m�6�D���~p�dL���n/�7�����?�o�#Ha�t7�b>�!�*�4CRͱz�"�މp�����^�:a�z8�=:���Z(�&�zo�#g�=讫`���{��o>�S�m���A�?<Q����d�CbNř�๥21����^^�9��@������Ó($�_����B��Ʋ��#��g�Ì�/�x��ɀ�8:����QZ��݆����$����3Ꝅ*�`V�0��^�	�h6��M������������Y�n�3��r��Ԁ�1f�8����N���+���$��-�9�ѿ!���%���,s���t��̝(j���5�~�}ߢ��t��=5B�H�t�x���0�u�|f��+�T.R�=	Q�^<ԨL�n�����	�t����/���XGz�y����pnbN5�Z�HtM:�������l}�(���&�2��f�=  ��B�FB{�-���|��R\Ӊ�M�/Hx"�P~dwgL�uqMJn������|�,v�с�&C¯����z_�_���DhI��}�<�l:� BI�M �S�E�|���U�ٜ+�������i�D�A5�5���5>��8�,�������ݜ���`d�A�q/@���-��$����z���Jd1�_�M!P�$�Ig-���cb@���q���6��?��P���o@�yc�Si�pٱr��u����x��"�����[���w��.��t������@��S~̒SB�;mS�oڇ�/3�޽I����X �Z�i��n��[��_߿���C��zh������<NV��;zT �&�5U\ �p�A�q���1�z��F9NV�/�����}�?��Mb2�[ �>&��N�/�����9��G��s�0���
���]-:[}g� ����Ҳ ���(�N+O&)��(w�����q45;�1Z�X��0�@����_������$��ns=8�s��V�1\�Rk�\0sv�ʑ(�6֖D�U����(���o�ez�~3��]팹�-����{���ri��ۍ��p:i*He����Q=�Z_2H��s k��Go6�2�䌙�������:�.(̃�#V�	O���k5$b�|�)kR���yw{��Y��P�ze�}�Kn������.Œy��v\-��45_L^U���[@v4����Z�J�7GW���N�?���3���7�b!f�0M��
7֦V���\'8�z��V%\k#�
��(�a|��Ũ�5�Z��ذY��r;�[q+��xD$R���Hq$bO>�	�3�`?0��[I#���PBx������^�������R �*�hp%	uǥ��lV�Cr���V/	\�'p����-���":@��c�'�*5/����*\�X�쐖�_7&|�{V�;^\	�/��M������#u�4��sF��i����!(&���f£��칈RQg�r��H�E����R��I-�3� �7K�%e�:��A���`�D�o�����Y��}�}��͉j�����Ӈ���]ぢk~�3��/z�A2��?�j�Y7��������ǒH�W����7U�/���jy��V
S��DM��tan���a᠒�Lyd��i-����.�x��\lȖ�r��ƒi��r~�˱��k:W����l&wL��>��S�{/6����6x2��~�)�����z�?�z����mR��C��WxO��/�dE�~̳*��K@�"�υ!ZA�[gi����*T��zv�*�x �|V�t�?c��6&�kctɵW������Q�����ݕy��hJrg�a���zd�����3H�Dhc�5�ja-�~�>(�=��|�0#O�mP@Z��UX�SPρ��@��R��p<o��?�X�s�6�x���9wo�݀��M	M�â��3��EJd����
%d�LO��J�s���6���3�0;?����a籁�����L�f�VP3MM�ӎ��Dc^�Q?NR	-�,�`��v( ���R����7�ͷ��m
�sI���G0Tl�R�?!�YJ��0{���*��㻀�Q�,sg���9��']ӻt�-\��#�y���H��d���o���"w�z=��ׄ�;	�q�3}��ű� 1\�_"�4519~�!� #�*���:�G<m��i��)��it�����U",.��gԟ�@w�����&O�v�&��p/܌�~׆�bpOz|�r�g�ND$���TZ�g���.)���2��O�r��O�>[VYY��ɗ����=�0'2��O��WË�.��o���F ��<���ީ�ĥj���}1��'p7��@w2~&2���1H��,�WA�O���d���HM��K:^�b�	*F"��,����s��Ou�;:*G��Ѽ�	J'C�j��}XC��J���q �G�]�yLB@��>Hg�#���S��5��	�3E��n�� ^�ʒh��*�� ��� )i��~�āf�Ā���D|��K뚃L���q� ����bRg��6�K�m5� ��[���$)�ď�c�}�����L9b����)��w#e���p�Z$N�̡��ib�JS�{-M�Og<gv����Ԏ���}��G/V�t̨�E�8���;���l~qNo�P* J(��[f��F���b���¢��t��m@��x~��5@�8 Y�^�~~s:�#����k�U��zqN4�ܴ�
/�k��h��??���h�?J�kؓN�M*hÿvr�f/% #2M&�Q;�u�|0��w�'Y�>L��En}�l/�ǌ�4�ߣ���<p�V��z�CNE�
X�]D8�)Mu�I&�
T=�OpjL*�]9�lx�0�c����6Ex�c0��LA,B���ˡi�.��I�'�YS���a�c&R�p�k��v�U�8�ų��r!g�E((��Ź��mz��k.o��b��ʚ�h�;��U�OL$W|H/S�D:���1!J���Jv�P����/!9����D�g�n�(ufGH�l����� ��;��[8gk����tE����W(<��(�!�K���Ǔ��~���|H�Oς� Qe�R�]���7[��@c��N~=����;��ˎs2������$X�s�6[��[����8����Fn����/�U�����1�C������虱D�O�΁�G����g�H���X�\&�Q7jz�Ȕ1����oh%4����T�1,#�P�C�kb�/(��ͪ/���?�4n��J��jΟ)|����A,�p9?(<&S��U���r���Ǎk��$ۈ]l
�'#^h8-s�J��
=K ���h�ŝV�јU��Ã�6 �"��%�s]��<��4����ߤs ��ͺ�x��q�6EL��T���r�U)�81t�q��$����ǜ�(�&g0G=����rQ�%3�⊝�[W�:_MЯ�nRj5?�VxOk`G?{���?���t�U��."��cϤ��S��!z��:�t���#�A��~|1&�b7�bg����Q�s7z�2�@�Dvl��S�C��������`p8�/����eV@�"J�Ո�l�]�}Z9!�}����Hc�O\](�(B^�0�r�n�����$6����f��CnP���5Η�.�����XEZ�Z��#������o^�J�}�U��	�'�U��������*�7E⥡�Ā�@K�W�'���V���q�zI�G���X"r#��{$M?�^Z������8��ޕÆ�R��C��9�bz�B���������*�紉>��0ic	�U��16ev��39�����쐣۲G��*�I��X�ϨI�����r_��	R��������b�j3��
�a�e��8
�\�;���ަȭ9i��Ծ�JnoDn/���~-�-���패#��@�Ek�:�D�GX+����"�v
����WM嗤n��|�;>5�1%{`��.��aB
���.I� D�z�-Py_��x����/j������*dtT��_(j}	k�W��X�&V]C�]���zU�GB���W�H�e����{��S$?�6(3�X:��D@HC��>u�:�7��&�u�	��@q�8+|�t��X)�Y�4k�~�PQo�='.ĭ(�׉L��p��+����tޯG� snI�+*�Xt{�t )���xWI�}Zž�v��C�5�hO�lG��dғV�l�6�/x�E+p��:q@���
����=����!�6�����o@c7U��e6p�b�r�>Ө������\�~P]x���SB��FqU�3]�ӌ>3g��P>��)�7��b>*����љy�Z�`��fx'�����J¢H�7f)�������f�-��Y�=C�hu����0&���B�C���T��<�G�'����?��]��x��*RC޿
�@eS��,+�,�:>�N��"����f.X�Q�;�Y����d��Hcŗ�WU�}=1 rV�A��Hk��*+a%��������ٸ��`�U�>�ݗ��}���u*S�zbV�&�U忌%��gV��D���#��)�K|m ٖ����N]id�������{=á�Y˩l(X���8>��;�3�u>��1�h�����AM@�cA�Bf�nIPn�2a�T��yo ����U^�ǂ��2hp���8�`)�����pM1�{�-0��,fw����MZmTp����՘O�h#Ɍ�㽴3��r��"�F_.�R�j��ܝ߬�M��yc����������.ooY�����Ƙ�]����.���cT�}�}9ج�r�K���h�8-Qa1?��vHv['֙��Z���`��S#7<�N�f	�4���~���u/Av����t�@LO�f� -9~ ,PW�B�����J+ �C��Qe.ɊJKJ�;`���5�:��6s�-`���J��i�,��Y�4����;�ߏ�����o��pm0do�;�ɶ��_&�]��g[8V��"�p�<���d-�&t4Lhq}�me�U�!d�� ����UH�o�L"X*΃�E7�Ee�$%�G�
D[�h�t�r���V,�gꔔ'D�L�M�W����B�Bl�J�jv��;��ͺw>'b�zk����/��(�|U����D�4却O�tٹ��Z��6TW
><󢝊����˛��I��ܴ��}�C�A��l7BqNt���,��NF��d�j�i�m�)~�w�5��'z�,�HrEZ?0�4���}X
���&K.� �B_Q����K4~�$__2x��x��,�{���+͍y��m��,����¶:>ٟ�2>f�1"���q��+ƙmt�����FR3����u�Tﰾ�OtI�	'����vfׁR��N2.�p؏�������h��p\s@I��v͘�Z+So	ɭ0�bD���R���o_�P?c���{0���v��Z3q|pq�]��T��4˘�Ei_��;t�B%�����nA��(�ER<��`�	%兕F�]��k��=Wp!�+� Q�7B}��1�b�n���!�{�z�������U��^���F��m\����?K�:�����ƅ'��ƥb,ڹQɧ��uQ�c�\�l��ǖ�u|*b�4�Dd�Vl��k~�T_-C
��suJ�����@2�ۃM��in�͈2��~�Y��P���SO����gI�٤�+����]�2���3tch{�x�4�$G#�'L L�h�U���7�7/e;�:��M�h'*�����A�gS��_2a#ٲōz�J���Ơs��ׁ�7[r^}(�e	�p��\����[�DM���kW+~�(B�T	��l��C~�Dfi&�� ��X&��+��������Y���>qO����.���-�x���7M!NҢ�W�O��������4��qzԄ�0xA�V�p��[_HA6-v[6�_�RJ�@�?�?�9W�]7��X0�bt�8lũ��Ƞ'�ߗϜI���B(�>_i��t��{�x�t������A�lɱYf��Vx�'"�7��э�//�	*�N\_�{M���ڣR�&9��Nxa���=/+������$��ݦ%��|~��ٚA�+�Cu\*�{�H^����'sXN�����kb���.��5N��8_��)�N�}@}e����i\	��-"af�������$]�axv$�b_ٖ��̵�yeNh�!�N��P���pG+�F��*x{�����a[��\���K�(��k@�⮌C��5�ʸ
���a���:� ��(�w���H�L�کi�%��4��~�vw R��F1�ߪ����?5��������vD	'�(
I��An���4�g&��̃��k�rѣ�t���X��ٺ��%����Ͻ�J�����WY;���]�R�fy�����d��@)�]��4Dw�� �����5�P�_u���N0��:%��o�	�=��_�*�^%&�Ǧ���o�M^��j���jq�t�>sV-^N~Ȣ�C�h �_&�4�1d5q:��k񛻰�vzu�#ԸG�{��Ʊr<r��^_e�����:p�ߵ���,#��),��J";�aЮ61�D����t�B]��E��УMn�d�����������!;�K�6$� ��O���xs���]�ݑ��V��Pm�?Q��\o���I٤�s=	���	�f��$٫�;�c����i�ER��hwڄh�Cr:_��@�2��=v;���ZO-�����?j;�d}p�/4��{�(�.�.]�����TJ�r6�:���>����C��B�L�;5C���&a�1�� �a��`�$��TQD?�}
�z�
>~z��e���"�	��ڊ��K�hTz�C�/��B쉝�����O]S�F �B���@2Kn�?��\+�'eN>�F�@ț,�*���e:ƥoC�Q4)0�t?���� ����Ŭ�z<�;��W㊢N�E7��nZv��A���"�B�;�v��'%����M���=���Ώ��H|��+���G�H��ŉ�(�o�5+����.ݛ�ފ�M���1�7=��F�8n^���M�P�������i%�3�q��G��:� ���?�ɐ,�9!�ܡ�e��v����w���u�]�M�i9[� :�|3�|���6:�<����)�� ZO��!�o�F��ُ��Su��I�T�`p'�t��A%�pD!_�-]�r���4l����X�Xڊ������j���y'�Xa�i7�k?(R m(��F�J�Z�lh�%�d�A�`f��B�+�M�ro���ST�����o]�YCYX��	�����AvV��D��i>&NNJϐ���E���Luh�Ȱ������1�PE#�c��	~j��6���X̗t��b�Y��܅�i�w��7��ґ��`2�`1���N�{���yg1��r�Lq$�)`r2�Z���y�ϩ{?�W������7�o�	�C|��SPCk�����:��W��j�(���\�)�!^e�����=�~�M��$�����Va�LIx�����X/���f�?m.��A��~��U������̼w:�?]=�̸uK��Fa�)w��u/�m���o��\m^�cWI�8#��AI��n�VE�L�vʐ��m�����v5/�!Pw�7E�������W��eDCؚ+�TZ�@���9����p��.O�o<A�>F�cށsaO�u�*�S�ې:It�Ё���:���Ό�"H$ີ1rx˲����"�����M��$q�&��㞯O����h~���r%��ږ�#[&���;Ϭ-���jDY�OJHla�S�~^]
}tWГ������^�adaW5���)%h����!�_��W�?%E��\��w���aHa��3������(�wߘR��u�TS=���2�'Ϗ^*s�P��H�І�`y�)���B�#�G��D�t��niBS����n(5x��d8�PQ�EaBش��ذ`Y�G�=���U��q��Td�Qˑ����v 5fD������
,�>�CD��dYǅ?����|����@����X;d͌��R��AW���;���D�w9Tc��q��1P�$�����!��u�"����M�onv4&̎"?׌�1BʨT�ڥ>��H\�?	#���87R�8U$�P(H�=���!c������� �b�����5������_ފOz��� �'j�O�B�|�K�Y@�`�L�H�X�,�gY������۵�+I�ኝ����=L��&��_F��>��,΢�kn,�!,jd)�%F�bi��FS�!�|ѷr�=���^���tО��?�l`���`��?gkI�E�S�t/�*�b�M� ������P���J箓_���K�43��<�i��B3���@X�[C�@fme|%~�	��/��	��Mof�g�S#$�l@J���� �a�.�	C��>4@<���׾n�F/}���{��N�@����0i�0��|}�f\��,��J�#p_ Oyd���*ٹi>�:�9���C*3	��Z7H�}�&.-[8|���j�d]��	�=_60b-{I�G���n�Nxv CU��R��R;d�7	�rf鼃�E1~�aC�3îk�t~g$;�9�sN
�� ���%�'���4�%��J���t� �������5�jؘ�6���_w�p6v�Ӝ~~�)Rj��:(�gWl]��R`�j-��îݗ���EP��oJX�);e�WR��A�	����c��i�w�Ǎ)�la��������>|�蝡���O��q��}V=-�R)z	ܢ��Y�/ �_5��\9�����S�Gãd��r��f�𖎄�x��P�f�T������pe��3�:���`����y�6��~զ��a��d��)���)������F}{���	�h�)��w��\���7�� `�d�n��Ө���ryU����*1��*�iU���Q���d�R�>�9�x�RC> V齶o�sX�C[����b4�H<9�f���MM��)'ֈ$��̰�[!��Ou	�fG�Y`M*F���H��ňvQa�d�0o-���ë�:�U���$sOJ����1��K�)��ݮ�^ȍ �Y��!L l�V���O�z��G��!*}��
0�g]�4�D��qNg��-���p@bވj[	�)�������'��q�d�#�-h��Q��(\�-=�:�ŭ	Dh��NC�w4A��P��0�؛\�!#J�]>�݃H�ZKkO;�����Z�"����{^߯�NF<�9��=k��F4�K�$����M���-�	{!l�>�����О�8ܭ:o�a_��ց�
h˿8��*a�[��n����i:#�ʞ�X�Eֆ�1�� ��@�e����ꔑ$\��H�ڨ��af�*R�M��/أz�c ��ׅ��*�jc��98��*�Y���S#.2�2NF,�^������&����O�Ƽ�g7t,��E�^�s�O* �7U�o��*x9Yp��-I�/��T�g��+��3.E�������Ә
�g�62 cf�{�s��:t���m�Uc�Ih2r���1"�]gylb�9�WfR�'Y�]���%bzm�=��ke��6eBU��1�#���N4�yȣ�1����(����]fk�?N���y]�<jsmq]����Ka:�e�	q�'Io���_��ǂ�C��&R�k�TY�Cz�O��O��F�.�'��iO��Y�
n���1u�}�Tmo+)_���
���+��;���ş�
c���_ۈdp�����hc+=/�{����8lif�5G;h�\�<��W����<�p���&}�����r�W)��Qpf�Z��I7J��m����ׂ�?��x�Y�Ei�ī;%y$`�۲�V}!iG*	#v:�e��M.��fK��t9X�I�?�20Vf�ΐ]g�6�{k�[waL�c"���.�	����W;�0�Sd��P���j��L/��株���F�ј7V{l��m ,�3)����5�e�μ�O�J*��7J��t�<��]��T!J6��@����f .�KZ�x�0�-�o�P☃���Xb��sV��i�r��x(Q��Qmτ����q��ҽ���8��U��H[e�ALp���7�o���7��Sb�ñ�2�-��m���u`��!vj���z���K�u~�S��&�3K���H�׳*�u�W0��S��ӿS�(�i�C�$�7�m�t}�,�o$1]�n�{���DG��|,��!;P��)��\M�9������(�Y����:��1�U#�t)G �������{�Y���o-W`��F��P_h ťޥ�a����s�	Xo�:O�o���ŗ���ܡ�mY�(�4CJ�$k���T�o�?%`|��	u�R���:I�4����"权�ڪ���^���yg(��\�O�K�w|p��J���K�>��R�_'M�2^�0b	��N|�x��:9�$�%��`�~1z�B�Y�����@L�h)�6���zm�M�AK���׊�Ah^�I��M���:���dXdt��/d�����Ͻ@���p�0�}RU)}���(RRg�^L0�͆psa�����p�"VVH��M��@v�4�3O2�� 7�^K��~"�|VZ�^k���I�=��$p|<���<�7x���)�`}�*A��yʉ
���Q Ѳr�[	�)Y"p�4@}��p��/e�)�/�Y�+���}�����{�4����-��6��IxA�}��"�>B�<���y��[j�e�8�2��\��K[����W���j��"�����8��R;�ˁM����� �$�	�Z\$��}�X�T�����J=Y��^>a���w2K"`{�5���v��ul�d�!�l�[��r��=8���q+���os03����A�' ��Ѩ/�|@%p= ��o�1E��W�Az���AJR±�_8��{cĳi�cG}+�!�B��E�l�kW�����]4��~%(�F��cm����{��5/*�C���G��D�!,�|�K�b���ļ]�d"J-]�����s�RI��f_��y�Չ�9����}�Y@�a�ɬ�b����@d;�2�< ��dЖ�LrD�Q���~L�`0S� ��z#�z�23��
~x>�(Ƴ�ˀ�2J_C���J�1�67*��ZY�
ё�����F"l]���-�=q�A��w��-�� VH���@V���2Z:̅��?$-?�v���K�O1�@�yC G��$1[2}�)���a�6^� w��e CHC#��r�:K����3��)�Z�a�AʣP/�S,� �kˮ/��h�(pOz��!�wN4�"^Z-2�*�vD�	������[w�����0�����2��[W����]P����`�6��)��P=�E��g9�x}�Я08SO#Zb���gXO��.15	�A���V	o�#,��M:�����D��8
E3��}��%�!҆�H��V&�st�pp�*=��{q�%.���ޕ��M��e%�Y���H�:e�jlKMH��ׇ���
h�ع���"p���hk�[r��q}�[���G�ܩ=��!ED����J�^L}��uR.a9�}�D�]���bdq��c���|��k׬7�*����sn����7c�ų��x	�WR��̃�v��Wb9`R�y��&}�Nӑ{"Y�2xWn�گ�%HI�%���\�����N��cH�**RF��/�c����A���gI<I�%�|7e��*=�c����)��V_������'~��j�#[����"E�����oCiS��Ag�u"dNUl�*? ����F

�a26/D���r����.�mN�҆�ܱ9���
��IR�� ���%�c�g<�|:��EP3����*��	ݤ�^ች�k�.}���]dy�uv�F�����"T�h���9
�v+���[�gZM��nJZ?�cfc�մ��;��h�?�����$�>���/���)Q���b�$��SȦ�� �d}�R�y]kixD�<��nl,Cz�_�$��;�ӛl�� ]�^߭e�H���د~�N�T&�EB�\�~�O�<�tm<@@Oq�1����n-��.a���j�	2k�5`ml��w43E>�Q���uqMXP��5(�+J������"nT�?�J�B"��JTmHG9ȍ����`!�a�?�����_�^��-(x<b��.�G���8`Vǐes�-�,ǣ� >X����U�<���E]��#�~�w���P��A���_GT-Z�Ӷ��L8dpu�m�
�����Je�	<�7U0۲�yK����V����od�F��;�<��y�����Q	ۉo��ROE�2�JF�W',�bF����`��~\�c��V\�E#�8)��Fգ�Kb�[���:jb��]��(6Ƙ7)S���Z�@>�� ����g�Ccm`V���7���4�k��x�j���g7����B�c���F`/��#���#B�'б}��@��:!�0�n�6������JйS+^z3������=���aڂG���P�*�^�!�����M*.���P�.s����.�U�"L�?��e6����e���� �GR������~j!(�W��e�� �����%E��<.����w��]DSۻ�*��6a��)��ݹ����zH)hV��RA����<��$L?|Z����)��oyS���cu�a��e�}��
����
P�c����ၴ.�����5���fQY�*��8�-D���hzT���B�����`1��YHEz2%+k鿖��s��t=�Vn�|�W������E,�H�Cm�e�&"�L��lh�܊ �#ŭ��=���]���|�XS=Xugw"��H�qd9�?ڶ����X�Ԟu�ldwP�$ǈz{>�o�\PfK�|�z��2�+�fE'h���!�%�R�pC�
/y��\!���g��� �.#ql���8O�.�}��1�)�ӀT���̐�\��5!���0(Ч*����+Vw��?q�x�����J�^�l��~0蘛��Y��'��91���V��L�*¶�J�̌{d=��>��~"F>~���d�ǔ�d�	��R�	�/�~	�����Z6�#B�"���/��)1?H�\���a� �}ѥy�B�����j��i��p��D�����SF�¾�Hb>:��^�cs�wQ?/3��Z�b��`�� ���a�6���$�Ý��K�I3w7�S4~g�ʋ ��꠪�âB�2ᯄ_�QP��+c�6��E�mt�$ܘ,���T��":�pM�#8�^�?�J��xZ������gh�7 aYe'zogt6J3E�91	��<p�-���'�û�YH�E�N%M(:7���� �+�D��/'�@�:V\[6Lt�C���
��A��'�j����KE4�l��k��o�"s9ߟ��#G�4�	�����GH̏�0�nZ1�e���%}�ѶUZV�b�Y��*_!������f$J��	%���YP:>��f�.�,���|=@���dJOd���r �@g��?䢊��v�)�xtqZ�?�0i(w"4"1؈� ��\P�5�\!�k&�|i����΀�����\���BϞ����� ���Yש},�"��b;!�[��G�A.��T�8mۢՎ��oܝ�+�,�u�J)`�Y�ٽ���L�-F)`@�R���A�,?h[�Daa����~��
Z)���g�*��	w�5��`�����'!xM��)�&������WWRw;�c����6�!��\���<rb�|��{,�hq��[/uu	���z��]= Q�J�(��X�}qx�zL�U���<�M�c$�0��^;?ۆ~T������x�tO��u tR� pV+R��m'q� Z.��=X7Ū-W�h9�ٲzk��مaf!H��^ ���[�g�Үz6 ����Igy�h���S[�٩*昣���˓\+a��Nze5#�cK~	�����s�ϡ� 9����w"��׭e|m{ĩ(���Iሦ�s=�a�2�
�2A����ʲa_d%>b��a�5�{������� x,���־�Q�^�QaP�%5�[y3>�rb8ߖ𺸆0�INwY*@Q���e�.G��',&́v�ĈH����ؑZ�QJ�*���n~�N��:a�_?9n�ر��4��kX-kt1�W'#����BK[Uu��]0�`!����ҝ_h��H,�-��-��WI$^p�b�%Fg@��j�ѕڧ�	ZŻ1S�@��&���V)>����VG��n���.c:�dc�s���+��+ybM�u��ݷ=`8rkoTDp�ͰkF�`����{��w�j)�dv��3?����˭$'���JFU����7�lu��Q�^,AӲ4���;�|2/���b��B��]�dZ��\���|��2x�±Ɏ��t�1���{��Z�@�S�?��O6�y0pGar�Q�����-+�jd�O*�F�7�P�� r֟M��
wx��	2�?���6�V�̤�^�d�V���@�Y�cx���F^'�de�����ЁD�i�f��B��u��h����,�'FA_��SiT2V%�g�*Ć۠Ɉ�/A�n�.��9��zG�r>��M4x
�DB
m�=k� e�+-�����%a욮/-6X$	�)��i:��gT.%�Q��]�w�/Q��>�����)}#*V�	��lCή�҂��>U*۸
C�rEnA|H���!�(QP�
��g;N���� Wk���AߤVɴ�@�Ǜ*W���]1����i˓��V����'�T9t�Ct�h*�RiG�`f�����,��)�7��q�� ����,<n�n[F=1N����;F��א��s�ͮ��A�O&�e���&�-Y��ц����Ѽ�b@K�l�:ݪ��Pv����l�����q��V嗍1�������:Jkl������ƸzMԆLu��g���KP"#�\'*��pXE��-�B������ٖ��̦=H<0PK�o��ġAw�oT;J�wˁ=Է蚫	ثDJ<gWI����rdn����Ss(�E�\�,�#'�I�O?������q���O߳dz(>���,�t�[�PF|��8�Ĵ�k
*�%��-w}��@`����|���:J9�1�O	C�v���5E*M�7�)J����A��(8�� 	K�yZwNQ[Nq�^�Z���/3K�b�G'���c�Q��n��%�@�&*ԁ�w[���@M�dFm���47��.[����F��_��6���]�K*�seBg���Y1�(����f�l��ݺ�"~��A�?��瑗c�r�#�>�r�,@d����"Sa��d�삕�M�/�.K��~�8x�m|um�$�l����ۿ��=l` �_���HTQZ��t'G�a����[����E߳���3v[{����u׃(y'��+	'0z�s�����M�o�m�-%��.�cE����~'G>d����L)�3������� ��6�46�R�%�JH��A3��ː�����՚N�̷.��zn�Q�U�HtN�sqe�g�w�6wkZ�6���S��~�K�w�	 D���2<M�/?-�����@W{�TPԉ�O*Gba92x��N9��ހ��i�6�nK.4�L0)]��)��N�e���R81f�2t3`�A�x8>*�+U�C;v$ԙ�Y@��Г
~�0zw;��k��v��^#�;T�T�g^��G6�\#�1�!ܷ��Ie��7`J�w�h� �p��%����_sk��rdJ4�0��\g4�>�:�;Hl���.��ҏ_�C�}�
}i�"`�b��]�:�2����	�z�J�T� u�*M�_�'*��(��$�ߪ��x6#l����ʛ�*�C�y��dE���L�Di�ǀg���hEM�O�I#B�7���.Rca��3��P���k4��w�@�|e�6Q��I
ai�᳒}Pf�t���q}������^�����,-[�ۓ�Ʉ�6%�8�L�:��>�c��@�Ǉ烇=$+� J���f��G����C�u���ΏuC����/���:D�JWګ��3|�Ӽǚ�#�� jfY�<,���u����r������%��G0��L�IK�u��EQY����<D�զe~���c��*l�yOQZ	�Bw�B�K-.۵KzR�\�Ontz'����<��%�䮒�!�>��b�F�%^�|�߉��.4c-z�o<"�y�Ѻ��`Z`����;�QVv��c�E��FleQzC�4�u�������8�d,�]�Oa�R����ui+��0]Yu;Ie7$9hj-�:�V�D���_	=�:��lPg��^���^͋r[��'��fؠ��X�=9(x,9(�U�����˙��/�D��|R��>��@-�3��Đ�a3�_�E�nm��Jq� �F��zSL��\w�9�b� ��N�M7kA�^xG��⡐(7�( ��{B�����Z�Ȭ9���کH�b�l2st+G"G ����a�]���e(��<���k�KM�� ��9x��e��>h�i�f۠Z�>�7�GA�A�߆3�i�^���w�.�U-�O�'$�\����J	o�<}�G�4�^���Ԃ)���1P&�hi _Q8���A�I�Tf}��m�x�'��]��K�ߑ
���~p�����ަ;�9��N�m�n��KZ�������4Y�c�D��:Kd#~��g��
��pZ�!E��ɘ�kp��*g�<�AB� @)�'���_��
��\ˡ0��y��MM5|e��N0]��m��؇#à���f���3pָ��;m$��{a|�Zl��]��q�Q�R�uF�~�z��������y��^���95�d�YEXt��.^�������%�G�?1��>]�$e?���6V�'��4��1�??��VI���U�`��6X"�*1t��RǛ��&�@���ⱛ
^�Ea�#)��#ł�-[J#{7�W���C.��m���KG�u���r?��c|�2K�r��ɩ�t��ˊ?u.Lໝ|���NM�VV�v�=R���+G�u��m�&���aW׊��E��R�l�mZ�?V��	�6E����&�5��W���Coe���cY���#gI#P��9 ����67�#&��yEK^�=ie��@�j�e�lFE�|-q��e�8d�xLC<(C��\��;�S(nn���u�o�,����������II��z����E ��^,��Ys��2�$�|G�Ny���"_�$�;��m1�$�����(�w�[?'�U� �����\���2�� �EM?.���<@u��=̡+�T!���:�Wƙ{jy6Ӣ�.d�zC+p�&5�5!�Jԝ���Q�G�1�)��u�D9��3G]�\
��J{�`�?��D�҃��$��G��OX�2F1����{�x��J�I����5xi��4Y�%3gp��i0�!
ϔ��U6����I����&q����o�8!S���tMĔ:Giz��pZ,���%���qh�~ڡ)�HӐKV{m{D88{%�!~�5? ' a�N��Ƞ�/�&K?�,$NFK����*Ż8���R����>� YZ�Yh�0��}�~Y�5l�du��=�M�V@��I*y�M��7���^���!#��5l6ֲ'��}2='K8ؐ��������DWO��-���q�}��bh���rf:ܥ��8ޢ��#Q�r��R��I ��~�$���u��s'�0;��J��O���fp��X3�$�K�2�LM�#�x�oM1��p�(�Z�7��5�-2L��AŵI�E)�i> ,�[g�?\m�����cŘW3J��{j�W[�����Z�j9�/;��/�G�U������d,�3�ii-^�c�c�n+���Jg�*�#z�!�X7�-���T,�R�Ł|?���+����
S޲���y�@�3P(����Qj�Ms��𱚔�v5Ԃ[��$��)�!�C���]~:�h��ιh���|3����c>7e��u>�^� =� �<!=0,��`������q3_"�� ���k�B�ǲڙ���G�H�ʢ��g�c4<�9]���ǃ���M�0�9�Q�^,���,�H��L���*����7�q�����٢�E]�ܙ�h��m�pC�X��È�>���B8Ńk���/7��V����ǂR�����e�/@r�،�Az�]�ot��X�������^r!´j�� �t���h��P��u�.(�!IH#���>M`��G��6�7�!�ؙC$��a�u�����]�]L�=s`�>��[�^��u �����b�f��ށ�����u2�<w���������ȏ������D�D��I�5��7��7z�E���XQ�͚?w�e!?����Y�A�t�$��g2�����t�53��gE� �齽�	���6_�h�Oׂ��D��1���<l5x�-�"6��/
�/0"��#���q�Zu]�E�&�9�K#>��9e2�������$=w�! 󼀟g���1}��[�Oqbf�P��@���[b�u��i�NЀ���fx�K�#	��xy���p�rf_�5�&4PV���?�㡱�p�+��2�Y�eA�!�j�(2��
��%Tc�l�`����w��
�-��ev"�^y�W�}��dN� e]��^�L�����Ĩ��SM���ӭvt��Dua�_hS��c��#�Z1�"����W�5��!�l�ĆHV�2[Q�!��w�}R�v������W;k�L�j�H{#�~|��Ħ�7>�g3�#T�
���\ ��h��*L�����C�e�OSB����Lbo�'�.�`��ws��%>kh�}�w�	�h���M�D��m>IK�t�Y)��Ρ������Y#�U��D�B��~z3ؼ����7�o0����E��W[ �|�����!į�22G��P��z[҇�<5��&�d7�K? \3�����V6���Iw ��P�ñ��r�{�bl�) 7��<�Ϝ}��c���x����k���E��I9���6�_A�1��ʑ�/lk�o-˨Cn{t9?��eЏ���1���$]g髙�^!f�M~�wz��M��jq����-�IO���@ ؉�ҍ<V�Ő�=6�
\���1�����?2�厖T�����=���(Q0#dj�ClN��d��^01�u�]����}A�"e�MP����`���<ꑚ&)Y��2������m�%�,rC�x�D7��L�l?��-���aL?ˣK�eF]���M)�ͬ�(8��KbU��+�K}�E{�a	���ٷu��ӯ�M�jHV�ĕl��M��$�z,������l��1S��(|0�뒥0�x��F���c�f��@cSR֘�ɩm��'@��-}_�l�/{��[ԣ�kl�c7a�:7D!�E2�����z]�s￭1"�M��"�i-�}T��ÔÃ�r��ך��������b?]CƯ�Lw�-ٯa��.�F��hC��BBJ�XY�!:ǳX��x�'gI�q<�Ѫ�p�k5��1����\lVb��Žq�FX�Ƕ���mH�޼T.���%H�/�o\Z�'�b:+e�4r]�哞���G�8#�.d5R�Ht�(�oUW.:�oЩ�F� �	�,~k_3���9�8���tH��@paq�q����̂ZWr�[YGJ���^�!�|�Nf��eH�����LJ���?�0�	k�3��Vr*��_:���j!�:{[��K�d�yv�hEf�γ@��y��ⱟ�>r ��ꃌ�&���ǉU���E�f*]��՘���xG�x#�j��FΣ��6��@�j�^Pdq�ƙ�ҟ���+"�#J�C
˽@_e�؜)���'�aĩ� U�?bT�^Q�a�����sf5�̽Tk�aۘ�.9�yj�c�����. l��4.�� ��5���kp@ި�_ <��w�qP�Y��������7�����~��'@����Ġ��TqwT�ű�v�"�j�V���d��	��H-��6�k���ć��N<�+���;�T��@��H"��V;��?�}�o�^�	b�ӥ������]	Ͻ�P�����-)%�A㈾X#l����ݤ��Aw�`�Y�=��������Z���E_����䰚a0��Bl�\;�^��	$e�̛�V"�p/+K��,�3FuG�X�m[�^i�ERl�$(���F�k�gs�	�|��kg�Y�ԧ���zƛ�А���ŃT��ju�'���9p2EL�/G��Q,,VEDO��F��k�T�
	�3�eh��!k�1u�N������d�?�ZV����)�z�0�)5�O�+�yY�4�����0`h;�+��.�J��e�hBρ�f`{�4���1� s�o��D�+�|=Rt6����r�e�>#�M�AX�WOؤ�i��_�i�6����Rѵ��}�o�@��M�����!�O����bt�X-!�_���+"�fʡ�bA[�%<GڝюA����L[���{S�SK@2ʨB����v �uu1���ى7��5��JJ���=�;6��w/���v�|3I>ոΣ<%[u��9*��r��N��0M`"�ٮɰkX�9) ,t�$Ӟ���r�ĺCk���>��Y�b�B���:��W�0]���` ���W�\r�����|7k�ݮ��.s<��M�S�X��T�J��\�]�|f�r/�`=�(�W�L�3�3��DA ��D8kT�Ε��(���ڕ:D���9c���d���v�B#�9.�A�#*�^�!����'����2�u�0@����Mޯe��<�x�z���r+��$q,|9�4��%��tW��]K<�ǚ����y�00�o��q��;gT��|�rl=����+)�e�� �U�AU���_����~�h6�p����WL8߇������${�ק_8<J��\��Z���q{r�6�Nm��x��x�(У���o��v�<�t�m����C���K�ϸ�K�� DF��nyyZ��;� �p�uBJ�k}Dt"?�6��Z�
�X���.2��sm��Gzһ�/#[`������!�����Lc�n��]�._/q���������}VM�w�ag�r������Ƕ�\�mKX�:.�M� =H����"r��N���.@�E�!�P�1�Lj-ٰ�U]�f�����;}����tB�2K+/������4��ܠ<7��P�s�PZq8���\�.}R���bv��P���$ۖ
��=G]VN`���/)Vѓ��٨Wu�_S��F�'-lǝ��e�?�؂�=<0�Z>��h�.�+�_+ρn��{0G���M�?����7ګ��/W{JF( �g�]�>V���r2�i<�#Ҋo�be�]S9�T��3&�SOB"�L��!ڍ��&���u���27o��$�!^nR ��0�,��ܸ���>7r�;���=�V�,�����eU!6��65$���p���1L�)�;�X޻-	"I_��
�0͟ᨮ�w��޳�����ǃy�!M}�6d>�Q��p�I�H�@ҭ��S����.��`��i@���x���k��h��
�䵥F�j��KT�S0,���G��$�@�𜤵���� G:�D�;�<���Aj��Z=��cg��?��7+Z�X��%��Ko4:�ո�'��]	�Е�ſ/_���h4s��ғ��)�4o���M�UƊ2�z���=ݢ��U~>�?���V7�s�1F�\��;R�j59kE�Ig��>N�(��4ϙ�΁�^�#�ɦ��i�%����	��'{�|q�<��u�t`2�r�� ~v��Д�A��~� ���P/꿨DեS�rP�܌��Z��h>�c~����������y�X`G(��A�����0����Ȓ��G���9#�L��j���>Լ�?LC>�\�vw�T��Î��� �h�����*>Wc� �1�=�,ڶ���5cN�\? r[m7^d�w| �e�lwJ;�&�'��I3n{���4#^BRc0��,�?mG�we�e�4���x�<��q��J ~�LH��2y@P�b�=gp�ݚ�w���)����ŞFn�V��A.F�`$��N��0?	�Yco1�����6�e"e�}/���	�n����X��FK�H���<�ҶZ�ۮk�i��p�kq�����0)�>��ٮF��L�#��atK�8JYu��B�R�
�M�a�D.mX �D��3�y0���/�GH�8� }Ƒ��ˀd� �E��`�G�YjߠfX��BJMa��Q6e�7�au���f�y��?ς�n�����]� �$\G����|��w�|�I��y�d �qz�p�,��ۤ��`/��{A�����l�ԘI!�$?8�^VX�����+�u�@����] ��2CW��4����O�p�rMѱ�D��?���k��y��Q�}���z��$�C�>�$L��xQ���X�D�<=���F�{줉��NAb��a�3b��z����tBh-� S~�uT�w<ҹ0��1��8��l�ю��Tط��и&mJ�R���{(Ԕ��ޥO���Sd7QZ9]�-�� ���|��
I�x���.��Z��/SM����|���ڨ��V��"i2i[��6�YU�"�J����Sm-�����|�D�@9 �	5�ǧ=:峓)�a~_ܰh7�c\�/�~�����RfP��t�_K{�=)1y��i��I5��s�Ґ0�P���N�A��8]C!�EZ�%.Xj�StO�	���<�<�S2x�E=P2
�[]�N##��-�,&7,A�=�������[�>��13#	�+�&��ͥ�{��@U�,�U�j�f4/Y]�Zoh�qi�I<��d�����c+'Q���b������^d�U�T��
_�t*�B�C*��NHO�q4�S9Aф��UE���"�t�_����(���=kG�'��=G/���s�4/�6؍Q0Ip�6���� �}Ǝ��S���*ա��K�h�P��џ�O�a��_�䆡 s���7v��f�{OuwQ���(*۠���fW4��**���V����}��L���c֦�\?�|c��w�Å*!C|��r9	u�`	
ٺ�詸=� �����U��:��9�\D�D.;V9��M(z|E)|��ꘅ�CcxV��7�c����r`�2D)?�������|��A�N�E���Fd�y��������)����"�J���g�EE>ap�����,,�� e���G1f��2���d�hk�|�{|����`d�ti ��ʃ���j����^~�����,�+���`�h�	��֭a��(�q*�Я�9�W�0�S&�9���o��wO��"_�펰�r��1+���mBW�:~����a����o��v�/��((7��-�;Թ���(3OT��"L-P}m+�,����ۏy4��C=�-9ٓ'��JS��D�U�%-�)t��+[��+�}�;�hu�2��c�C�ݭÙg�J�����C2��K񨤱8?R��+[�&��aΐ��9��!�r3���� TV �h��M}CD�|���a��r`۳�?A�_���l���N��]	��P|�P���x�uٜk��.�^d,�X��=�
{�U����4�����X��wj�c��N��#%����'t��RbQ�D��7v�'� 0��s�8��'N�3�qӳ�����8U#�),#�[p�@K�>�6�=�S�](˪c�2.x!��Z ���qH�Ta�&�j�'=��S֡�0?��k���r�3�'a��Uo���w�{n1�����S9ZO |�`K��/>G�	���T�d>w�\� X�g�K�V&-%*��t��x�t�
�1�>�����t�ә��3l�u�1 �w�T�j��-��>�U�h��S)���T@���eA��8����`�)_��j�x�sΜ`]ێ#�w�k%�L�l�xX���Z�5A��^� �~|5)�>��#oyP6��_�:&��p�rT�E�p�Ԍ��n�4�����ʷy���1��\���L+/e{EaY>��q����QU"^��+��\Nau��M=f�Abv��+|��E���lU��k;-��@/�� CT~��ƋwȜ���I���Y�v���3z	:�i��ߍ�}�E���v�S���H��Ɠ���`Ɓ���HGP�J���F�HO��c�p�2K,�\�#.e��.	h�fӕ�F�kI�-\e���y������`�u�����~�?118�E�n�*'9�#h�[K�F���m���C*����f������wU�r�HL|a�cɴ}�+~���"rX�����h�m�jٳ�S��u/��٧ͼ��+�T��' b���#��o;�'Z~#�mGF�yӬ;1`i ����Ή�L6)ۖ�#�w�%��ͳ!��.m� }6nã���kj�<$�ڨk�tY��v���KZ���ˢA�8NG��1M�j���A�n�9�Ҭ���lv5u�'r��,���ͫ�tR�p��w���~v�eT�X��c�Q�"}��Ĳg�uЩRy,ʇeP���w|꩒�ӡ�D�HL��
X�� H*�W�ǐ��RG
���H(t�~��o 4}��t��)h�u�Ju��e�F|�n���2����c��͞y�o�*Z�[b�V��m���/(P{�O
pX��pI�R���6\��PE�����0��׸EA")�q��M��.�FK�~�K	�t��E�C��v�'�曌�Inq�+%
�rj�QG�b蚳��K��8|RsK9��`n&�zOV�/hD*�kͩC1G�>��(�/}���ZL�w�b��[�}h/#��Q$Hg��W�GG���}!S���[�V@�u��x<N�hOqKk�P�nw:�6����p������_��de�DE�W�� �"�9N7�c�Orܼ����?��Y*�e��������X��v���`��0�a���&��k �[i����T�����W�ח�^.���X����6��k� ��g��~�Z�8�Jҟl�T
ǫ�0ys��f�уY����,��nD�����/��_�LnW
�:��	W������d�s��5)W*�����øh�g7�0�eTb�u_$������1��ŧȷ�B\&d��7m�1�a6@���<s���wd>
HUV�uku�I4�਽ԚA�Be��L��f4hLؽ�I)���h�է#�?�ٵ��?@���@EJ��D�U�����i���򅉙�2f�/p~?-�{�
�eXS
���륤K�ۻ�簩wL�r��PjB�y�4��ׄM�}�&ujm���ɭrպ�c���uZf*[�mhx��,wb{�!��C���ǭhFn5L����_�]4*�4{DF)����^�G[�8�!G)p�p�F����|�9�)���vMR�툚.����|�'��zِGCP�ҵ$#�ز$
�����k�BV!�����[M����w��:=�nls	w�W=���y��2=�ͮL¢ϊ��;j���e�l]P�ixP$�N�	+O��ʻ��C�\�@�ζ��hsM&7��,f��~c�&��;����}�F��o����,� ����C+[���~�l��Hʆ�C}o�=zT��t1�����	@+?�������,k`M��l�߽�� �E�E�a��I��eE[�J�1!�0uf<:�y��A�)L�Br���1q���o�[\HW("[wUl֟9�l�6e�:�o����)��y���.�Z��"=�����KA�,���T��hDeȸ/�/	g������y9�۔#WI!�\��1��ҾQ�\�Q��2[�D��C����;4��B!p���j���͹�P���2ɬ�mPq�wZ��Ǵ3����Vz���
΃����#�i�-�B�_�O&��귭�@J
7x�Rpu�9L���"C��]�y�19�B���
l��؜��!!�ķ�X"���7�y�Y�(5��r��#!(�ю�H�1�������L�R��%yU���J�26�2N�p��@"Ŀ5|����d'7U�����O��N���*KၨF]�2Q�G�� ^��ĺ&]�e������pvx2� �� pj�|x��bӶ�n!e�&p�}7%�,iVÂ�iUd�� ���I1�TM�w2��+��JLvGۋq7�x�=�%���&L�SX}��*6�Q�d�5B#U����0�(ʿ����c��]��յ��>�-'ǣ�8e����_�LF☗o���R��L0k�������͂���u5�ɞg��v����y���{?#DET/�[�ͣ��2>�:�I�LB�xt����!��
.C��Ǡ�ϑt����/�v`6����څ>���3H@B��(�u���2���|@��b���Nr��ƙT�5��f��$���u_V
n�����;�+��8����/ŸZڑ��Aگ�uՖ�~f�>��Вt�F07�\���"�H���ˈ�X����*���aٛ��vr�A-�u��DDC��7��ǝm�(���~��X���h�!���X�%�E����6��?IKI��?,�+�>#�����3d����<↘m��@���?wȠ�q[�P� 3N�6�Om�50�����<��g{K�^?����\Ή��3h%�$��4<�J�����������Q��`0���L9��u��2S��Z6c �Vi'�K�8P��>��q�'e1i��1۹�ӗ^�0
����}�\/�h1d:^b��$�	��'GE@˺��3T=���g�R�.6R�sc#?�,�+~�dX����}{Ê���(f��`y�DWD��x2��I��^5� p�9�����zh3��Q* ���h���qwG����*6뭉cވ� k�&mU�52c�2ӿ,�4?ѷ�!���PA\�!��-6��2Y���o�����n�KJ����==ǉժ�'��w�֕��P���-��e��v������JG� ��`{4B2�v��k�R�cM4&���=�C�/�FRv��N���|E��	�#�Q�f��s҃��y6O���$׈�i��TDh�]9݀sE���!��j�)뵥Iwα��E)6�i ��3.O����P��h[�ٚa�d��2Fu�$D�vr�t�̞ip<u�]oٌ�>�p����91g�^d�F�4i�SZA`���w�|ZJeK�q7����aS:��|���6���pKT��~e��YJ���+�}I�dj80>|�A�H��hF(�Bh�j:]s!�v��8E3b��uR��c� ���e�= O�n}��
I��Z�N
�d� 0�w��]2Le�>���U�=��j����+��Շl��d�i���:�{=D� DW�j#9��	67�Qg��b�vTR�� �ې��N��3+�F���fe�eR���@���Us�Y�1��Z(`ΠO$��2�!��=@Bf�v�kL��t˦/-t}����8���J��$�;�Z�h���Kw��`�Qט�X���C�����I&�r�T�0΅3�� �T�E��@���;9���*:@x:���P��c?
E��xw�bOd��7]���O�����r���w-��+�Ϣw$R~z��W�ݍ��2�;q��TgɎ)6,�j�u�`_�	���9��*������Dy���Ar�4�a�5Ӎ�';��$xcA���fH~(ƣ�5]�ۏش��h{Q#�?y�����Tn�&���[A�'�+���JT�S��je� ?��ʲbX�~k���2�yHF0��ݶ��0�>�dσӎ�͠pKc5U���T�3����q_�������/Iu�'t�nஶepյ�����~�*O����*�A��,"��#��Z�[�a�z3�2��j���oud$��yP2����}�N��:b�m������qi�X�oմn���k�M���+6���AS���(sF�r<�7#��wyqӱS�o"�Q`��IH|��A����1��O�G��tcDT�{EW��n��nqV�49��KH��v�R��C��N&P]��]ۿ2�B���O&�m+'Q��W<�^�\�V�I-�Δ*��p�;qC�t��8�C}&ep�B`ll u�Jk�Q%�[�8W�<����/t1���b�Ç�,��}�@ �>��:�{x���ƪW?���7�kv�P�e++C���~�`ڦ��5fee'�pMn�KNi9*��;�dU�f\�s�T�i�sb%A��_݃����v-�B�}�&P`�uj�+���n_��b�ɢl �f�����l��T��'�AP�t��F�@�2�C�:�(1v�'x.�"��u�V���"��I�iM]Yd�����w���X�i�`�A���㓡T��.C�4v�2�� D=Ke���U��%zK�7�)R��T
;οtR�m�D�MG�u>"~���%[N�Ln)�)άu=�)w�w�Q�������O��a;?���KX�����-��%ɵޙ�#���ln���'����7�(��{�1�um-P���>_�!��C�<�|��ĕŅ��_��i��!��`��F6	��KMξ0��
��`����x�z��,:LeH�T`��I��ʒ��w=0���<i�e_��=Ȣ�y*N�ʂ�8�}����0�9e^�Л继~��@/�J�R'�b��[M�^�-V��f �+hh^�E�+�.�25�����u�q|9�M[���l�;�v7�Q��Ƈ۰B<��y{m�4e,j>�A�$H�$<
�V��jOs~>�<�u�]��$Qꛄ����ȗ��ə������N,S�L&��[��*Zl��f�������a?tZ��>=�L�&�r8���L8X �D���8��v�\n&1�ia%���k���i��i"P2���[U?S_6��y�ն�f��0p����]eo�6�aT��=����)W_1�dL6Ε���������xc�I�ty-��Vh��z��~B=w����L1�@�y���J ���k����yb��n!�����*��cPf���r�����Ƿ^�h{Re����b�\�d� j��z���hF
s4O�w��o�}9�����}v�����P���_-�6�ΰ��5J>��x�]r?�	Ѫ�G��Ļ�Ě�"��M����N΃ްU�r���U2���� �L�&�v��eS=�~*� �3�a^C(6��B�96�+��J?��շ��9�Pr�9^j��
�Ap�f��������%L"���%���c�`��>SA��>�p=7�9��yq�-`��r�;�u)M�v�P��YAIo@)��מ�H1��`�/�e<j]�H*�(퇣*j�e��.P�����]�T��w���šӜ�k罐)��f�
�!D{��1 �:�F�L2���}&.��ѹ(�eCH�r����Ԑ�]�j��a5��'K�*��O8N1�QPiZh�h��i8���l���w'����UzƸ����ԓIK6Tȗ&iq�6�i@M�֣�����`�ٿ�S�_�eN��^c�Z��Q��	0�q!W��9�4��.�eS�{�N������&7�ʴ�v ܮ��m���JY��r�u^Bظk�H�g+)�8�H��Yo7�<(b�+j�J��fP����f��T];Ɣ|Pܩ�����co6�;i��J�qr��Mg�Ua�����EKޜ_�e����U���c7�����GH;_R�(�ꗵ�'���L)���ݏ��+���8�V30d6�5�F8W�-�,)�s)\쟙늦J� 2�ƿ<�\ FP�O�E�|� ����*�0��x��MԎ�^�ZЬ��Wd5�D�*˵���>IW�_����&T�����^KcG̷]��W��A�݀Z�j�YX,\��_����[EiZ�F�F�s�v�u�n���q�l�N�cO����>B֩#�<ͅ)	^䐵c��^�g�u��+�R_�V!+�Z
8a�|���e����Ǚ������.8�`ٮȫBy�g2��RS�ya|E8Ĭ���d����ss#/�}���.r�ë6��5�ػ8ل~U-'�+��u����aIz��p��3�ы�r������9�E�|���|�(�A�4�QM �qI����<��,-��
���Ľ^9���ǿ�@G��r�t���%�$����.`������*h�c4��U�X�c�̼��f��z��^G�ǹ��/u\��C���!���&]���7$�D�� V
D����$���He&)Z2�G��ڊ
��;?����w|���v�gS	>Η�5��B���g8���h�n������K`4��z������نk�����r�����-%	ފ*7�
V�A d=�'qO�S^ok0�T�a���\������V���/�_b��Ǟ�������ӕ@k�Gu�c(ll��/w�dϖ;,��ի~D��q�8��TF� @�<�����?imD%6Nq$ܽF��	�ҍ�+c:�x��eU#�]� �L_����Ab� �=��aE���%~a(1��,[Kj����M�y�$��+�o�v �!fђd���'����>��{��tt�^>�"�g�~��f�v�n��+���r7��yx��m�^Ɔ������YQ�9�
�e�'&y�mr�~{���L ��w��8��_%��9�)O�n|�Ϧݼ�T�Y:q�'@��V&JA��-��+@�iw3��)�/o�p���j��C�,h�lvy���x��*%����Tw����P?9h^�pǇ��B+�0���<�]�8�әi�N�,����veJg�!F�W�*�������CzPh���|�O��L�����*A�8����	&>Nu���,PH��>3Z�fRk����v��-��&�J�%s]¼\��B�Ҭi*���ЕZ	G)�n�=��hz���;��%�d?hcnTg�L�v���^#�H�
�����'��*-�<��[���R����F�ܮPiyb��j��T�'�]� �y���ml�ဿ&�wC�:�{�,����G)�����^4��X D}�Y�R}7>�Ǔ�Xw��CL-SlT��;�`@�>Z��M�ov��������8�9��k�QfR�VE g��`����T�6���2ن8��r�G�s��>fנ؊�]PUp��w�ePu�-�p!����슂�e�ibd��-=�86�,��{X)Z���0�(�=��O*��E{3VЋ2��Ua����P�4l���)bf|���~�;\�6?ǘ;� O��o�~� ~`���~��brh�%���L�m�f��ŝ�FZ»%�,r O�YS��%��PP)���q@+]AB����6�D$NA��J�m],�0�5�:u ��+fЋ\yF��5$H�;|�$o��N����a��4ŵ��{�~t��_d����)���Q�螭�qV3��V��-E z�GRt3�gsD4X�؏�J�dq����;B�K�^O�٭x���%�-�θ�w)�:��9/sҞF5���D]�2�]��R<���g'3+��K̀ԇ0I�@�Wc�8r����Umr��FV�w�\��!���Ȗ��*���E�������E7	�����ŒRj�%&��Z��.o~(@��w)Y�νK 0�x��Ӥ�����b�x���p�����~�O:Ƣ�Rg%URL�f���"-Q�V��M�񲨌����$V+r����)`���r�R*]X�����T�?�O�Ĝ�в��E/�2�����)��v�r㫑�Muz��\�0�oY=��R�"@�Q�%��z-���;&��`����R?�@L���-?~�� �J<���z�c.�e�2�ں� zn�U��]��:���d��:t�|[yJ�ϋ�MVmw���ѧg[��p,���8��Xv�C�CϞ�wm
*˯!+M�~h�#��I�Y�#k�0$V<p�Jcc9~�_��kM�)떽C?Z��X��PMT�7-&١۝�ǄK�=_I���ץ�s��Э���n��HV���'�*G�໸�p��4D�Aƣ�z��q�r%y�sV�/������H[ȍ�O�|k�� ����91L~e���������[�E�K�L�soj��h���V=f͇FO���24^�\i���Ý���d��F�m�Uy�d��L�&����F��`�lROvf�U�0b�N���5��]u"���Ib��s�"'�]SIA=�N"|,{'�3��y�j(�b;5�"��tIxŊu�}.J��k�'B��P�!���/%��Q�v����so�`������8��!���4��Z-�y3~v@|�z�AȔm�
SXi4���ޝ���]s��Ⱦ�������7����ӻ
�A�k2����G�['�7�"T��g4^c��er�AF�x�k7�o���{I��^k��%���=h���a@�|>{�H%œ�#K���[������'��U�{b,�^h���ic��?L��#�����������2�_�\��:@���Z�7 ���Jrz��J_�y���j&���C TE
Vͮ|�R�)͏]ӧ5�3��,ܛN ?�p�i�7�AXTH�1��dܑծBR��Fvc����6�t�-j?B�9�P�Ѵkɯ��S�䂒b�0J� Up��x�<�/x.��$8��IG_�8�6��PX�1�ݢ"֡g�	,��t>�{�����qT��^ @�ۀ������T�v�7ؑ�`n�O'��r��b �EG"b�k߉�b1�&5����3>+C�����e��V��ݽ5na">I`�Q\�
Q,������ާ����\�E�8���X����<�i_+x�4��4�\m"��߃R��:+A0�?8����(�b҂0>�@�ָ���[l�E���,N;�*7t	*9o���&�4(���w�U�ԝ���d_�db��G��E��#'�$���ơ�+&�k��Qd���Z�S$M�@�� ����i����5=�{K�Ԕ'g���'R�����Z�o!@��DG@ �:��ӭ9���4���vH��N}~��?0�g���$�+�Sh|O�&5o�e+&=⹹�A�sS.�uTsE����hdu��`9`�Q�,F��7 V�nc���c�3�p��#���]��0��d�������?���{f��p��/��2gЩ����<��T�}'�lъ/��/��m��\�)��9��c�	�>C� bt�1�����>w���k���B�`� ���!9wo\�"/^@j��j�K����El�3"��������f߈�;%�2Z���{O:�����O�!�5�u��S��n�>���h�sz�DUAZ�o�b��6&U?0�c[C�P���H�Qi� A%;��u�������N�i�4j�7���?�	\4�6�ih}���_}	�7�<��<�C]��l���f�\:\��<uu~)��I����ud90�2�@���W(�-L��.Z�a�����I�&5
*��1�1@&��u�WFۯ)2�'���d���WS@�(��J<0 ��H1��oþ�Kb�zĜ��fmJlh<�����2K.�9{�+W�FK�������N����|-�Um�Q��u�\ʒ��mvp3��7�g�&��%�4�{��hE�l ?������X�+N�c�r���a��&��A:
�������Us莩�}����b!z�A;�Pi���Ѱ/eR��+;��-
}���`�������b���r�Ǧ�e�H�ZÏ�(.�~��ڎ5���"��`�bD`Ä����Qp}>����פn�_��\9���͒�^�`��v�����)��r4��*�ެ��5��j�� wv����X�G��;:���m�J��F�(�k�y�G�_-�*�sX?}'�S���$ ���m�tͥ��E 1˻�]�z;�"�������,ώ�������~:��6f�h][��Xױ�IO��u�� �
	]a����� �AI�*f�z��$�����g,@��6=G��Uu�ZR-k�� gkY�+<�ւ�:7!e�jO}TM���Тy�spM�H�қ���:z�.�z��ʻaЁ��`s;��:^eo�� ���_�沵��NMcchsp&oT5"��Ty�ly�{��mq�ӳ���΅7�@ƾ
����[��fc��q�x��o�ʿ@=����P{��$��e{�q�M�͖�i�^�
�V28UJ�I=�4��n��_��qk2[UR�v�C�V�Z�Z�@%�@�\�T���M�5R�Y�(�G�<:���+ E
�*՜y�X���L�UЉ��Aw�vɪ B�G}��a����G���x���稘|�)[�z^hGĿ�)��R�郛�������-f@
]�"�N�P��s-��/�>���_�^^��}����m�m˙��zD(Nꑌ�N6Q�e� �u$�׾���vN�cs#z~�٢8�*��fZ��@��O��L�(�u��,�{@lS���\22�����w2���+F�xp�Uc�u���k�۬����3�� �;�|e��:��#��N�X����
��:�P�+�����>k��bU[ch� @����w��N-Jh\�^̆N9���g�p�(˕��YO�0�#a�fZAB��O)���>�(�4�T/}[jv|�]����	���ѵ��6ed>���lU^n���Z�����!���f�����W�4��I6��:G����x(d��Yl����������0�ۆ��5?Niɱ��K��"B�{���5������`�^��bBV�(�=Ǐ�ӕ|��i�F��M��d04&h_��g#pQ�bI��K�b��\�ɨN*�4n�	^�x��qk�j{���4Z������z�!�Ɍ11����=:<)�����|�ٚwA�\z���.�d����EK�5�u����9)~���r2
���2q�V�bS���&��Z4��9k�6c�Dc��-�+D���CnQ�e��9/}�,�ޓ�G=���Ug%U�8�!��_wXç����.�X0���� ��f�ؕ�7TR~�w��!vJ���CH�X�q3��X�E�Տ�º	���%�3�Zn�^�`��6w��K���uw�}���	*r.������_�5G˾�q�Q��B��@ � �}7��1�(���Ho��ⵋ��fej�|	*_~����j�qS_����[�D�x��
��FT��0����=��������a�Рz��))���.�!�8� UEk�Π(|ɳ$�YK;�M�UpǸ�IgS��_�_Mg:�s����X���y����݀dW�󄟣� ���U�P��?�mvqra�
`�,�Wj�ҭ��ZU�t�����C�FD���z�h|hi1Bv�SF���\wB�m��P2BV�1k�{��(�a_���P���b�q�j��SM�Z�O���[��0�8�zj;gk��2���?�lf�	ϝT"��C��eH�Ωw�=�����<ͬY�Pc�0^��eovƐ&�"������s,
ө�Ima+h�&s%=���J͓ˡ�^.��	%J�ռ�<�g�/РC��ꚷK��,�#"���O�_H��I�L�1N9�UO�&�ۿ���������>˩�8#c��+��@g2@�Q�=���{�;�p~��r� @�=��
���!N�G����\-���P{!z��ń���0�hOG��������iG|��'�$���.!�0��%�)�P��w5��M��)�R,��0�2�G�Av����6�C��$�6�����N؏\���pϷ�o=�iW-ڿ���)��H�%r��C��sWW�Nk�h;cuf�G��;�<2����B8#��SzP��M�碞�H��?��!=9��V|��I-�Fj�-�S Q|k�o���#�c��K�&��'��Wu�_���EoR�L{���ΜeƐ�����nq*���X�L�P��E-�g���cH�2cOץ��$Ԯ�f4i�^�	#Ǻ���5����C��������C�c}T~���'�X6�Udhy�,��{�����BO�9����9HN5�*XY��V�b��o�+��Жj�'=��63�j��~>�Hs����W�(���B�F��縓����GB~]?b�x�װi�F��fɢq7"F����=�M3��wewP`Ym�~�i�L����t�l�X-���tZ�/C!Ձ�h����
�$���&98�#�DP8�׼��.�aE�� 7�{��������z�܋Su�ɷ��J4�ԅK���]z��++n5v�����aI�/p���l�(��s�dl��r�l���ۭg\H�e�HC����gr�`;E��0�1���#>{��ۜjo��KÍ���sd!��<듞K�\E9%Z?^��t�{�PT�Y�+x�f�*?�&��e	�O� O#���~����9����0�Ȁ�EC�z� ?7N����C{`]tŅji��S� 1R�.F��F�~O�ǀ�{��-e桲�g�п�����B<Xo��W;I�F�&��3m!Sڇk���?{���!ZO�����'�<
yS�-)��9�*f��o��Q���Tt��|�<�!h�L�d�*����ª�H��,Ps�2�L�w�������D�����h�gU~/��c�L��j�4K����llص��(��N-O"�9�lu������p�BJ}��,YC3s�,�uy^A�V���y�i�9\�ņM``_��DRB�
~~� Hm**�H��f�x0=��{��8�b��WX]���>��?"�)�kt�ܒ�q;��"�vn�#Gd��G���~Gb���r��R�.���P��{����o�\]X���.����4n����z��8�aY�%Z�C��7F?��(����F�����wVތU�=Xj�v!�=�L���}��w:0��^.�F��QX1���}�ԇeB�^�j��68�֮!:��fL&�Q90�6�{�� ?�X(͋Q\�0���f��p�I��9�d�պ��)q8���>�v����ʒ��-~����
"F��!CBz
.)�s^�0HvN�������j����6}��� �c޹6��M6�Q���A�����%�L���J��ֺ���%3�9�Tw��k�;B{����N��$�4KJT;�\��\CT�`�7�{�-ē���2����BҒN�9��u�P.�`�\����`�Ǔ�����E4���D��veI^ ��o�U��\`DP����&��* �m?i�m^Fu��}`��"� u1��K;�K��C'wH|�H���Iz?xF�����34DhjDi�!�N��c!�0�{P�.��Յ �Z��.اޠ�����Y�{�^�ҿŔ��Ĩ9|<|�:4���w
�g�Ų���>�Y.5�¬ro+PJ��Zk+{�	� z� 1��0���X�W��c��g;�#wxK��]J����5V48&Q�qU&٣('ߐ�l�8Y����\���Sxx�b<�N���������>�"ʾ�{!6��H��y��6�=۟�F�}�~Z�U�+��d1/���c6&6��ghե j)1p0T�'IU=dWD�S��3靀���L��!h��B�hp��[�nGi��1"�b���w��Z�dzc��ڶ^�m;fH[>�<���}�q���BlD�Ջ>���1��eQ���F���&���C���3:���З�m�JS<�mP��6&�zk�hl�F����xx3�U㏈AE�*�=;��#����!�y.�5~�mp���6tKZ���}uĩ���b��1������â�19����~!����|z�~_\�&�#�$�h
B'��#HGOӬ��o���f�&�iyD́�'��4ISc��[�����#���i=�Yk���ޗ�v"�N>ɐ@�8<VfLòT{D��p��T��l�^C �<DL}Oo��퍼����tq�jTٓa�ݓ�m]�ڲ�/����4��Wk	*b�"G�G��A����PRÎ���%�ۃh7�s�􄜹���H��H ��i��H�nZ<I3a�rZ�X�D�QE�M&*�D
���$y>�������+�޿hJ����KeZ
�Fz�}�����=�1��`�\�(9�2BI�I�&)�0i6�����I'���W2�6�:���f�����d��X%��x�Ń�
�:%�+�u��p��%�-ᚕ��� �WR�G��}�V��W84��/����E�>�d��l�d�m� ������Cul>����h�6����p��>�lB$6+n�x֑P����9I���6��W�O;�E~x�������xM� t��m!81����������q'�?��4�Ar`w\pl[�L��-%�ߔ\ �J(�N��.E�`���Ǿ�ek�?c���e���CK�|J{#�֏�����"[c-}8?��|��}w�;=��,��&��@��G�89A���!
�օH�`�J$0y�/Z�㑦~>H�ƫ�I�k��EV�Q���3�/LsѣWFŰ�,�5^�m�e�AbQ�	���9;�̢|nk��Eni�`������de`�+�P�5�rӖ���\���K9�����Z�&B�
��)����$��e.��_��Y�����lm��T�/�b�d
��&(��};�XH����i���ZR����"�6kr��qA|Q��a��W�:�����tN�G�}��J��dٛ4g�^@8@״�t�^��S;e-:?=7d��^-š9���Y�{�Yzi�ޚ���{�q�My�x�T8e���|S��?s�T[<�s��@���y_q��k�U�PK�4���'�zN��[���j�_��!�Uڪu�ު��r��fU�q�_>�cOT��atN��N�:�%�?Xz����>1|﵂��>�_�&�#�����t*G��y}�Z{��*w''�ԅ;z��C��oZ�t���?x�;7�~�X0�[�WY�������:z�V@B�1����Sa����Y*�;r����~hq+����\H-@/i�*Gr$����43fr|�"��ķ�q=�Ͻ�V3���~��{J��ýv�;I \KUNɃ>���3�Y-e�!�=�a����J�s�����?$�$�ery�p�'�$-v��@�0m:3TR	{�`�1��w�tύAeX���n.Ҵ�Q��Iӊ�!ܣ�Ns����p���س���zA��~��\�:�Q��˩q?��"O�;;À�#�J_,��K���Ū
I�V)I'��D�U�P��4��sa�l@/�y���E���k�c����tX3��h���2����}����V�$l�6�AC�|5Mx�(�(LA;lj~}Eݏ���zrU�K|���OE�."�g�E�igg@�N�V�:�W_װK��I��5��]/�����_R�n����o��~fH�ӵ7{�(��\�ۡ#��16�q c����:o�*�����ss���u�ք�ߩ��ٙ��0X�H&�.��5 3�Fu^>���`�i\�jH�H1��~+�a�5�X�!�`���v�	�9�V�K0�V�o|�w��i9���ϰE?��y� P������g�y�g`?�Iϩ.��i
b&H��<1Zb����o|v�`]��T�aR�_���q"sLަ԰A���G�
3_[�YclJmL��<&�f��QɣK���I��]�)�p#�*ɯx�2IC$��`��݆dٯ���-��8697�*�D)�;GZ�w���>�cz.�7���ګ/։h�:'�Ҿ#����V؇Oz��K�1�0�/G���t�8��Wo������Aom�`�2�Y��(����Xtr̕l�T]
"��_����T2������Q�6*��Ax��o���q��~# �0����?��A�$v�Ek&��U'ew�LV�@J�A���f´h ���WT��/.φ�4��;����	�B�.fكò�ۿyMV��~9�R0�۵S�h���T%ث��ۈdJ���I�;N��pz���V��/ ��z<�}X��^c�H�������\������E����uRԧ�fQ���n%;�0+�J���kRb��e���eډ���N��D���\1�`Ĉ\L��9C��*_fO98JQ�����5Ǣ�v%���'�s'ڝv#��+|k)O�Q�#�U�5�1�٥M���up����_3<�,='/�z���b�+L�qQ����ۻ6P_CB��z�1�u�Y�Y�>�њ|�[�
� �_��ù镦SB��{�8�����E�3r��FY5lr��`���KHr�_?�������C�_�ً�i�)��"��(F�����CCD�Ns��u!���!n����#a���v4˹!{�#�_�>���@�H<:V�wGD���|����,SGV<���`MR�R$�7m�[?m�Y۷%ѱt5�Β�T*O�B5ƞ�pfTo]r�ͅ��5�n�����Uca�S��<��n��N���k]�\o��⢌��5�� x�A%�"z"sU}E,݁f��>�}�����w��ak.�����<,GS��g�?&5Rǝ
�
��Dv��4/�XNM�y-���s�.&ԯFɍ���.�z�N�O�~ږe������O���;aR�1��ePtN�,��izvX�:u�r(0�w�;|� Vv@�2�=ٿG�ezo�L�g:�ݷ��3p%O�*D�΃��Zy��>����qn�.��&��em��b]^�$�r�"��a;�=l���%Wz1l8����1��wZ�u��4����������r��T�V�5�p�{֏b�e��Ǻ-Y�V� x���=D|�z�x�P�n��?-	 �"AA*9���I=	
N�	�������qyr��c��P%8@��~�U'�\v���66�@N��g<�ּ7)?7��?Nr�v�۰S��\f1��<�J'��kL�X졒�6�4��뽷5n����I}�	����.�I�$��,���(6b�f�A;�H��6Ո��<���6��(d@��7=r��I5�B�b��~�3{El:F4��̅�F���+Z<h+˳�d�Jy�2]��f��X��B�ÊF#B����t�F ���\f��6��u��iO��r�[��vtݹRd"����	�(��I(����, ��[ ��k�7�s�k��^m/�=���~p/����ľ1L��9,�%������R|��_ -���{÷�Y\�P��2Mm��9�	@�Yxћ�&DS��:�T�o�nI�����ɵ�u���Jް)�
B�&1��V��[d�T��U�_#k㡅��%A/X�ԇ��K�*�)�ٻ����]0\i��T�H��F��7�
b��u,��+n��X�h�}���*4�u���.��b~լ��5Z���P�4f�9��z���B�tJ&�f�� �	���C�S����Ѿ�a~�ȗ�l�M���Za	��6T+��f��N�
X��ʑ�����H��O(��/���S��9�`��qd���}�۽�YZN+�0���d�����ɝ�J0K��q�̬�w[�UU���an9�$)�������T� ��4Z�bS�`��
�dL�ֵ7��a]O_�b�c�HhCP�τ��Q�����i���=C�TׇLDp�ݭizX~��	"�P\�m�r_����q<R��/��a	��+#��-(YM0Kzٽ����V��y[��j�gn��g�i:t8�����SM7��T�n���pO���k���(���� �� ��x���k��T���PB��%ֲ��~�A�@tT�_#�R��
��H�"�������75���qnBׂG-¥
7o�KƜ�{���E`DI�2�3.-ޣ*6mvӸT�G��k���H��݈(<I_�u}t�w��?&n��ߠ}��u9mw	u�˽-� ��z���=�f�Nu3�Ō����	�A%l�`0CX
���_�&���&t��A�z��ְR�ʲlBSY8ݞ�cITeVBA�����U��,����.:������Խ�_}�c����>��3��iI��i��qzjL�N��?��+�/�&�d��J�>�_a����Hj��[6)�4;WӒ����}�LY�t|ֽ)m=�'�$�Gl�	�|e�|��L�;���@-��ԶJ��.��ԭ�X���{z�}��1��$g�U���PWKҞdhʸoG~Vw��������>R0j����#,F&$n��n��QG�H��!��(o�OD��'��������QC����{��s&j��5;��8��2�N;�C\Ǜ���8�"3��?��$�I
#���ڵ��2C��26O!)�HKt��4n��r|<�.��#�]X�#�ũ���`��7k���T����.!"��\�Ұ�!��4�5� R���`d���]٩0�X�>;�$
�ȡ�o�����GQ�4�O� Y��qZ
�^�¶�!!��v���9�&oj��E��8�2gתe�Jb�4N��5��%�T��%i�������*��"ҝ9\�3��b�B�1��;��pp�$4�i,<�	.��8�WF�"������_�u����Jɰ�.�&f?w��_�����kw7>{��Bb�����^IpD�)%���\���a|��[N��\�N��H�8���P��1�~W0��L�݊���⏙u�ޱ7]ͦ>�i�ʌ�!���[Jގ�ֿb�-Qʢ||���	`]����-�	��1p;�R+�0J/��J�|q��}Ǉ!N��<rL�����,c����Q������X�u�*��L�a�����/E鋻�z B�&,��E�%�7ljnA�6|U����N���u��ϯg���}Z�a��� V�pzJ��T�7Q�-����>;*>�0F	�VQ?A&�>���q�����I�]��0z_̥�=���4R-�!}݇)�N)��Ԫ[[��u�Ѣ���E�<�E��i�e��0
n���;d�M�!�z38��';�`��$Ӆ%����I��y��h6r�ދ��"�� Ț7��ᣙGV>k�?�\7���>�m8��{��&�=5���[y T�V��8�B�ZH_�w�����\I;��C��:�=v�ǌ8�|`f�]�o�"�j� bO��[���I��F�z]�`"�tu@Ϋ�ɧ�7,pɄ�0����n$h|Z <����ϲ 􅥴�VB{��	k�@�ٟ�1�];��z�m"ߠvW_�;*������*p�A�h��ڕ�yO�+�p�BD����w���OB�2��fm�5�,	sf[�
�/����C�S�l@_��Ui�cR��Ժ±2�f$]gT-�%io�����bA��Z���q9� 1�A�Pp�"7:���ְ��2{\��NM~W����L���%����@���H�%!�]m˒A� �3�k��3���Z��uo�no��8Bƅ�6��@ӣHO��A��^��g�e��th~��D��Yr�߼~r����b{z,l�0�c1���:��\�DJ�Ӕ��n�8���R���:) ��?����遌X?3���gxIL7����l���p�*IޔkcRB3ܰ�X3��b�xw�;^sU�״����LD��R#�CCؾj�qbTk5{�C�*����~%�rܦ�9EEkN���opm|�ܤB��c��}�m�����+�v��@Q��͹G������K7����i>�k`� 	����Ye6�����;�H�ŕH��wHvp�􂢱e%��-����>�vjO�m K����|�}�,�ikx�+�Z$��L�¥>9�T�h���u`V��TH�(ħ6J��%#��GX�މ��%�SO+6X�uy�7��bC��S�5�O�HD�P؉��?c��b�tZ��L��T{�0+�o�Cy�_L��ސ�.�\����3�t��һ��X1]�DR���o:	��r^�,�ܲ.=��]���Z��4�8����/9K���T�c6��Y�-ێ�U�?D;g��0���C�t�W�W�j&M"s�)	q5��	�P��[d�5�	U����.R{��)��D��I!�R�[v�ګ���1n�u،�&qLh� M�g;:ݦ��q�Lڹ���}����kޑ����	}*!	c_��.����+0u	t� �27���-��>
�|�;"��MayێÉ9P�Y�Y��2�u	F��DvB��Ҝ�H��dd4E�
h�r����%�=R41�PTmW�h�
a� HRY��&[e�`}�o�A~�WO�h��9�SҬ�B%ޝNg��p��0�J�<���	�G�W�35� ێ
:å�aE�o`.%��Qo��å�5�[��D��%Ud[)NFMݔiGD�]�̛$3b�r �h�7�D�of�[�o�i�U����vl�>!O���`�>&��5��怶z�Y��O��Y�d��j�_v��F�\D�Ǔ��C�eB������ntP��7�	��3ui�n�/yt-w����Ȕ��Sy�su�R ^�Q}-��?�˲ ttN��I�c��M��\w+�����Kb?$NZ� B��eeimн-T�NxG�̱5�L�F�X>�y��ց��{S���^�g��4t�EA�Ta�@�'F�vl�KA���%3L`S9:J�4z�HqZYd����C�܂��Hw�kgL����t{\�F����Qx����N`2M2AN�FJ�r�׆�٣]��j{#��W�,� ��:�@TO��+�:tCf��/��܆Ŗr�'酭�}u�E136�P�JN���h���u9糞��u��4�f|��!��%�#�_�yHV!��M�x8"�XF�q37 fF���4Rph6 ��>G߰��l3B�;AU>�(��$�Րl8���\s�/�a)����v�}������q�^l��?��9{v)�X��Bo��RTa��4I�E��|d�5E ��e ��ŵs�Z鮟�J3�{�O�|�2Y�㗊ѯ�|ir 5)�$EZ����D-Ũ�S��%�Z��R3�O_�H�l5.
�,GK�	9ũ����|Ae�����M}��S]At^@^H:"���j6 
���~h�4@��.��A�0���R�+ڰ;���A�M�V���,r�5p���h81E�8	��͉c�`�0��Yi�H�$���-�OGR���Ώ[�?@2k����)�$i�=��$��g�%�.�g��ܤ:��tqw�K h����R��!�b9�*�6c�	9��c
�\��,��'	H��	����B���T�5�� k�I2_�^���C����4�Х� ٲ��T@1���Ye_P�[��&V?�s �r?Dsݯ�U�'�%�-u$�{�R�߬�ذ6����}j�5+vh�2���g����b�s�j����yA-�t��};A���o��ݺ�͟ W�0`0uvR*��B�_)�X@9�-F�ۆ���O�m�����i�0�o����^�S�2�>CVނ���0� ��v���i��a��2aD���c���{�wA��8A��d��:�c���6y��#J|\�&ά��+ ���QԞ�v�=o�����Vӈ��z~�
���@m�|�3v���^�6����p���cm�䀘Q����7�I:�ae`��@���oH@"Q0<�˯�w%�w������Ơ��,�p�l�����ev^Ag=�����b(-��S��N�	]&�aWi�o������+��4\B[��<�G
P�dz4����ѪG�GXx"�Q6u�,��:ƓtjzVw��M[�|GX�������e<�i�qq M��b�=U�d�C@Hi�#"�=Y2-�ߡU�����(���+G5��1�=��@=�m��/�0&��X)u�����k3U��ķ�>�I@��W�S9��}����_n��p��ީ�Q%	k�����29�!�
S���E��+���Hy��F�uX&P�����ɣ�i5���p�U���3F���{�m�&]3ۼd͝>;��	�T:3.b[{G�Oo�R»ي�R��������c�x:ȩF���B��GB��u���C/���h�,�o�Rŉ���!�}wA�Ft<��Jf�-	+����D����СO����6�����;sYT�7J��gC���B[TI��%��C>QyAp<YO��_�b�O�Z�ᬿf�������;%0�����ow�gzқ`�V�{�W���NSw?	t���[�Ti�9 ��L�xCk�~i��F�\aCw.�އG���� ���� ��;
|v�nt���V>7�T���S�;8r����/�Q��ԃ!�9�� D������c�Q
z��A~|�K�̃����	�4��i��ӄ%c"��C�al�N��RƍK?�Һ�I/z�����1'bbF:AB ��ԥ���@"+l)p�,�>b�FZ�ge�Pm�C��x�~�h��o�/����cw�s4��]zZI�O�l�����ֲC�l� !L�b��ek~���Z��y������޻����;�`��V:SOx�Wh�x�Cu�[��������\�rn@%��G��OO�� �\�lѮ������3�g1V��k%�&��#?��fca�(�׮�1�)� ��h�W������za�(�٣����O��������GlFX=u��%w�n߰?'�p��hs pf��_��@�Z�F9��K��v���&�����1<H����=D]��	�Y�-km�J�e$D|�����>,+�Ə�gYf�yZ�Pl��R�b��9?���{m���ľ��z��	V��t�D���'�i8tlf�筀z�],�+��G.Y���z6�k>��8w��H����˻C�,�Y���-�v~&���Eİ�uϬ��G�Jު9	��{�HiJ�XI�)��'I�'�#��kѪ<�����#�=�a�ʿB�A�'�CH�s?!3���l@p�(u�<@�5_X�;��'%R6 ��l��pypU��,���]�yp�?��=����yl��s�Y����Ct�E��T�w��tVZj����A�������dL���r<��|����{E%�Z��|[..7��mX�zQ������C��G)�O�	��'z�yBEgKZ�+�T^8f^6���Z��ԥT'X�QP9�O�JW��Or?s^�/ƞ�4 �U��-'p����h5�5���(�q�ɿ�m�m� �O#���F���܎��k�±Ɛ�5��-��v��dBc�"��c2E�]܆���z��-�3&,�����;�B%�b�
�!..�w�g�7a��2B�Z�z��N�i�����G)�ޅ��s Yh�z�W���s�J��, w�'����y��5E2�ӳ�ا�o�z�<uJ�Ǝ$ǆ��|uhmU͢0��Ŷ�zl�>��-&�?o*>R��:2�]�%������L���쓂��ޖ"��"ePZ\��M��ň��N4�\0.:R%� �TO���#����.[�X�规	�烜�7�)Q���6�o�+��A+�C��3G�%è��3j:���Y;{���}�J��~���\��A-Y�������.��)���tĞ0���ex�����'0�EX3pxF�t��"��$nf����C�s�,:�mu����2J�$�u��e�xй���w/�hO�0K�Z]�X�".�C���;����=�����^r�Þ #M��O�Wb[����2aQa֞"�[zuδ����&q�3�ETh��տ�U��W�X~Q°�`�PDvT���W����|b��a� ~%�xb��Ø���@0�*��V7����^�;#MQȤ|3w��~I�a�-�������u�7�]�k\�3G`d�]���T�e�a�����Ά����z*� ��z/Ø��� �lLW�
��V*|��6#��EA�g
��crT�`�'G��R�]�.��[(؄��+6�'��]�cp8�hk(�Y�R����L�W� ";m`O~��*˫�ڼ�Q���T��4�I��}�N�i��u+e ��1�5�Ǿ��Ay����-+��L5�F}=�p�D8��s��w8Ure��(�;�o����\�Z�q/j��yc��wg'S�d�Z�a  �g����d�+&m禞�t#n��pĶF�bZ�Ǉ>����3�R^�~4ݕ���)^Y��h����	K���*l��C!��hUÚ-������*�aV�V�>�����m�H��_,��zg�ʆ,r'�BsG3��<e㵜w�_M� �������"��f���Ա���{iD�8�f7]~θdZ	�E��jX����\�ԇཋ�f�~��ٺ1�
�<����tt�/^�������/X'D4}����BF��qJܹ�����<����4=��j�7y8�`X�H���V�#���Y����z,��`'�AJ�|u�l��xv'o�Y\ ������[�G05؃mwt�p�$��_�%�&���|���:cE��]o��������r�����ڭ�b\�%��ma�� �^os��-ԡ�S#�>e��ן��/I
H�}�3��Bє���A����z)H�\N��䊹�r���r��h�~�_Γmt�2� ��+���� 4��
���:m�>�hv�)�D��2�MblV�2�h��_�U�L�;WO��V�/^<�$��?�����ܙ�:08*�ܴ�s���CU��aQ& n+R�,�,b��a�p)��s6'-F�����l=T���!�����8��rn�X�9io@L֕X�6t'؅k�5�}��g=ӡ,#�M�h�������ʨfX47K u�U�w�^�0�^ꕨ�)}9��RnA�tRVR��Q#h(NE`	�;���t��Ó�ˑs�@��D?��y�>����j�©�\�E��C	 #��ic���ʘ���n��{\�1�$�.��.�u���h4e��P���F��U,�R�S��C���;0�f��4����%�6��d����v4��`�А���������"���l籙��M�q�~)���#��#���������o�^0��?<����jp� i�*��Q��p�N F�2P(�MQ��*����&թ����]M�����d�ޏZ1�vץ-���o�Glб}Ճ�<z6B1��2�\�D|�t&Ӫ�1mLgk��י���M�����v�(��:�j���NNsDX�J�_���W��t=�;��J���@�K:^u��_]SS6�@F�Q��B� ��&�Qf��W2�	�%%�|N�J��z�K[D���2J�\5t��V����L�,�{s����:5��.��p���j�!���%u�_>z�7W	�K���k���B���<��.�Bv����zB&n
C���T�"�#����{���9�x8� c#|=��czT���9"�{*㬫����;>��/��b4��no�Y�,
�ԕ�Ä1�.IU�=	����p5�WL�c,I+=5=H1M}��Ƭ�+(�a�A�G-Ae+��
�FP�ن���;��:a�%�|��m�3}� ��O�1�XC�Lqvޓ2fl&�ԺKᨱ�~�ZR�khl��{��3}E]��S��_�p��2L}FMGz�y�43!~J�0��]��|�����ɏ��V� V�I�y	@��U*5��1�X��fr��Ll1�Yo�H}���z���qQ�5M�܅�"K��^>���<dԒffeo-:����%�cR�dÚf8w6D�^V��T�!��A��[��� ��'�iv��_
��1ZN����)`�KB�����r���\jѧ�|�#qkE�d�	m=cyZ�UW?�a6��1����Yb����]�ڒ	�D ���(�%geV�v��(nmk+�Mޱj
�-�����I�(6a/&؉��Ȳ��!�[��!,t�=��)�sJ�>sj/ǣ��ޭJT���}�m㶀�Pm�M�!�S)����?bf�o�~*��:-�0������M@j�O�=�ZEJ��y���� o����~��߬�B&�Q]�Ir7<��{*��,7b���eX��|E�{���/�;Ҍ�rq�.EM�i���X�T������5q��'��6���JtT�K艟���	�22��G8�����L{*����܄F��AŌd�j���@���(�a]h�����$��,Nz{���k�%f��F�kd���\���ĀE����p0k�y2*d�n��O����h8!@L=/k�V�ɪ|5�ٸ��[�� o3<�O���?bnuD����=@l �4+y�����Z@�{	av�F��Š���`�njR��y��d�`Y��kL
$��h�V�G�<�G�����d	���� ��),r:��v�i+o�C�"4-�$���4�o��/�+z+&.i#o�� &0�\]2�e�e���ܺq�x��� /�����vϧB��'Wf��#��S9��W�u�"����;����&9���#4av.�2�xF��cf�>ۀ
d��W�v��+�����-� ���N�6��.�X�#���u��3�!���黑�ϫqM�ⶊSy�Wrl'��t��j�q]��fu;����ũZic�gqf#�BO��'Vh�>M�\h��¾A{��M�*a-\��r����aQ��9���5*������/���1tֹ�b�"x�Ng
2��m-���Ր�ݹ�<f�>�����[��Ƅ>��Y]�����p�V��.���%B%��*�t�ӱ3b��C��P�+`�*oov�����ލ��[��SF��� �fO����ʆ�`�w�y�O��eo{�Jj����{���:�	K�_���h޿lo%)m�Y�EHz�O�,K����{׍rH�V&��IN�,���Ҕ|ǚg�/[|11|��azav1zҸ����Y����1��Я[�1"��/���x0����c�q��� �P��G,ɨ]%�_(���-F#]8�G|� O�x$KZ�[eqU�C5�8ڶ��#�<B����~@���f1��2��G�i�c`q�YM~��>VS,[}f��Z���Д�6���`\�۳:?A#��8�!���{c�spxBh�T�/��}����x��
�K�8�Q�ڷ8pB���a�L�rB�	z����||p�C^p������ch�S6o��޶�E�̓�ѥQ�F�=І�
If�tJ�ڶ(�0n��e��V�E�i+��p�7#����rT?1��N�Eww������@5�P�R�g}u�'��A��O�5;���r���������M[{��<��'\�ze��N�s}d��A^��C&��yfW<'¸�B:og6Ђt�m�F�<ǭ�ʐަn[��3,?Db��*��2� �W��W�Gp�Wё�꟥?�^|Nⴖ^�Шz�k/�(��`A��%Hł�qĥ��v���`z�Zg����\�/.63*�
���9�,�ҢJ�
+�A�X�h=y��H4�0a��B��,�[^K�;�AH�<(�o9��<H{M���PZ` �(+ ��w9�
�4�_a�X��'�.��?��H =Ľ��6q�~��x�
0��gT�$����8k�(��.8�9ՎN#.O%Yֈ87*4w ��&�|$Ȃg)����"�,�s�ׯ�uP�v�uQI=R�m٫�4a{�a�
���"�p��Ӻr��D�����R�+����I�w罃�����+����x+�����zf��NF@������e0,�b�܏�Qi{"iQG������sz���p
O�<V�$>h�Pz��l�)�WY���[hA��/��G^��{�r��+��&�w�ۥ{���z�|��5歷�6 ��$�XY	=���&Bѵ�\��(zVOV`�`��M����qv�;X��jF�݈fd�=O�H��U��E0B	��r��t�p/�$X���~�63�4�Us�yC'���DӚ���U�w���A����5��I1��ݧV��ps�m$�f�&�"�5��'ٕe��e��#`�)_X
�IjvC�N��n����H�`���� ������lw��P?͐�m���_��"��c?3f������^�e�������e��-�Q�Z�IK�g�3�oՕ=�� #@�\����f�O6�QԤ39�	�D����p/ -��.2_p �Έ^]�6!F�
ޡ�ֺX�Mi�Z̎�k����j�Z���M­,���[�G��f�-?�Y��qh�����u�dm�gB���u��S��b�'��O�TU^�c3�X������>$H5%!Ǌ�6f�u�yU���t���nQ��2�S*;uN�'�����_!���ch�q��c�b�	��ˎ��Q�'�� ����'�<�S�De�8#C��j[^�SI	2����^�����yp�ً| ��d�e�ip�ُuI�A9�#J�vf�$�ڴx����0i�Fj��({���|f�n��F�_��=��<K
&�2!�.F�4��`�<G�G����$�Q�����	,��^�xH3W��׭�V���A!�즞�P���Pb��_?�ko�*�؂����`�&3�a=�רDa*�>��.�i�R�C�����׋�FW_Q�)����3�?�U��|�����s,j�h�	wd�Pm��#h@���0���apr��5��%`�R����G/p���,�I|˸{�Y�� ��Y�r4Jib2l���*�9- ��t�^E���Vm��:�'�!Y�,�p��1���.��g�=9�D ]��aky�@(6�.�?�@��DJ5��Y����;��`�&�+��ͤ��Ky�q�S&�H����\h���q��1�]�����9����I}�H��11TQ(��ʥ6�BFt��+!���s���>ғ��TL�.�yU�mWJ���J�_������X�;]Vg@�Dv|p��R�@�!zf�\�:��ʤ�b#����I�#���I$Ӵ��=��T4P&^--^
ik&�ڧ���� ~��OeE�K���R��=Ԕ����_���_> 1�������{x��.:C���c�O6\<9�"��h�Ef|7�������v�@��x�Q�-A�Y�>��i*�)kBI�k��8�΁�	?fp�n��V'RC���y�ӯ���3B�!ao�o��O�w���v_�r2<g]n]��)>"�A��8�`�����Lv��[�g
:�껛��@
=(���5�g�DT�� �aͭ$�I���rZ�T|�4x��4	�bĘ�U��Od֛-تu�$����v�7�����f���i�I�(F��X�Z`�-��X�O��Ժ��|l�uΧ�b�l�by��-�B�VT�;�&sQ��jg�
�CO;��.˝2kA4�LX%��
�|�l+���`	����r3|}����fV�	I� ��.S�W��,���?��+z߰���V(��8x�O��(R5s�#��M�q��<�t�To�|���%<3bib
� xNOX�q���%��Sg�9�z���]^�PW��;�g�>#��F���V�_�;���ߚGq���8H�܀���ݳ��a��~�'�}��z �i�.���[�y�g��������չ?���<δ.O=���Eu	˞.��lR+>��<�Q��n�(�����m��&�"����:�
��l]A�A�}dg�{<��FlN����2?�)U7�\�&q��5�&�����]n���X����V<�d�ή��`ȱ�`������ۡp�P,�MX�G�<�v���&��n���,��=1���C1%�1���	̷��҆Q�������� �S�D��X&�?'@G��,;�/\�#(����:)�����*C�����U�}��Qf��ƀ ���
t��_�}�g�@*��%��WO�jq�����y�j��
~�ق�B�p���p"Ա(���! �@�	a�D�˖Z���,K�N�b5��A�:sB���:����WÆ+{]�"�f���
�O�D�{zUsf�8��M��߆�O�c́��\S��U�zA�[�H)kϿ���x4�k(�.���Bt!m�R�:�:�7�"���*��f�YB�&VjM �*
�2��S�L�;�s�F�0�N�%��ex)��\ꍧ�Eor�F1fki�5�#�����;b�JcY��V�'>[W+p��m�Çը��o�Wc�d_�e$�s�ĭ�DQ�{v���/݊Yp�m�BO����<e��&�(G�{W_��V�Ƒ`3}��f=ԑ�v�5M_�i��t}�#���:$lXq�H��m�:�k��ת�R��v�����p8�ݬ�P���P�v؅k#�C����~}���"��c�E:(F�`���|Fr`kn#}�( 1暳�Ffm�T�\�4�ಱ|��3�F$���g����6Gc��sG�0K�?iA�u����'�7�p��~\e���� j�[�KX�P�R\/T�����ϴm��z�H6NZ�L{ 5�7=T��.���ÕCo�A%��Ë�L�nn/���-fX"B]���eq(m�~(�T�q��W�m����@�� �?��:5M��A�7�W�fߓ���U����i��NQP���pc#�_B�[~�Ic�B?�l'U��R֕%��ә*d���f����>i��� y��l~�s,gͺ�'��j�J7��cX$��l�*y�0��F=5Q�,˅�����'�D�L���B�#��4�
��hT8r	?n�h��jX��f�8��ϝ���HP̍�&7���I�>R���^��KS@k96�|XoT���ݤ��a޳P�^7�[��#����x����:)&C1�űng�Ri_X�o�
"U��m5_�v`����}Z��yi�n#�5S<�i��ra�~��7Y��o$p��O�� ����u��)O��CT#��b��5���c��2��GS^�wZ�3,�;lꉛ=��;��bmY�N6珯'aS��;��ܕb.C�o�Kz+Zw\S�=�X("��K�]Kgm��b ���6�	p��@�(�����:��[������.�Auz�&�����hX?jY�-�o%9����>*�4�s�ы��
��*�'f�BjSCI��(7�Ex7�j?��{:x����ɼ
-o��������.�N
s��,>�z�S��{���?�{�l��X�C�D��;tC��{x�g�@3�^9���	�yߋ�' Cր�*dz���#X���OO-�MG+��\�bz��F��/�}[�^^J�I��0����7꬗�M?�X�ҹ#H�G�)-�����4o�o8w*�āl��'
<�m�*�\�c�>q��AB{_��H O��&��zU$���ǹ 5ʂ�GF�9w����=.��T�^x"��9I�:d�����3y��u���x�.3�h�	uwU�I��;x�x��n#�#�K��,�N���KZ����IE��5�Y�I�ꓫ[�}���Ķ��ژ~&�>�l���0�S�H4�Eq��=d���+���I�ӓ7	�W@� s$��j=L����UÃѱ��F�7��'NP���*.��I�@E�]�� 7a�O/*������>��h�wɾ�����r&�e��OStu����t�V���Z�4�ҩٖ-�-��|�}t�4�+��cΚ$c�]�wo�N�&�w�)ܾ1b���RƉjD�����`��e���+O����K�������%xE[������&�|Р�N<�X��1�D������֘jY-czŸ�i֣o���"EC�����mT!�Ky�M� �c5�L���9e���l�,p����NA��z`���?gs(\-H�}DV�@�9K�yzx�P��*&v&� 6}�`��`N�̿gV���=cdV)��!�R�O�TY�
NH�No�n��7	4���؛�(�K���ц��ďŞW>Ў�O��!����"��FtYk���˨�^��G���I���D���m��/��߭!��Y�'��mc����)��¾�
�󊦖�b�_��C�ake$�) `����ve(?e�<+f>&�n��Ti�Ӑ�J�pE��L聾�;���v�7���kA�I*\I���ܮvm$&ۖ��O�O�Y���M��/�q�@�{�x�TX[1�J�+mp%�n����T�V]��\�M'���W28j�E�z#9>�6v❮�>q���=�J��S�oO�ה�mGYt�?.gbjɻ�����lc��O�ysa�`�g��nm��-�/+=� �fL`�9������[���73�Y����C�)S @s+W�!!���ʾb��a��\ց�r���B
�cz��w� ��UQϯJ��+��J���D:3�raA�>X�>�1��8,���Z�uy��-U��R��jX�.��k
 @�>;��g�у[��J��qI�����w�󬭠B-�t��q=Ip�C���Im98���J..�B��8���Z���=���^��)����ȏە�>�샲��Fu3Y+�ۧ�5�1b���HÈ6��AW^�����L�����+�I�)�cV�����ihA������C�^&4�M�ω�S#Z�����O����s����M)��]�	d8��r����J`H/�U����nH�����������Z���^6��,��.|��0~�R3�ംOuI����X���-�d`�W��6w�"�F_spu���΁N7Ѐ^ѻ1�,c�7xer_#�Mx��aQ�vK˵�uz*�5NՋ�;��
tU?��hlґ8Y�	bs�
g�q��K��{Jf�ڬ1ZB[}�6�ݛЖLq�Mt3����\�A���@���U�����u���?��)p��mxy ����ʇ���t֞G��a`�'��Q�K�p��^-�*kQ�w�F<�ټ� q�����I�c�י`���-���T���?�'n#Dn�Ix�?�w	�ː��iS9*�&c+2���5?�ΛT�@:.��:wON=c��M�fRg�X�j8�;�=�El���m��aQ.�A�јDA}:VH{�SR�i��ȁ~��4��hO���MqW�c	�ߒ��ZW4F������B_g {��v(ZWC�N�K؊���N�E��\������$��p	���I�ݖU��+5�~~�p�Q���Gg5�.��\֒�`񿏜N�/��Ȃ8*�8�`�-4�7q���+P��vZ�����"f�iֽ��p�v/�{��Ԃ�t����^V���F�v��ai����i��*��]r�������bQR�W��ǌ�F���� z�ч=}�Y�5�Cۍlu~�kgtp�փ�m��pmV�9���6�WH�������aS#�Ɉ~�QJ�H�D���żlA����5��T�㹲�,T����*�|v�0W��dNM�������V�;$�lzj�2����s��I��}�mM�=�{0�~E%F4Y�oIe.y��'�5��|u�p{�iؕ�\e8K�D��-a!��/'�K$�����Q:�\�2\����y 0l(�0K?ϼI�g���r�SU����<n���G.޸/:U���NJ��YZ�[��Ÿ/I{9+P���|4�
�"���S����>s�	����#�ٚ�� (��B�ݛ%c��Q���4�����xi�Scf����h�A���Jy�ʚ}����<]jJ��S(;'?��;M`_��Gg�;���E����s)q6����D�^�).D��Sˋ��i��ei��s.� K�Z�b5��L�a��0��� ������w䲑�1X���5��.�K��hK�K�l�� <I�s|�S"�_��X��\&#<&�����:}!�g��dRw�Ϋ���IE�{�*
���������O=��[�D9��{N
�1Y��F{P��w���<c���S�;������Ao�`D���є8r	���KW�t������s��F�� %����7	;��E��|�E��LH�q \b.��DmQ2˔S͢Ei	W��S?'���7mi(EӨ��7=��ã�v$�Z�����?�Cb �c����>����	٪�K��-�ELK6���Ti!����R�,�8�����ZJ�c�`:8���j����~,���5��R�g5 J���� c�j� ������+�҅.�˧p_���s-�$3.f�@��(pTkl�a�r�>n�{A�T}�	h3s�M�z�S������\RS�Uh:p��Shk�|��k^P��ߖl��#�?��/k&q�J�%��0�=��1�F`$�Gv˄��>d������������WZ��w�iw��V{߆�x������|k_g��83��f���F����[�	��P��Ԛ����0!����ֳ{��K.g�u%�$�s�zWs.$���,�d�����ʇ4�����e�F��n�){�tz[�Д�K�D���V8$������4�$��s�1KS�F� �Br=�S`��f�`��D��dwQ��Tb��bJ�۶�:yQO�+-4g�!�W�����������AV?$�m�7�F����7 ���+�s��L}�mlVjê+�]�H���o�aj�c����@DBe�k�����%3�2̦8#8��2kPĞ-�!&�wuV��rcQID�5nZf)�{5�b=�A���x ����)�"a�qu�[�d ��Nc��ǿ���I�vG��2���-�a�ZT��Q<D�
Oԟ'*��yK���zA�r���9�dK�~���_W��/s<���[mW�]�j��2����r�wB�KO�1j٧HA����Yb��|S�_�p���=j�T]��̜3C�
��i�N�;��<#�&�\XO���J��B����B��o�8R5
��}��PMk.��ADbNB�Vݟ�ml�A������"�S�Y8=^ԓ���.��?-R\�#=�L�]�D�hఴ8)&d�~�>��f^�.�>��]y	�n��c�&�l*$aL>9!�0yM+���U��J��ӝ>P�Bx
��	ׯrJ鶯/��|��Jį�EC\\�J�����ŝY{�+Đ����z���J��u�i���>G=���+��>��H�3,��s����}P�R��v-v�)o(n��߰/��T�cT���j:����e
F�2e��pi�&p��_�3yu���$�:�ܑ�۴צd�	U[3@cG�����%�i�M�Y�Eۂ�v�x3_A��zn�`Y	��\`���E�dJB?�q ����r_��0ⱀG�"��x�qMo���S�Ia��t�*$�5u�9�D�hwp�YYRq��9'b|%���yiޜ�yQnq=�B�Wi|_-��:4W�xE�X(�m �x-Q�zM޿,Q9c2�����w��g5+{ڒ�WS������
�-���'����`VK���eGl�=6��5g�2P�/G������"B�-+���Q�  �M}�z� L����W^D~�C�F;W4���E��E�ejh�خ�����B .��~����65���>p��x���LE񧏫v���)��xf�|;�ɦ)�܌@�)�2RV�������&��Z0�����e�̡�#�)Ї�-B�i����D�^�e�K��#����+��q�l�_���j��3�!�EдH�#�{�I @�&�:}qt��HQVz��s�u��%=~� �-H�Ŋ��9�0"YT�l7�i>/:e�|�|S�+�7�NJ���ʱ����@�����Ԩ��j>#�h����nF������	�/�$�2hp�P!]���}�ȹ{��R� �3��l�w�"��2�Q�6�b�_��/�Y�'�;^�?�^:��������Ae�}�;0$��I���S���� V}u�����`iCU^�%�F�F���liؚ?�L�z J�q�c,2����-��
����o������s��KPDFL�ā=�%1�W&����r�[�-��V���B����S-�}XHjaoE��3m�F�3Om��
H8����G�*@��4����hrড়�h��9����OV5Z1׳�獀��`e���o�yr��fօo.�ul����7}�Q&!� �YɁc=��o&4Zz���5,J�!���J�=7� ���PWW���͏���̙S2��H�{XYJ�9����h(��K�
����m*�_Y�	��z)@�HA����r��5��W���49�i��0�	<w@�װ�5���YW��"�P�S����Dǃ�K����J.sΈ��,���A��?���J�c�"3��T/��C3 9�`Au�^e�e��vۥd7ײh��S(u�	/�&�i�w��-1Z9���B�����X�9ؒ� �{I��7����p?��%���PF~Y#�۸�솩�»e�ƙ;��&�ϿL�ꇰO	�L��AV�k{��y��Md��h�Mc.�>�+AK~�dcﴶ���ꊭo�:ڇwq�0��S�=��<mo�+͉��ݮc	$�,�O��E�Fe\}8��W R�/�c�[h9���U��Wl����z.�׿`���;�-��`��T����QΗ��N�SuMy�de���ˑ��,��D�j�vs�nZ��5����]ny�~e
�E[P�9���N�q!�B>��
	��8D��W�"f�F�^�φ�	��c��E�'n"�ϒ�=���M ��{�3<�&P�ۓ�FԮV�[m�	�)V	i�ʤTD��J�����0N%r�Y���x�)�9�U�=�U<cE�y����g�0`�37AtL����o��IjCh2��������]ܕF��A�Y��)���B�I �
HSMTf1�����?�'�2�}�$ܡ��� ^H���r�DW��e6c$�i-����|a�loA���Ȋz��J`¯�j�<ӔE�8�� PY~9�y,\���c�{�R��*����S����V�p?"�HO�
,��c�YD28
2��F����p�_׽8� �7W���xhޞ��Ig`-�x�^jhvA��D;B��P#~v���,y��O���z,P�Dd��,�"z�Kh�G$���o�,w���&�Q�4��|�Hƻ,M��Ψmux �)�_���BP[u_��!�a2c�B�䯸O�3P��}��.�����Sf��~���/�Y�q��D�ȌLC���@AΞ;=ǧ�\~*,w3Je��Y[�Zؕ�bn#��%׭ґHq���P=�*x�9�~�㬳̟
��|�u��ޙVi��>X.q)�����l�Nv��#l�)������A�p�,��S��|�� �����LBg�:~.�4�HTR�	\W���
ݸy;��f:V�-�����5:e�w?���S "���ɵ�E�c��^F��l�L�ʖ!na��p�l����!�T0���ц\[����X>;��ߵ�BX�q:��c|.V�B]&�ҟ�-�	Zo�����`P�tl�l�.;%wo윋�c-��:s8ͦ{��vbϮ;�k�n��zE6h�J�5%�͛��*�۳d�U�c�}�/���u0���Kg�f~w�	��APf}e{G�B��"��)���~"@%��g��F������-���'�=����U"���w0j|�/-w]��<"�S��E�l������ ����\~���9��^b�=�Ec�^��(dx������R�uf�O�]c�z�����3�s��7du2�X��֬}��v����$�����Z��c�Ys�k4����w��6�}X�/�W��h�(��i�uH��0�UMr��;
�l�i�o�Ӄ�� �'�����H>�(9ڛZ��6C�J������^���C�"��\�TzXs��B��[�7���o��v3./�>��G?�.���7�\b�Č��2Y���e���Ӄ_�Ԧ�7$�՜���G,�P<�B�q�
��2�j ���{-�'��#	�EF��f��;����J��C�T�~]j���̂�\k,����YÌ'�'0 D� @z��k�B��S)�(	͑ )U�4'��b�?6���֊�S��0�~n$}�mr�*�a�%���b���Uq�`��7���{�0��B������Mgh-!QonK�I�������#�9����/��p_sl�)���)�w��qҜ���n�E e�,.��3�;ne�#Vc�%�E�\V��4��:BD(�B�rp�y�[&+�t�l3cd8+j����hOR�C�?��!p�������mtd��`�C����}��*@���+��G*[[��><� �^p$�����[��L��`���qs�9�d�*�v3[N}�=fgR|d��q'x�0�R�\�r!~) \g��8!�mC9;��X:+�����{���(=ٛٸ�L�v���gV�K��X�q�Vsc&�Y)���'X{H�%x⌂OkNq�t����q<�s�%����Iʮ>���B��a41p�|4nG�֛�p�d�tk�iz0�~GmI���&��]C�s�Rh�����"��C�JHZVL@S�t:v.�߹d�V۸m�qg�Ě���
�~���#k��2�p�1�)���?@���(��1�[B�.r��>K��-ڀ�hD��ӕ] 
@�:J&7����cGΨ%�hFP�_>�� �m$� v���,����)t�e��J���$�J�Y�${��JU��d����L
탊��1�u���?7{Ȝ���~^4rSA�#�8)�M���2������3�U�FnP�h�� ��DU>}�`Qm ��b(�"{���-L��d�B��E+��EQ8��˩�٫�N��H�ܸ�u���X�@
n�z�B��h�棽 1Kū�-��I@�#�co���'Ӯ^���ny��(�Q���X��:v/Ov��U\�	���Ҟ��j�`�l��-õ���7�]�Pq҃x1Ż6�/H}�<+�@nw3��3��9�ò��k44h���j��#x0�k�����E�GH��ʙ���}v��U�;+^<I�b�g��	\�/y~)9���e���+�)����cJ�W�A5�9�v��*�p����0���6��`�_�PRpx #��أ@-$��
���oVCżV��G�t�1�Zu��c~Z����`�a����Z���y	X.��q*O�>-�*�vf�]�!x��_
m�JX����`�qL;O�k��U˘џ�f���=�5�2����9O{��L���rE'/�w�&����KپV|���\l�%$�3�d�����Lpj�^ �	
 e�r4,fS�J�9Xh1Pi\�uAw���-p���v�I�4�V_@�fI�2�p�����!��o�]�V������[�C�E������ة�,LN��Y$�h�����-.������;ԨNf$��8s��2{�AI&c���Q�fe:���nw���iR�h<ٸ^�Lx�"1w)�Ӊa�9�$�5�i��D�S_�堅����O����m��Q�;�{���Ř�*�����sY�sv�MK��j5}�*��Ѐ|(��q42<Z_&u���"�}'t��S��	;��������(�8�9���$���TԻ1�Z^H�~����ʧ׾�%��|��2���2)��k
c�g�j2��\�讇�q]� *���N`h�g��6�ݣ�?@�/��:��濍�B�*�ʿM�g;�j52�O��߫��n��w3=p��jt��|�8�Q���"�%a��'4X� <� �B��A_���i��'X���Qkz;�騀�0o8Z��W�]h�D{e������&U0X�d����ݕ�N�o%��H�U	=�w4��35�U�����fr#ޓ���z�ۭf��%�i���[�?#h}6���KQBY����)����͠�ýwk����Q��γ��
9@���nػ�E�aj �%֖�O�$��R��:��d<�N4�U���RYo;����H��NQTB�ˣ2]��ۇ��g[%���Z�J�z^d��}2���*��]Ĵ14j��6��],(עL)Ā*ϚPCp�>��W�!���E�eJ)>�`I��e.,R��2t�DUl���=�1��-����Ι�s ���;��!''>@W��v�kت��mH�A���@:�U�.���0{���޸��f�IZ��l�5�^S��N�ɑ����"�����O��tT�Ŵ�q���V.Jg(��zCJ��[�Z2�F�o�E}��OUR��)�5�g�ږ��"�\���E�"��K/
���v�F�-������?H���p5��lokD��Ɇ���-$�_�J���X���7��կ�Q�{`gK,>�!�"�i�A`fF�)3e�F������T���Al_�p���Рk�^U!Y&DM�FP���wbm���`����Q�ńH�~Ur�n��	)�d��^R��K���C�pz���ӽ"Grzci��2�����.�O4gn�B�TWA6�Å�������z&S���~��د+����7zN�_l���#+�Gh� ���_�}(�@��T�N��?mm'�DSQL^�kIUEk����13���;��05	`У�5 sD�:����Iǜz�Z����e�x��s�wƻ���`�M�H\FR�V>��O�+Ey
������/�6�+e� �eX1�L�'/7Q��E;LZU/����ȉ�%���&Q�.�Uy�_�P,m�j���h G�[p���٫��ʟ�I^g?�ѥ��k-���@1��/}���;E��f,Ш��u��}��#��l�(��ޗa$�}9 �g��SvMA6V�5�x���f��3� �D+	���p�:���~w�yH�1�I���v<{��]�)�h�sMђCn`�&�L�TΟ����/�;EF�lS�v��Jw��_՛c;�������rҹg�H�;��aÀ<��[��� 1�cǳ�c��Yx=�F��s3o�Z7�Bx��s>�@�4F��-�woߍ���6�w�w�>��ج!�Xۥ=W�L9��ٕ�� =������fa���=/���E�E�R�?�:8퓻X�?���yzL��7Rn&��o.*UE��k����̝&7����Q��a$s����d�&�@B;�p"��L�ɟb�RE[�Yuu��Wj�L0��y���A"��D9�T�g���]E��N��[�Ruǐp�'�����S�d�:��J����1���X�N�h�nB�Z���'1�9��;����-��QG؛}�6��x�"�&��]���g`����Gp�4�˫�!�J�|�'�1#��E~d���̏~"����0R�eW�������]���p�R��Z�K�t]�f����Ӵ��x5�.�Y����@�םE#uj�Nh��(Vx���ٰ�ϳ�
��]Y��K!�T�~���?k~3&KC�$��y8N4�6��y�i�+��c���AP��c��7��]3��FGA���b� �C���z,��4s�[r��s?!�r�e��R��O��pK����}�*Y��J���a�WcN1	t���e�q����R��R��֝r�R)����E)�dnJ L2i�dH���i|�f���lc*`�h�Hֵ�q 㯕297K�[��b��:���ܼF'��Cea�L������5���?#��~9��+&�up����7�����n����7��M�U��VI�fV���۪��G�����!���f%�/+v����j��� 3�$����`����g:���`۳*,БwY��U:�wQ	�2��Cf	9�=I]�|��4������$p̾��_,�+�/���������@6.N�Udſ�����A��	u)�w�,�~��5Q�j-���u��V2�>y��+���Sw9.�����*��-MBf�bO��D0�1[�i�?��p���cZH�Y��ݷ���F�;���m0y�|�u�J�*�9F��w���\�������0g��h�B���U�qʬ�Y���?��jF�C�g��*v$��0/�Қ7n��!5n`,g�Ή�����b�{���5�]�4�"Αd�?"?�tx���m�r�(���~�y��-�_a<r�R����a�lh��y�&+$��/�,2m�������R�2�˝���~TW㐗�\�~Z�3`U9_N�9У���Λ���9��T[�j�I*�-;�93� f{5>E}rc�<O�,������;P6����a|��I���q���J�~����y���u�{���0�	-Ev�����T��{�-��Bcp-F@�љj!i}�3���@ӬX䚍�9������''H�4��t��r�y��nT�}�ڃ�RI�Kt�=�� ��y�T�|�p�&��>l
ŉ-I��U�dR����9���A+9�E���m�+
�H{]h��+E���v`�8`3K1PE��*�G@=w��%����x���ѽ�����f��|W�
"*�]d+4�C&�Q�wCM3��T��*2����w�H�-������49�A ���4BT���a`Eז5���4K>Iax�9L�FY�������>����9�*�_�`~DX8���U��`hw@x�x(�{}��d~���[��,�\�]�]��0Qx+l����E���3��U4g�ܰ$BC�k�F�e�^F|H��,�c��'�36�W�PF�AzUy��J���)Z3�I*	������:F#��mr&삸]��A@���xJ����l%���.�eZ��O��Z���Z�Z�6�'����B}��I��K��5�5���n� 1E����W6���@�p�@B�\����>���{ԣ¬;��2,���3�LR鸬\=��Ѓ��.�C&F]C��"�S���PR2��7&��֡�mrOe�[�PY:�ĀbzЅ�nܖ���7*��q��z��#3��	�a���M�-�ah�pj:���;'@�{��g����0Q�3�����>���1j}��~�h�ɸ<K"��৑��yF_��yʾ�}Z�9I~���,p�5Y�e�xǜ8�V��Ա��z�w���0�{Y jW�� !�7��c��o�ENECiqT�/,/�DN�GZޖ��8�:7%��,��
���k���-� )��(hd�(`@��z��V���mQ�V������yG;H')���Y�F)e���2�6Q\Xbg�@S���y�f��*�z*�5��F5�|o(0�</�k�kp�*_�W� .,� @-	^��	�	��<f#_n��_��ې�ռ���r�ڀ�}́�g��ɧ���p+�3��Q7Xzn�*U�ߞ�?Z�mL�c��ݼ���JV����ٌم��,.
�
��[�n�x��w�̮K!�&OJC��ne��"�7��f���ȥ����k�<=x�}^Z��xF�L��پ[ �#kR����<t���g�gh��O[n�k3Igp���KL9p��X�(�'��EMA�T��W��wUon��T6�}&�ŒF0k��|���V��S��>�v&`M�"R�E�oj���-�5^$\���#�z�� �HB� l�]��~d�lUWP�G�1H��g�d��Έf���h�ǻ@J�]6(R-��m2��_��S�"D�����9m���d\��2�4����bY&���PJ`��]���1�!�`�n6���#�1���2�P���3��9��R%9��B��h��=UDN1,/|)���d��(�R�-$j�±Mo��q��e��y������Z,�RR���c��>d��۶���4�� i����xhd��c�N��k9^��t9�S��e�\�$��˟�L�ͅw��Y��R=����(�W�毾���l��5@\�������k�&�B�z�S��m.�����'	�^G�U��0��{N؟�޷QN�Lu��*�:�ǈ1�U��O�x�s`�O��z�i��*��������Ȗ���FB����LRG��	�3��g--l���r���D��
��&KJP�a�LX�K;x�v_?�Y�v#B�]�~y6��A�����-A�R����S��Gt3�X��(���g`e.�jl����NBD��-�t/�Թ��+��~ݣ^�͏�ivb���U2�~�$�2�<�֧L1<�n1K3�u[��f<�w_p$!|�@m��š�<��L��A_�"x:k�!�m��y��[�ؖ�]��bՋo� ��^�3�:-mu����x�L�t��҉���U����>^�S��
Hi���7��$ǹZc�~�~[�͘km�w?��N� Drz�t@܆M�K����00��S+_�B�wq�?�N�CTT�5#� kJ��ӫ��Q�H�����xJq/?AWc��KFT^�[a!<��q!�O9i#���������+�ZŶ�"���F��G_Ow��D��S��Mw ��T��?:��G�7�Rytǡ"���"V�iv���|�	;Z,Z�I�:@�!�Ĝ6Z����529�FB���| @�Q�a�I�/��d�0���	���wk��6�,��=`ϑ�h4|}YQ��[$E��zq��/T�i�ޢ��i�o�FJ�~��1�����^���P��X�3S�l���t�1N�q��B�L�9����YvPaW������M��
�xõ;���[��D#�#�EC�U�w����C�3��٪�v�5@l�8CW?t>ۓ���<mM,�q�>$ �ҹF~o��VX�S_qe�"j�ѧ�*��?q��L�~�p��B�}R�&���iG��i��*�p_UeXj��)k:yW�2|"�;��l�±�!A���q/-�� ;�zl��;��[.��Xa�c+��}J��Gg?�Ox�C��9ȑB����B�8��^��ce�A�Y燃�vB�`F74��>���R�D��O_�.Ō������+��c�����,�x����R���|����%Ŵ��$me��Yj�����6�gI��6�c�: q�1;7�P�cN��d��\-{S	�#�K��|Y� �Լ>/�0/5�9�~^v �"κ�G�����/6�������=U�G S�'��%��f�����(��Oao��.�[k��ӈr٠������+���5��\��b����~7�>��a�c���r��
�$����
��%d8�x}��5!*e|�\\0(�G�����&+2 $��<^�������]k!;�䦡�5=��p-�n�/ %������E�?�X%GJ�X�{�F�s���
�:�*� *(�Q�?�7���j��l��iO������������Hs��I���L �Cߙ����@��95�������8	|�sF��+��;���!ʥ�HYGI�|��z�'+��?P��B�P؈_b��g,�5���~-m��6v[��w���HUa��sۤ���(F�C5,B�,}3H�����6�!A�c"{7�I+�D�,���!-H�g�����gCF�Ug�J>S,b3:P�"s 61N2q�0����p?qN�z��{%(�����K�!vJ+�W��vwY�I��К湄`v��&a�;�U�A]��C�s���ޅ߳`)c��n�1!I
������S���AB�%��b�����ɵD ë�����}�D���,��7{�FnB�ݭ͑��a�Pr.�P��Eu8	]�otWN�;��g��(^Ѹ��<�3�}=Ϊ0�����ǩb�L��W̽�O[�J|�[�=�0ܝ_[��r[DX��~���U�c�;zj�W�7�x�`���n��<E)�Al�}��=q�8ӦW���(P		.����H@ɞ���Lh�x��<X�����	�ř�\{�<����?I$q�*գЖCI���D�H�u7����& (C�V�B�t��DJ���T�ϞP469w��U�&�|�"�*���Ӭ�v�D�Y���]�2���DIN�E�b�/Hy5_��#*��.����M|�&��MG���ku� H�M���y;柣b����)k"5]��K�DxVnv����;�"�el<�.E�������m�j��y
;<�#帼f+L��C8��R�)#^C1N�RaȻ�b�Z9��h?T[�` !x�{@:�gO���<%�:f=�쬾�[���lo��2vhRc��9�E�E᳓�����2p5��548YI�����E�w!:�P޶8��;�Y�	�Ic�d�88t�Z¤jߊ%�H<�i-SҖ1^����)�`B�������e��T>-�"F��z��o�[�D'L�Q��A�ZD)HO���J/������m����A������������}���Dϳ	��a�｢�æ���s��ʂ�b�x�����s9uۓ�Rn�M��p�NH��m��ɐ>.��>RGv	����y�Hě֔7�Co����C����ݝ�t�5��Z�yo9�}h�pϝ*�[R�cB@�;�O��0�!�I�6^;ݶ��w@���!�E���˞F�E�ˢ�ь�ځ�ɵ(�A�G��]y xFIc�"WRi+a�����)�;��5��k(�q�)�Uff)]�@�Ԁb�{�̂"[���΂���#��WhJ6C�Z]�J�!�i\z�,m�C��Gr��AN�*�F��Gk��4�2/!6��/pǥ�U1�y���e55�mv��u��_s��l��$4p�9p��XpG�:pB�gR�)����� �(-c1L�*&&��; i#�Ze�W弌wqk�)6M턊����.��k�(K�̟�۟�.Ҁ!y`���<��L6$]j��1M�����K�,�{&y�7� E�"	�䔭&�L;�!�F�V�^��+Z�w�*�dD��\
����N� O,>�b��Ώ��`�6�+J>��lh$�]ǫ�C��A�ʇO`���D5���ve3��l����q��CS�V0]�Y���\U.?Ŀ ���i�}��*�ǁzʰ˭q'.�������{_���>���ywk\�^�_�^:��u�s]~`�R���<*��}��A:z��*�ŕ+�C�4��a�#��l`fy-�AW�T�5"ɭ�MI��ʆ�E��W9öG�$�����w[M��S�N���*k�� ��w/��;�t����ݮ�~i��0��*�z �\|�9��>�%o�z��R�3L�O��2G7�6~3��aC]�����h�f�׵��JÜ��-sD��q�S��Շ-H�ɓ��t��W�&p�:ɩN���Đ��>��G��~ԙS�\���#��*<M�����a����9dLû�7C�+���ی�&GՕ��<6���q���aaG����~�Y�z����-�>���YK�K�Ty��9�w�ԗ+cT�������>����?$��tN���ET���<��f�V��p�<�4н�*�����R�S��(#>m�W�n&_��J���N}����p��>�j�<ʻ&!��-U��#[k2�<Vʨ`S�7�z�b�o�.ə��D��
��ީg�U�Y�LaqGh��^�J�^�Q��wi�����h܌r$$�ӌ$��Y5��G/�%��w�_�����?3�����z���ɕ庄���Q0Pg.}�w��|������q��ۅL�fG��p�V��T�:98P�>�QlTʑ�.��aw���)��X������c�"����I�)2�A��!6�����~7��Yh�L�n%�\B4p�� ����Fd���1�G�A�ڸ�����݈K�:����Wr�z�=��{��AYՁ����i��Z�aԜ�Xܰ��ǜ���cf�lYGEfv��G���)�m�/��?�EX��+v�Tvz�����ޛ^�c���.�iy|�-͍@[��Rd��aT��]	�)��EG�o�
4���])h���+Y�<�s8��[GȊd���$�$3)]F���9ڼ�pJX�l�e��|h����O8f7��K=m�o�&�R����CW�H2��0��o����_����HbK������{q7��'�	14�U���^l |z����U��E�7�6�R���s�DB���F̾MS�H&̟$�'����q�3Z<�i�h�M��/9y0c���kN�@������u��@tQ�@�����f4�uO��Vy�R@Gq*��N�C�L�������%���hO0���pw��l��BN��t��n����0-��Sހzn�f�yb�����ә�r� T��N�ڨ�!=���L�\N}[]��Nݍ�L�}Q#��e�+�r%�2Mf�������y=`+t{	8
D­z֜�\F�X�q~L�������G���d�@�#�d��� ZST�}�Cf].;_���zI���Z akL$2�{������'��]ظC���tN����U�z��;0�hgl���
��j1�+>5֮#(�ȧ��u_c� ̔l�h��&�f�[+��`��/���5���bc����?��Z��$��L��*�Oe%[�t�+.Չ��Da:,����R&�Yr.Yq{2��A<}����y3G
�j&1�w���22ш)[��%&W���0L"c,�I1Z��O��i�:@����`��4E�C�۰�[OU<>_�O���	���=�o�X�lpA�E���vk�ʴ.��$Iw$[W�9�@-�� _��N;~hK�XE�D�����
�i�B��9������{_H�p<�i�ؙ0��ʣ���}[����25�ܛ�5�eiPj�vk�w$G{�{�w|�ͪ���[��s.�*l�:ޮ�t����O��-O����9�tfz�6#М%���q]mKC��Á�S�%H��Q��_w��:-2uӨ���� n/��2�*�5j9h9�|���-�y19�'py+3���.���p�(���}�NO@��`��Ċ ��y�y�A��H [���1�tNE+V��g��TD�f�����&[J��7f%U�Ycf>�.}�T�-G%�ѭ�q��"E��:3�pS��K!�E~�8ܨ����J������p/�B�ׂɺ�e����R®��{��E~|�߈��~I���\�Eԁ�bD�4�k�N�!4����������
�҃�8ӝ���b�����(�Fz��m�{QN
���TH�Ř��)J�׽ir��Ȅd�s�M�Ki�v�4�w�7���Hk�����H�A����{h��5���U��heҍ~����]L�J�o�<tx�  ����i��{�_��9���n4��v���(ĝS%7��?��B!ƛ�z�;�r-����=ٙ��;�x�zm��}[f�&{S������:�c��ϜCm����W�Q#x��
�ߌ�n܈��[7J����6|xV�����Y�K��s��{��0u��)*pN�}`2$���d�t9ty>��z�Y�rލ�*tU&����\�S��B*�7>O�
��/���ւ.��W�}�$�Ԯ�x��*]�q��d��r�n�~�<��,O�iVlp"�k���I����h�/'(�x'u��&�s�!��� S��[T��qRXt�v+oʘ�i��F���[:����P�0 BIW�����!�S����Ծ���u�Ҡ٥]&UUS�RɊ�[�c{�-k#��*ب� �s�����ʪ뀫����(16�\��y��y�N�7���&��i�ǅ���/�o_ ����Tڙ�H�+�S9�p�sѮ��U<聯�%`t�� !F���%��5zi�q�a��$�('b�g]z��'ƌ/���;����xK�M�5|�C���N{�$N��iH	n�nm��M�ҴN.�����0�}A�M�h��>2u�V��+���ς6-�i
rY��W���C�xf�'����o�OkU�/ٵ�U�I���q��S�D�D6�X�I��G�4��]*G2'ϑ�=��\S4%�:R�8�6_�E�M#2I�v�!(����(z-��;�n0�ƔT��P�؜Ԟ:�y�`K��+�J��$G�a���u���V�[��q7C
ݸ��\�RVF����� :PD��j.r�D%��V�[��s3�~1oDJ�G{
8g	���	�Kiv��D4-�w����AP��LoL����߷M�ⱥR]�I�8�xs�I�p�"8�s�O�3��	Du��C�X����1KF4z�o%<�i`�k=p+��M�V>�3NV��:Q+�
*|�X]MnxuU:��!��H`hǶ(#�a�$>�w���$G��Y��%L��.L�Eo���MU�����A,7ʄ0�+92�YQ�f�����8� �Mx�:4"������ڪ�ⶐBa��/c�le�����I�s<j�ʚ��S��ަ��N7kl����	6��+� #�Կ��[S� �kr�<�O'���B���9��[�۴Ib�Rz~Zo4S���}�򿲏?���T�U�ᾸUR����ZӲ=��/������$��p�(�9ՠ!�0�����`��*A�(�6�̠����k��d�
�NPη��:�h�IxV���X= ��`��S}|��{� M�g-����⽢� Hq�NOݍ,�}���7����6!�Td6�uekK7»�5��"0�T��X����y8�?t��O��c�(w��&���(G��P3[��{�Z�S��w��"'R����Xy}�Ӵ�㎔c�.��<`;���kG�~7Him�A��oR9�1r�����#���U� "}�tq=�#��Ŋ�Q4<���-08�����=�d��қ�"�<���8���k�SS�uΰy��!���a1x�-!����Q�l�����T��簋x�^ޔ���9`\�=d t�-�f+1�[<�џyR4� 2�;��"�iF�9������Wر��em#��zˁ!�7	�V�&�M�� ��(o��\��bφ���D��O�XX���ͦk�x�ݗ��,ʒ.�%D�=	$��t7�c��/�ɤq�����TE�\(li�ަ�w�aC�gc� P>��S�!��w�x�����`�����P�O�]\���� (O���,��$���k���%��崶��M�$9F���#>�<�<dNT,���-o4��j�1#@��!���_��Õ���ɨL�ֿ��;�x<�1֐��fy6C֌�����_ړB�Ƀ�O13��᠈ʀ���V�o��Q#)�-\���}H@w��+{cꎄ]y��c3R�0ϼ�=\�I
���3?�),��^|��:E���KjVB2��]�'_(A���x�9�N`�J�[qy3�*�����LP��f��@3m�w5ȶ*��C��
!6ҧB���+L� �α(PɄ~�q���g<��� ����-m��K�xmWǠ�s!���'},e(��˙G���ƞ}��Y�ɥ���9��޼D|�1i�����N'+BfE����-�"�Eu�ÆZV����T�՗�C��F��C`z���x�Ḡ�����&v�%�ʊ��ǈu�q S���$����\m����a��~-I��i탿�*��"GR<n��I����,�I������U�h�^���>d���j_�gYו��YB���ڶ��[+ֽ��בT�DqM�0��w��=9��n�����uK�����<(�*)�L��v$�I���Mu��:ن
�\F��g$3��T��u���%���02���[-/�9l����(0�k�W��e�;O�l!js�3Pqʧ=Zr/�_ܝ8|�&�	�G�N
֖\��(��{�ӣ��º���NB���Sx���6�7sD6P&�^�w���G��
C׹\m�x�ăc�#O���r��yHyv����_s��ŝ��-��c���8��^����@5a""�~�!{Ǝ�}B��s�(|Vc���r<ݘ�h��E�i������N��:���ף���.'!���0�{����v���I5��Ѥ��s��?��w5�+��
/��<�=3�>����^cvR��>	�.�� ��t!��͘a$�Mi�O����oE_o��W$dY�(x��|*���_��ې:!��^�e6X���}{A��M6��x����kKa�D�6m�ቂG��t���'���0VM���N���@L<������̝9vק�z ƹ�Z��,��lk&�V1&���RP v=��K߷rK861o�3�&��y���b�������F�)�Ke����H�&�Aԩ�L��Bh]�j��q
��>W��9�KyY�QU��[K�w�O����=#4�_�ةn� A��Є�d���&gh���~��
G9w8��,�C��m��h���
��_��x� ��!D5S���^^���'�ɭ�WءJU�){��5��P�*��ą��L�]� �Pnෆ%�O�$��*i��(G�q:��f,o|L��B����9y�w6�41Bs����a؜J���sm�y����GX��G^Q�Ȃ?AT��ĺ��#���.]����@�ι�r�1���zS7V=�)'�3V)�l1!��,/RN��Ƙ�<�t��Q��nBZv*��װ�����X��z����O���17�ʀ�D��Ի�3d� ��oV�k`��;աUP�s�ʼ�o�Y�n���\PiN�S��ܭ�:%+מ&��xp��唽�%�JB������U�0`��Y6@��C����1�.�=������Τ�K�	�:�k�Ȱ�Q��ir��m�7qD��I͔w(o�ʆz�w�.����S��Xz��e>���-�.�����<�!=��Ulj���U_��{Is�]���r���@ջ*;6�ӒJ�[���&��ۗ���H������d쩚N�M*����yQe�Y����.P�$�]ڿx$�J�+��I����I��iSW�m���G����u�#W��ӨÇ�Ve��kvbI�
F&���U�|2^x�>o\��bs2�2�)�H��/�̳� }�U��"�	��IPhck��j���Y�T�U�xt���ej�d��2��"�����[�!�'����eU֌�¢���
�����oÛ'�*�Yq��*�g^�'��K	-}m��X�B�f�m��.X<������N�)��b/^�0.f�4Ư���M_%y\����_J9v^����M�"|����
���Kg�p7i�C:�4�!d?��7.QV/fnX��)�2�gd(4\�e\riHB��˃_N{�ó�$K��P0���Ks����k��J�V��]�����$\��\�<�r~����S)��;�Kъ�2P��p��.dו�S6�x�g�U���Jj@�^(�t�8#:�{�'RJW�(�\����*V0
��Y�4��'b��i.ٺwA!�v=��и���d�l#�ň5�C+,e9 *S
ӌH�߁I�oww���_r�o4O]a�Ě����	Ry~H�&��R�7ka�o�O�
����.6U��&�_�4�����*Ω�����>5*g+�h�5hD�X����;��|[h����q�"�� ͗A�.yc�(Y��-
>$�l����3OΒ"<aU��Q��Q��2����YZ�Kn��lq6�ǂ,���<���6%w@=�уl�D�1�7+�k6yY�o�$�s���f�k��5gsX�;.`�����h�	���-�)�#{���vo��Sn�ks챈ޣ�_@9��YeHcr%6��xȈ�g3��d�������SYe,�bC���Y��b2|����U��O�Sz�SMx�A�Y]���sc���u7B\[��)X�[*��xA�4Y�����LV����Ց0�^�w;����7��B��n���7���?�8��6�,|[��UF��w܊4	=�ǽ��� �>U��F��i.h��̻�/����w0/����4���vR!G�z�o;�Q�eh�yq2�v6+
�R�:`n�Q<tP����+q��%��	���2�Ǐx�/~*VFsIِp#9=�ɚ�a�RP�8�.�S9Eb��e�-�U&�������1�o���P�9�/\?����	PDa&vI�L�n��\V�"R��7����<�,3zC̚��XxM_D�,����F`Cj�����Η���p<ϒx�M�>#^mV5���:�@�lH��5|�r�8��_ȅ��c���]0�>"V��Ƃ�sZF}|�u%϶��x�	�8,bV�����kM�6�A-?;U�Iv�4�P��gM�,b�wna��-����h�J�].ØH���I�gH�
�L"�C�j�1�G��ѱ`���������E��&V�"�Xy�d|0���[���(���n-]!mӦ�:`p9#�^�>��!CHJ������0��>�6�x3�w ��n'��t"���!S7?,�v�bn��e�s�78Ҳ�_��6��>D�ZlQޫ����Hb��u�����^�4����N�,���4�x��٭�4�Iy� �%7}ka���U���� ��I�jU�$�i	���֙zc)��\�jS�M�Q���;T�"�(c����!�z���r�[�7�=�R~�I��l���-���g���y��{{ٺƺ"PՒ�҃��8=��m����`�QN0cK�b �����*p�
���3��>���FE�e�:ghݜ?���k�|�=S��~�t/HY�&�+�[�ڞP���h����mAt�.X��V[��2��$�`.�t߹vKs �S�de�f5i�Ǥ��+����1f@�>��������]l��W�}�Z�!A�aAu�R:�P=1�� jL��`_[7&��Ɯ0�a}�[���+wv5:n��K�v˫x�
��?A+m�KRs��z�ň��#K�ug��-��~��d��`��KC���"e�yȼ�@ؗ��Դ��
�!��[�;�$���;~�v��3;z�f��%���������"�@Mv�V��|&��d��]Z��/��*H�G�D
J�������*{+�U��J���#/̅�6�c���!���	[���^5�ت(�{�ZO\��[l�6��pf(�PO�������N!���7\�q�@����Y@����d�f�v��]����l��w��ed�� ���N_���М�G�P���������6�.�	!,-4��iqU"S.�J|�"5�ژ-�XYġAs�y�ӌ��-w�!��Q$S��m���Ř�6�߂�V������<��f��:0��҈r���G�U�p*nv��8���g'hۦN����),z���dK�]ґ���8�2��K����k��I�^���U(���|S`�Vv"�t�ۄS��B���j�Y��Me��'D��ˁj�.MW��Xd�J�T MV�c�(�0F�`t�w=��=��	��.����5��rgyf)�t�������1P=A�v!�k��W�c�s֊~��K_�B��`*�^; �+^Jg�$�ˑ*dN�Ϸ6Ky�$Z��1�Wi�x��%�#w��$ju'CJK6����8%�u�����"Ŷ"���XY�WJK��9�� =�������L�3̜�fN0��@DPlʃV�xs�C.
��y�ږ�m�.H����`!�Ev![�ù����o��W�Q����K��E��eC+�J��@�C�`3�B@bj��d��t:�~I�@����jw?}���@~,07B���%\���(\'��l�]��4��q��Y���7�_����$w�ɼU5�%,��-a�� ��h���H��mD����;�\kK�n��Q��	e���������9�x9�{�&�[�[�R����X�oY~��ۋC���\�k0Jve,�7��� ����O�6u���%{ �ږS��|�U�B6�>%h����S ��&jj(���6gf���|=H�{�瑋̆�o���<7s�B�����%���xm<���v�TՅ��9*w��p�u4�#���q
���NX��HI�=$\�~rߙ��ə��~9n
��Zy��K�uV��0Zz��3�!!�-s��,RU���̰ih����`{$����j��^n������Ֆy�m��?A�����+� �
����V_o��ZK��"1�����Ԣ͒�^?�M<��V�Q-v\�α&�����8�Aٹ�' ��	�?��b��'!Ϲ!�ٽ�*����ǵv�>�ע��p?%1����:xq��_��|�[u�b('�uN���hT�����;��@����v�ލ�N��:�Ƹx��3���4j\�V�Sǆ������жk��U{�+ �/8��ml�����[�s_Ѧ/'�>l}z�n���,C���4K%��
����o����)N������q�ݎ�S�ݔ��[HW⎘6r+X���G��I"�M6���ɉ^���<M��$oES��QϺt�g :��-O�㎤a\�I���ˡӞ7z��6���<6|�MLOHB�����<z�
���c�?X����	�<���/0j��ͼm"�v��W�M_.|��-D��d�0�]��h��r�Rpr�o|�೻��HX�
 _��	�7�9�>֊��s�����z��c�V׫�K��K����o����~�B9��]�V��A�I"Cl۸����kw�"~8.��������ۉ�5d��ӽ_�y3Ľ�Q!��b����ݠ��Ώ׈����r=�D��Wذmª�n�cϛ�5��/�e
���k��~L���Z]%�bL!ݜ7a�/@l�'�@\C(�ϵ����@k9@�����.h��r���B��$i�j�+ի�]F
��Q/��S�ӨǱ"��j�ۅ1�Q�=홷-��a��a��	&����2p�F�)Y$��
L�QΚ��H�9�c�@�4OïZ^@�ef��������y��������I r$�VW!f�ڋe{D`��3L����=B�!��S���+1fU#�1bt> �V��op}kԞa��F�(������v6�KD�W�_X��ڰ�%�=�w�%yH��b��n������I���J��o2EZz$�gv�	<t�'��B�G��Q�Z�L[���%��W�y,�����p���HӨ��ِ��-'���4H,��^ԅc�	ȑ|���ne���g܌�����I ����t��zF��9oU���c0�v�m\Τ�����V���W=C@볓��c�E�Vv�V�H㢝��\p��q�a~T�,0�2L��L�T��r� �<��G������=��O��G�y:<>��s-�t甕�i2�^�m;7�
<�w`���EC���\�h��H*8�LD�U��ۘ�Sl4�NM�ZӽR�����Xtt�waog��"]Jz��8�Gz���1#��D���f�n"���p�MU-�PZ��tcA��/hM�f�P���D6���z3:G;l���n��j܎H�sB�!����f&m}�����!Բ��,�q���ձ��<5�[g�0��l��mj���>�`A��4H��lq.4,�A��]Y���L�x;���Z����Ə"�&����1C�hW��k�XN�%[��?�EY�TzU8�ĳ�i�ڄm
��z=���	ѐj[���Rv/&�ZR�W�F"����8)�K�eb�������2{�Y�1�N�-��u�I��V��~�5mDB��8@����)��G^�J �)��RM	�������#|wsB-�����J��v7&�^�T�r�}V��8��Q�Α����w�q�܊l�T|'a���b��f��Z���v�#��sK�U>�Uη6&�0޾-`���lo0�� Ct*��G�z�&���qMU����L頿<�'|�:d�hv׫�$�,:G-;{|�A��]|md�;�B�I�Z�[M�)潭��Y�/,}ۙ=�\�UZK��dO]��Z��.E�h72,�^�z��E�Φ_2KU3��қO��tX������g��~�/Iψ��P-&�Rg�=�ڬJz�����)B�N�e�RF�@XGi�.�%(���f��@��=e�4~ڷR�c^Gh�51D`��bE� ^Ug��o	���Ȭ�U����Wΐ�w�˾�q����Qj����A)<�+'E㭰b���nࣣ%�9��a�v���R_B��Y]V�HemƖӭC]�2�q��P;[Kn.���&�U+"�OX.�ʮ�{���4=^0��a�"*�U˞�94d�mvJ�A'=ᥪ�/�}��,�1�~	�<	b?x�bքܕheԀd��I���t=k���Ȥ�q}m�p�ז�=i�ѾOTO_�j:.��Չ���	 ��!����mw���Q��E��ǖ�.�=p1�˭Y)w�`W�~�w�䴉�#���E]���ɸ��5;�LvV��p���6T�Ϸ~[���g�(8H� r�Ao
��KDp]�!bH��.f~���j�	a�~,�'�M��*�S��#;�W�zֳ%���R	&^f�����̖b���ƙ6��U�]��_�q�fLDO�$5hn����:���ͳ4�Ln���6E�SC����g몡�O�
&3D�p�����y��)��l�ڊ�/T�ǖ�k��;8�2���D��4rP���9���6h&����u�yo�I��x�zXO��P�K���u�#g�;����j5��nY+�=��Y�wy+��n|;[P�j����M��Ԫ3yM&�MqI��>��5��֢Z�֥�f]_ο��j��p�?��1yCV�OSN��T�xHe�8G���vCrr{\Gn�a���'�;�L]�.@��Jy�XkS�L�{H���:	@���ߦ�R�w�4����ǂu(�RQ��ֽ����#��b5�ڻ�܋/N,�#V�x���U_昖R��̨��sT@���ϩ�}�b�d-9��l���h��M���)I�A�7;����{�n��-��$p��6VD��j�#�!qTH7�쌝�4i�SE��qzd�5�]��O�.hQ{vk�/�!$���$`-�g�& هP���:���d"0�y�P�N')�����	hxT��������4�}�@����O��j�^'�N:����{�=�e���aRvv�d�Ա�F`.�mP{X?ҹ���>~���;�o,!3�zd���`����W�[S_C�.�uG~��r���ᗘ�&u�a����>,:"�(�5"�� ��0H��>����H�ƸQ7tcG�*ť��`x���l��au�i��&�0���u��r:'ݹk����I�E��ψ��� ���B�E�r�R�ϩ�K'gi���¤�8��[�6�VD�a�Ž���^k,��E���֥�tr7M���a7�-q:�tRQ�$�����魙d�D��vi���Īװ��[�@��$y����V��Yp�p�8?5�뼶�F�6�Й����l5Ӊ���kA��\x��sm�#tx�,a�M��>�I�����pu ���.�L�1���kV�eؽm/o��^!ۺ�K����M�ɐ�G^w��i���Gp$q0���B-���b���1��K*LX5����5[HzqOd'[[b��Ȃ-̱͐b�� ��lu}�l�z�����i�o�Ռ�1�o�{0Cp�Q}�'GA�>C5�L�G��H@��r-���y`�0lZ���K�I�
]tف�.��cq����,vK��������܃_;k���C�;W%����RQ El|�b�,&f�,7��Op�e'+V"k�]��%n��|�i�wlLp�׬/@�� ��D�%4d����J$�Wm�v��@=0 /�|�E���U��)�7��dB2�4s{B����X�t��������4GM��7�0�o%��*����UB�����Jb�c�����7����!�9��:���'��
G*��&>t�.�	�V\�ڑ���&`׸FRA#[��vc�&�(��D�c�C��:h��#�ʖ(������A��fNw���?W�/��7�Xeb��T��B�tڱ�n3����'u���q{2%;;0�8=9����a߿��H����*�A4:�A1m����o�ĐY#�M4;��C���۸~D�UCg�:Dx�
�yr6`��:��tl�ٝX�6��}V���pf�u&Z!�B�<����8ɖ�@�j[�Y�+�8����Yb�7ߙ��d4<Xg�Q���'{1=�r�.%	������"�U�`�Z=�_Z4b��i�1��k�xP?@#�y W1�+r'~���ߒ��Q@���p��1]��%��C0����-0xə�������KǛ�O��~?d&�<r$�I�![���y�0���-��0����������׹�Z����=��l��5����D���,QV/���Ջ2�KZTD��[��BP�ؽ���XwM��V!�P1.W���VlE�Ul}�#G�x�D��௙�Xb2��%��`��3rاe�=X{9b3+��,m�-��މV0���#�����q�I�u%�/W?B4`7��G��;��oH�0�0e�എx�'*�Aˡɞ������I3�D3��R7wt�b����>Ǟ\����\쳽�dF�ǀH�_$�!W����-ϝkl�|޵�O2��\BC���&%ms���Hg�|S��/�8,&";�ji�H���B��c��r-�W������>��〡�~����FG �4��S�<0(��Fv��h6c��j~=��HEۗ�����g�޾�\�v���b����$wb?e�����-e��3Qc�=� qݸ�a�~�`�X)�#3� {&�����!�Pf¦KU��![��ͬ��>�ydSI��萢��ǧ5o*�!��!-��A�i��g��΂o���A�Q8�I��A55���cS~vQ���=SC��J���:������q�E !�Id[�Z3��y͋�Pˬ�l.x{�����D��v"�Dc�`��AV�l5����Ou�XTS�����Mρm��lt�\@�ڶB���������6�ݞ�J�r����U�pc��J���r]�ބ�$0��j?��j�'�r�Z #ğ|���2�_��n.c
�次�!CGH�<� �d}�9U@��x� k���e�_ї�h�#����h�(�ߏ��5=Ⱦ_��
�R�_�"7�	v��'���1I��)���	��Q!�#�֠f�!3Y*u%��`=�7�^}PR�܈��$���D�-���_����״����w�f������0J�E5?������ܪWk_e����e�9 �$��m�Ճ�A��ޖ��>6���E��8�3����iߦ�E90Sm�'�|�}�[��[ �?����od�s���,�im�F���E�����1��⎎��8%<-�u�Ti z�5TZ��~�&�!�L �(���0n��1�,<�}����+?�+����tղ�V��ݛ�'~��B��ϫ���`�G
0ɨ�W��	X����$�����a�\%�l�E^�s����nc<ćo{3���$Q'!�9c��_��:��(��Kev��'��z����e�ŉ�u�u{�:8�V��T1�V/2���;���B�����O�L3�OR�	zp����߄ǉ�C�F��{�,��iC�6���B+XS���(G��h�|M��䀵̸6��5x�ik�苋�|G��FIk.��w��\4�?�J��3��S�����G�i)���AL�k�u��O�r�i2j�Ѵ�����Hg���>)H��ulYe�O��OV��,�S�R�����z��D�o�;��Ə[$]��5��|�����8�!�v2^���T��}�RT�3��u�`����6t�$����O�f�r�Q��N��ڳQ=�Vw~�͊N&Vy>��|��7�B���Tm��7ug�#��r�����.�����|Eq]=��N{��K}����*u�?T��`4�yC�#�@�ʨ�)M���%Ć�~H��%5G��2��
�2�*�_?U�:�n�_Ap�����N|��Nʚ���������l�9P��*ۙ���wR�c]$ͼ`+8�%1�`��XpصY��o�W��[ ���owץ�����#l[x����_{��"+�����`t��8���H�W��g�$�	���|g�HF�>�Uu����Q�3���i��3�`��%9��й����M��=��l���<�)88(�Y@�c�z�ҙ��>��Κ�eA,�ƔL�{����v.t9a]�����iP�������5�URE���.���*���׆F	ÎTž���,���M���R$,�Y��Ҫ�EPȵT�$#�"�8�n���-�at��M��{�XT>��ʀ�g�Wc>I���C|���-������:�Xn#&��(�r�k�� tW�7eЏ˕�a�.Ǜ�!q	Z��x��q0-����CPE��Qq���M�t^�c�.1І��yc����Yݝ:�YbG�b`�YJk!7Q&Y��8�c����3��S3VP^��m������jL�M�q�	�|b�\3����v��}���WJ���e�UlR����:�qJ��_=�NǑb��D�p��1�B���]e�j�;@y`��fQ(:җ�]��� ��M�+ߕ���e��Тk�#0���c݇�QG�Pg1aEm-Ej<��0·qۓ�L��BO��gB(G}�Bl�( 	���f��a;H�`��Ω��`e����'�_�
�吹�����8T�N��D�����rJ���+��8.9%�9@�z+�9Y�O�'w�����}����vl�ј{��=jZRA��/��a���^kU�ޜ#��_[�7�k+e�WR�TI�ow������Yd����Q�����~&��hM���y�u$:ި��}0�2.��������٩�ʼu;�8�b������F=^1�V|v2犾��lw���c� �Jɳ�FA��PKR-r
�^\i�y�+/�G�ŷ$�p�w)E�P�'*黦�X�;a��#�F��`�.߾<׳ o����D`��b.�w^;�p9ݧd�+��^��_i�*���7�ǂ%{Beq����.{���ڼ���4�k�Dd�g^Z�->xE��|����������`��9������]Ӥ�R1�νh�v�G�:�@f)��A�lzʥy�Ĭ`.�{^eĲz#}�/֟w �ys{H����b q�ɀq��J��;CoE�G�Kn���i�D߽��������ג�FM=]�k�G	�QX�i5�P�&����w�$��s�4Trϣh�:\�{���B�Z��/I��D�m, ���K��7b݀�$&�?3���o	��1g4V�"z
������>���a���Q���V�.�@�V�1�pяf骶c�5ע����$�r/��t-e�B�\%��\�D��AϢ�J� �{	.K��D��q�#�*xb��Ρ�H��֔�NhU/��:-H?�]�P�<�l�R���*��2�m�A���wQ��dฟNA3"Ύ��M� �${t������RɩY9�N.�a�zmz��-u6YrD�nE1\�O���=\�?V�R���{���X0�I�>	��҆ߙ�'|����K�7�S7^y�
$�������A^�!����P�<E͐����VҠ��oF�-y��[A��w�sc�mPj���J̞�T_A!��P�q��s��Muf�W�e�������.r@��Q.��l=��4Ph�Q3'����X���=��e���%r	��YP����A(~O�m��w�q&te�B�����2d�x	��@$~|���_� @���-�"��q�������Mo�q�����n�)��o$y���'��%���� 8:�&����O�Q�W��	��UCEJG��F�VrXD���u�2��\ m�53$g,����T_q����īt��QB+8�;�8��6�I���U ��n�P^��L'د�b�W�`�+�t�Շ��
�Z�hOR��O�#o���Z���9c.�`X(������pQ�U�@��a��|l3���h9'�D���݋���a��^��x��G���K@�T��z���ς& �^�^�5F�8�fE=����R�:�ş�x$~%���bPt]߬�yT���9�x q�����qX��E-�J=t���(�&�9_�W�]kzQO>f���A���s֓���W�[�i�hDE[^y\䚒E�f�^����S�Ԡ.n����a�K)BA �9��H����:�B���"d/q�]�
S)Aj.���B�7=鹸�O�|�90���2�O���p]����� bG��i˻�(k���~�>�G��4��� ǋr<b�����圭��(F��ކq"u�s�!K�Z:ΪD�e�y
(��K��U1�J�����*���淊����OxI�˘�,� ��S݈<��޲m����Ǉ�4r3���@z�_����`���؍ a,W�>�|�׻2+���JL�!�,ٛݢ�ŗ�=}A�D�:;׫�r	.���qk5ڟ����<mw���hQ�\7a�A�Iv�3�|�"^=�D�Qs� �`Y#�	�niO���w�3�G�C.��aF<L�R�RNg�ynuo/z�屌�^�$b���T3��iP��0���5*.�}D1�����?�n�S���q��r���esR�-Ky�÷�EL��	��K�U�va񬴨��"	y7'Ԥ:8]X�?��."�?��f�b��[?��N"���z\��>o���lH��f����Mˁ�7ѯи���=K
��$U�m��Y�:�~D�~�)*��C��v)���������j\�[�ѩ�T�������gP��_}w�������L&죥����`��*7��g��b��§*+����^��ѭN����1��F��Ԏ%��M	����/���so��b"�L �|����XRO�LW��(��o���]�E>�[�b�<�#_J~�n�I����N��-��F�x.z�f�φ�!\�פ~��`\	���Q��fq�WOI����U� 2��~Z�\��Xӽ깅��L�r��:����:��sD�r0W T;q^.UƮi��ύ[��GNO�iu�"����Ϳ,/�~u��O�iNE����^������kf� t��I���L"p� =Q�ۓk��#� ��w��7UA�y���A�&�2w��vH3T���F	��ϩ�����9�iOV��Ғ��A?�PE�ײ���ʘ�t"]�M�
-S�64h�ƴ����st4�\�߭_���|�X��3�!#S��;Gr�����g���������&����M۷�'�=��2"�V�"�|���"v&be�N_�H��^w��s&v��6t��(뤞�i4G�=�GH�ö�4�tU�[����B�Y��sN���t�)������o��2��)ͺ�R�=0��L���.hR"ջ Z�,X�=G�K�`�ޔ�7ZȎ���'.�x���7�c<<���b��*�u�D2�b���ҁz� ���S�f��;���E7������t�1�E�ǟS��[��O��<n���Cxv��k2e�P��#�և�nw�W�g�LPPe����� �����r�#��A{bm�"�a5�'\�G>���+G�m�9��!�J�1�{c�Ģ�e,��y�N�\�=�#�DÃ�u�<�0�f�/'�ƍƼ���#s�-���o�-TF�l������b�Ś�r�~�-��n%��A���v Y���0�����R���`����_�kIH2�$*�lj&q���|��S�g�#@�Jv1��F|���'�ѹ=铠�~#�q�� ?3 c*����P̜�G禍C��K:.m�<=�sW�ޚE�Nt���n!�K�$.���0_c�a*�{��%j!aT�t͑M���$5ĳ�p	����/_�,� ���t�k0�3)��߆����<�~6�S������:�X��GP�M�K�{͗�e�lj�� w}���/�g��J�s��:C,�&�F?��.p�,�U�
_�!�ܙraq�)�H��8�gl���,�4� ���^ol��e)wU���)񜣲L���ZT�y�O�@�w~��S��9�I�@�w�ֺ���ں`F{����q�ɺ��-=w�8~�.�*1�O}Q�)L��m@��I��N�4�z�e_Q�P��"i�7�zA���K��W\�|�[�~Pݣv���1`bf�e�۩�a^M��^����G���z��(ّ��&����F{jt�+N0���2�%�{6��8[�Q���8�)kK�~�[4jkؗLЏF�)z���$,ϸ�7���k\�1k�z�~�zN��y���8A�eH���Q���
��&����:��yʐ���&���tИ3�$[s�N�.���:��S5��
�1�*�H8~B�{"-ܾ̕M2�ݼ9黻� s� CO���}`4�(B�o1U� � hh���16���3�v�1WŔ)��hZ�l74nd�I?Y�7�J,*��HW�[?GR���#�6��Q;���=�d��)r�$E��^�t���7��o	������$�!}��:��}��Z��.m--LK�ߑ�?w�z8~�e��Z���\"p�REJZ�W��k��PcǢb��x��=���s���:�x1��Bw�����y��0��e����yp�qv�z��6쾘=wW�qՇ��>Q6�|e��Te'�R���}8���B���m���g�cx�S��Mv�(��{����V~��ˑon�~�������Xe4�de�i}wq;z?�(�f���%ձݠYd/�-{sj��-5N������"Ki_K�q�Hnb���z��$���s@o�G� �M��G��.brbZZ_>��ă����hcK������e��<(�՚h)��̳^�M���
�����|fH�^�咀C�&79S��K��t�?W&:�41#�ab0}oD#t��h�1�����L1���k�����a�A&0�2�)�9�ɗ�=��ًk��.�W �w�s� �P���ϐǲ0��Hg����65��~��Åzez���bݶ��cHA���5}X�z�u^h�=�[��(�n HO�s��U��8���h��7���A��$έ@��4<N��J� �Ǩ�q�#R�,=��Jȓ����Z����E�Io�c{�I+����z�_t\1��:/�J39��CY��B@�N�2�E���	�sj!i^׋,������0�8zUxVZ�A�4ה)���^���n;���/U.����ҷ�W4ߏש���b��+�~#S'����Nm� ZvN����}��=�y�{N+��0,1ω���N}��)S�L�oՃ��1��R�6L�~cG���zڎl$ ew��Jk�
�b��2�Ҿ0�����ѽn|FA��矸��~3l˩�)Ծ��m��m��u�%W<����,�V�����N�˶'>R+��MO���[c�Kn�e��`%dr�nĔd..��zBe�K����"35�&�}��è����R�Wbݖ�]�g7�:���6Q�b�U��?��϶j��L�x�om�!W�o��YU��S�f��`!�*�8�v�2X�ذ�3��啛2x'�ѵ� �-Z���S@�b�(�x��5�-��}^"����æ�3bL�`*��U���� �F	��yNmN���k�ݐ���{˾�Yj"}���R�����&^���Y"��3�T�5S�4��І�-9ni���.�[�ApI��b����P���R'���݋�j�.l�>=��:@����`�k�㘱_a�t9��:����_��s_���Ϗ����Y^a���[*M��Z�aۓ��M������i�1�]�/)�u$�������8�FO���"̓��,�7��|~�Br���.���ݴ ,Rˢ��@��T,�ƍ���L�����5�x� �P�\0���¥�8Y7��g�8��CIr�Om�՞���s�� ��qa
������Qh��+v��QqNr���<`�{�Β0�Vp0E#�vp ���$B7d��&F�D�.�-)HD�ĄRR.������q�U�b­�&bҟS6�d�?u�n��/q�gl�3�
:��h�H-�.寜&��܅{n",��0��Г.7�J�3"�91��t��]�Y���1ܢ�̘�W��>iG��R�1k�ԥ=�o���#��k���&���!��G�ϟ��۶4��8� ���TT+��P6��E"���-i)ޥþ�V��٭�j&�X?�ܦ1��F�����7�4ݡ��R��k����g��WM���n&���M�3���H���9�[�3'}�^�Wn1R1&C�e���|�,3c¸$�C����*������e<�w8��kVkg�{�N�h0�%YעB��ό,!)�
�em˝��խ�'���S�f�-[7�AGx�X������:�)�M ���2b�)&1
n\t�/����=t���m�x8Ӄ�&�k?�q ��o���^I7pV�F�͞�ݴl*�W�#�0�6pK�y�Ș@r��q+�s��<��%�"}�>� ��t�լ�M�\��W�x�-�`#�t�cJ���H^�+�8�� Jc����t�2��e����~d�r�ĩ�?g1�
����M�$�|	� ��]{r����c��F`R�,\m�
�P���?�l�A����4>"?��`�ق;s�����A"[ٶĸ]d'L���=AU�8���j�����y�CmS�_oy��w!��-�����B6]N���=H�F�.��]��Ì�'`SF<ɤ�{�6Cz��Cm�0��x5�׆g%�@}�"��:��+�\$�)��u�1O ����b�2AǦ_9�F�����bn�B��FUN��`��&��[5x��Ǻ0���Ø' |����k�#Y-8�SYE���A����� ���҂�b�� 	�g,ɂd���	���{���0s�o��^�Y䑈��f�v��1 par6�牏ɤ�R/�dhs����鐾�U3_kX)\k{-Yl^�!8}�rj�07������̞\S��O�f�N|�g�.D���'Z&��$$n�!>�,�p�� �Ŵ1k���c�đЍ�]���-m ���}
ʿx�~��2�a;��ZZA��
�a��rE�]!�UB�~Iq�ȼ�Z�D~�e㺿�����ۦ�Pˠ��:��/����đ�����B�W͘lw�w�/!�,���ڃyhn�6�A�~5�o�h_���N!MJ^��K�顥=��xR��'��=B�Lj�q��>��Z��W᜜x9Ȝ��-;ʤ��R��;�UHɿ͔�}�C�wԷ�����H%�]�p�,^)d��	q��c#�I��ΣWɥ��y����͏n�<:�+�܇-/�X�)��O�=E�����6q5uсگl���a�	��n�e���g/|�;�0�k��LX�>� ���8[��`�`^�S�ɽ��'��i���StD�;�}���ׯ'��%7mB�u��s&A��:��CES����*V�ΊM���+4��8$�j���I������m7#�K|�=z�x��h��V	�V���IE*��A�\8G���Ƀr}���-���c������]Kh�L����(�IHg���i�˴���c�-��瑃���n�k�֏�GF��H�ܝ��x��*C��N�8]&��h}�I;�A6�N���d��)�a�����ȱ�'7�2y�����)g��ݷrJ����.��/�-y�P�	Kt�I��L/��Q�f�]����}�L�����\q�%���s2�:W_���������mS1 �̏�6�ju�{���ɱw��I�,{�n����9ܙ�t'��ƣ:���n||L������%�����\�����3^�TQP�,��|p�d���B�Ɖ��=R��Qi�+5J��Q�fW0J!.�a6)��^��2��L��_h\6�����/�ε�)Bb]a[^�{�B����9�b@��U���)��zG�D�#���*�������)��V@ZU����fIʧ~��nP袳X��_R/&�t��.>re$�H�4��Io��B�NN�+���&ժX�rW�""l�amXm>?=�do�� �|N@�L�:,��!�ԃ���:�X����B|�䖂[���ά�r6�: w?O���(W����#ۓ��N�<����@e>����N��R$M�,ْ�����E�>�=�L]����Ԯ�JSQ�7g9����T����!�f̞W���Ǹ}��
�ƯWl-[������ޒ�}/�k�~�:��0c�BE�Ub\�JM��l$n��:( ��J@&E���	�mN3�����!�k���a�v�W1X��Fp���q�,R��f!l$8\���0��%�^.d�L��4�e��;�|�HsÈ�1�&ϫޗѽ�ic�dj1�*���t<�6�-qHӽ�R�D�_2���JْBx��LqZ.�L���d����Z�Il���6ߜ�b�=���g,�#�1hY���魛�Ti�||r*�B�^.p1",d`���,p?�E��!t��}�o^�H�^�MY�D'��C193������P�]]�B9?�H����z���v�VD P�1H ���ҵ�ή٢��17��bH��&��<q����e�"���z���Hk.�(>4D��a�K}��=&	�'�u��i�"��O�v��&���-쾀t�vr�L�l�W,)j'Z�OF�[�.P��;�rrk�Z�{����+��F0��hzX��ԮX����s2��|�s)p��X��}t�<ed��V��PrΑU��l3�؃��4&ᅅ|V�G��*ZZ}=�_��
e�vG�!#.cEb�4{�8���h����Ӷ�u�����y�i��!}�Lf�1߇Д�.�Y�Yڿ�~R��	^�@����Y����&��'����B��,O|D���ew#�34��h,B��[���`3�=9]Ny9��{%l��;k'��@��+)?-��!��H�Ә,���-�g�:��ry��ɮ��yeg҈����	հ�A�h���1�1��?TP��w:I���y=��99�-~V�.RA��3[W���^���I�Vd+�D������$q0+)LI~�-LC�Q-�<�M�
V��kVCL�:�P$��_�!&oPa؆������8���j����l�v��.-���.��k��B~�[&G�W���G�e%���lv���5��"�6���![�ucjgh��uƏ�m�.�alw��s���:zY��Ak���wH�wm�<"�.��Ո<��S�U�>uq������p*�X�Qd�t[�Y������o��R�h�5[�Ѡ�_�9X�a=y/i��=��A��S���Ʈ"��*�$G���j*m�����u�֌�M���DF���(M������8�/�OA��r|��;�����L�Dr��sOA%i�ʚ���(��s,�d�߫5��~���fu;�qxoF����Z�7�b/��М��"�t]������k��F��7${��]Ea�p�b��U��a�3GI������*P��p�*5�6HŃ(���A��BB_]'����z�?ǹ�+"y+��0�vm��������R�kdFToȫ�UY3��^�
%n�['�|^ f�j4�{~Ѣ�Q�򏹕B���	�xD�����@h}����N�m��=F���R��<X�u'3���=��u�a�Z�*Ӷ���gؔ2��(�P<'�svj�@��%=[�.u�#��2z�t1��5�U+s;��7�vڵ�r{^�ӑ��es���z��A&�����v"�Q�&�m�Bm�m���l� X��NE��k�6P�R��O�մ�[H��JEYQ��N��6�����M}�	Q��@�od�tr9��tQ���<��~�
xj�Iҽ� � ���j�ݏc�VxNcxW����wL3���
��Q埀 L�Q��s��� ���E� c��� ��9&(����$���F�;]�nl���%/?����o0�2
�J����~�j�@w�1�gY����<�|��<�PM���V5Yv0�G���{�-�B�6#���;w�]�fk���|`:�	֕�{��l�e��U�e�Ch�V�%h���QB��p&��P����� >��ŕ#���ڨ�W�ER犛�I�f���{M��4����/'|���)���Z�ͽ�u9�D;��z����9���eTl��T�Z=Gʻ_����'k?�(.��f�P[o5)yS���$���^�yM�*5v����"��k�~�@ѲF��x�f�C.�����9Z�ԓ��)rj�����^"��&d�tkv"w�L��o"Sj����Br�x����:��q8���V���S��1�i��,��o��9�e��Hg7ki��o�(#$ձ�!R�$(�t5�.�L�l��\+3�}�ےk����?��IѬ�}Z5���'���lZϏX�mII,��C��iBX��AS�=1�$D8J"�6B��EF�!oYT|_΃�8+f9��|�ì���쬜u������:��5��*w�i��E6��V�<A�lD����:��~'a�ƀ$ۮ�%�ҷ$���±D��so���1�]�X��e�V�&�C�apG:!��5X���\$3[��K	��!g_����?����)��<%�����S:��Lqr�~�$��������򛢎P��y>�l@i�2�Ag���.I�r8?�҈xl�2�[Y�!�۲I�,+{b͕�3��(,�,A9`$����*^]��u!=y�rh��~d�o�S� ���Y�����?�KJa�9��5&����#�`gyp���|�<�h/C��\;-���
�\:��k vރ?��2��Ъ�@��x�j�t;�D�X�����!�4T�h �ճc5�-f&}ST'(p^����_ ��ç�cCH�dA͒�Ϻ����՛-/oÝ���h��%�W���>p�Jg�t�2���,�i3��J�}RE������3/c�ՖH�;-�1�r���5�dK�l�� �\��K#��(�����"7��y�0fL�5�X^'�D�/��c�d��،�$�NЯk<�_"��Z����eYA�-�J��b
����H�08� � 9���3�����6E�@ �c��� ���mS�:O����G<�HR�p���1^�Sil��^ď�=�q����j��vs����/$G\�	J�R�y篦�zy��h�V����!~j�QiZ_���ED��ڕ�75�Ţ5g�D���%�[���h��$m���R��U����UP@����!#�H�t������iK��d��>R���K=\����rO5|�\�\9���+L������ڎ�j��YB�+ �"@z�ǂI�r�IЊcEz�W}B�;��B�<����A�H�w�J�|I�@a�&��P:�U xj�K�$m��8-��>ߥ�(���Q覒�פ$ueәV���U-���Q�O2^ ��o}�F���U|�"����D2�|5�u$7����;��ڞ������f��J}N� �NJ�4�Fυ���"�*��UUQ���������#Y+y�?�@�*ހ�������9PR�z��ո���6�RY��߅7��޶$ڪih�kC/f�O������m6�L�gG۷c����Or�?�0P�#l�K� ��ZĘ���yr���)-9:G����/��G��>uz)"�û�s���~�*���&��H�Ft4 {��v����"�0г<�AE��W���?��~1�c�Y�83N/���!(�e��J8$n@��z|���mI#��wP_�HOy<6��O�ek�i��ד��9������
&�>�,����N(A���
:��d%}�����
�f1B�&?�V�Mg5*g�#�;����̺��2$	�9w��\{ҍ� �����U�K���������3x��קy�_��I�����}��hg���Y�_����&-���|\)E��|�Tկ�ғ�\��
2��s�1+��j���D4#̲3u�LS���}�cHd��B��?��g+P�c6��H��lP��6� h]���_�#fO���g�z�'��?@��zD�K�iv�\P�W` �v>
G�Խ����Av��}���R�**���v.�N�ϳ���;�L�т�����%�;��_m��ߩ��'-&��Ř2�q2�Q Y�)u^��nQzi�d�.�kЄ줅
���c/�Xɘ���Z��+ ��D*�u�ӕ\�'��� 	���Gm��6�?�==�U�ꘞo˴ʲ�X躐B�Ʉ�]\c�1+�O�m���6�8`}tYk�P��Y�Z[�k)��d�2_b]�ue�̃U����o`������h!�8�pΎH����]4�<�Ε�,���?;��J92n+5��ކ�X�������*��KH9��������ݨ�td<�S���SJN.�oKHk���l�-����e��@�E���P�F7���'�#:�^�M\ܻ/#}�y�!���e�X��Y����pn�4��f"r˂.ek~��$!���w��J�G�oa
`��!�BT�����^��VP����B4g�ħy�zQ'҄��I����u�d@H�P:n�I~X����~.� ���篩V�>
Oq�#�	�\��ծ��׿�*���RM�*M�Zo'P���x�a䷞\�oB��5Mca�68ӡK3O���?�*��ν4��2��{IUI������B�y���z[<bTnL���;t��q����t����~�O��2�y�DG � E�h����o��*�K�_-�6���Sd��,��
��2ȫ���=V�/68FbmHs�湂���j6ٝ���F������a=��r�i���i�K�D��e~���?֡�OL����6��nv��N "���Z��U.�wsWG��M���.��9���Έb�.G�6+���K�.i�� @
�a�hu�*�H�V������ ��fR��2o�sexZ.W!ӹ�X<o�ӏ�n�4J�ӽ��D������k]�G�)M��R|"��mL������Eh�n�{�:xT���R�-l���Ny`�m7)�)ֳ����}��8��.�``�Ǭ�_�o�:����4��t��Z�_$���o�L�zE�r���f[�m� cn 1��v�=g�+�O���e<��Y�D�&�<�7@��(�8�#��'D�=rAY.���j�I=7Vo2�b�Ĵ��>���k��8i�.O�R�eqŘ�7�kۙ�]&$*'�â��v7�*L�=퍡d�"��{{Tӑ�tL�͘�O�C������:�f@�����_Y�;'g�(�$�{wE5��q����q��">0Ks��?5�ڏX���{�r-p��:e�__���D����ْEI�ங�K,o`���M�z�V��O:���6U ���.�f�����I�3��_�+����Z�mx���AP\v�9<�@�X��>dq��e���\+��N��2/���I$[a�z��b�[,���E��v�3�Pk*�vMޫ��s��O{�8Θ���UjX2�9Z"��r�7�N&uȡ[4wa�LѮ헆(���O�-����Sp��ٴ��?��(V�x��*Wr�:s�/�ԇ��@O+U���T�.v�>�|�"r"��f7�	����5�3i�������He�h����g���L��.�F����cd� �[s�Y��J6:�t/� X**y�/D�	H�P����6)�d�0˩�J��x��s��J�+�c�ci��ٮ��<�_3���[�}�=h��MP�`o�u�j���o�R�G�o�^�c_YW>M`�%|�5��LR�0t��JX�v�v�OaaO�����d	ˣ|&d���<RD���U�>����(̒`6P
��C�չ='}��o��!0�H���	���~r��qܞ�ُ����)��,��.$+�8��A��ߖ���v�37�]�c�Ty�r����x._3Xz��y�V�s�6P݂�R�լ8an�/9t>5_4�AC�8\~���E�뵃��O��1�;<Ie�9k���j�'�b:�|�Ћ�g4��v�\���%����gI���M�ꚋ��.�P�u ����݌�9�b+N�R�5�=��if_�υK��b�B/��v�Ib�(�@����>���L���?�{�A[\��P7h���f2��#D!��Ҡ��xZJ
�4�/���Q����j0X�(���z�X{)�Wq�F�!���⸿��������S~���`149JL Nd^����R�������rk.�*=����1bF�;k
k�x���p{`�P���~�:��4W�{.GC�ޱ�٪kZ��#�r��D��M��9+̛����]p_zvԫo9�;&#�YD���5��W�l&���pzx�o�u�`#\N��<OX��UrX��!�/��_�w���°�7���
�;�'C7��VmcL��:�e��Q!�#!�.B��:G�p&!?>�N��.��mʼ���8��~i#�t�@�����[�`S�3T��푾���R���>�U��x,��f�C^L��0�\d�+\w�2e�TT�o�m$F�_�z�Yz&�q���+ Á �F�|�R`[�6�!:ᖚ�7ݪ4��*W��]��o��c��T0=O�w9&��n���L�(��\�ktL�*#�k^�aV]�����o���J�2�ړ�p�n�⮪Z�2}t�o��"~����^X��q��S1^�7RF xkxn�m.Lr'��W0>?*,f��βF�2�c��Hw2W
bVW�G7"z�ī�HZ������:m=iZȚH��r���k!
*�\c��-k.�;��8��뱜�w�����l&�n5~<4o��ol>7S껖%�ЛT��8��u��'��e���p���wV�V�X�	�j�4�?��Aw�hY��.��0K�$��h�-�� �G��;(��~�*Pח�¤c�En��>��=�8'�B��_}*�Bl1ͩ|"�PW�Ο����,jf!۬#�U�^�NK�t�NL�:up����e�&A���gN(�8���"j�@�{����Z�����G��A�(p_�d�VeBõ�~���ۜ��d)̂�H:OP4��!F�w|
lOպ�փA�4keS)���ho.e��oAr�n����������2��?/ ����RC*�P��!�$����!���r!^�2�]�U����*]��Pj"2
|��`�8��6}�u.�Ͻ�8��e��1.�;�m�@w+��p3Lϼ%�2�:)u[�r�M�Ct��Ě��VhT�uPtx��!Y(<��O���s�!�آ�N@hb����q��Kw�A�^��ziE!�cL��f��YN̩�ؒ�V�'uG,~�8�XFn�@���`��BH�Y��x�r�N^M���']���
���:?���=slaھ��x&�*��k�'n��xi�]:7�(�AB��H��S��A7�L���w��I�7�����	�T:q|/�8����,�bt��M}�/��b��0���E� ����J�	�ȧ�1}�A%g���'�� Ťʾ$��ϐ�2����s��D��^����wܲ'����#�b���hx����Q�)��+뙳F����F��a�I�I�XP�ǹ�='���Ȃ�Q���F�o�,ƌ�T �rV̕A=Ka��pi���f8q��i�Vf��=���#_�QZF%Y�5��R���_$�.�OL,�����ܼԵ���"�/��2㟩��zPt�����cvǑ�uN8~���x�K�eו5��@G١�E���W1���U)c$4�v�9׏���&�mIz��.H\�ԧ]XFbB��i�:�+G�1�D0�e,܌��d96D׆�)"��s�+��SI�wz6pC�aX��|>��hc���s5�&�8��Pg��	�_א�S�����}>��yy�0��ձ��J��r��3���M��(��G��ǍfW<Cj�C`��@���0E�����r%��g���SQ/hk�n�����s�e��]*}�`�W[�������#��Q���t|���`����G��ZL�UD��ڜrMK�q�rtr�)�W!%s	}$V�5��4�=I<;�u���L����v�/�W�OB����Lq����}�ΰ��¡�cK�7����#VOj#7@E"�6LY���@K���9;���'P��x�3���J+��kqatdë��e[X��hD�|+��1H�g��q�i>���k#9�pUV�Ɇ)�2E(L�Y_
��˫�(��~z&���T�i�-Z���ق��{s����֏�o�C��.��{���p��[���>���ls�i�lGd�a�,K[���\��m6
L�(����tx��7s�/y�;j�/��U�篋���m���0'��|�7������`ꗦ��8m�S1��ɕ�ud�t����	�>��H�Xm�\Z���?YOb@��~��"�$�ƍ��^k�7���lA>ZU�刯T�s�x�l a��_��
9���VG� �(A_Ȩ"�f�W꺵���ܣ��Qvl,߃�d���W�Aj�6V�2��o��S8 ��1�I���ɰ'Z4MX�e(?F�D�svzp�!�OC�f����ax�T[��DeȘv�!��rZ�ǐC��x�jG�Z��5�߳��d��)��܄�;�s���{���Tݔ+ɹלL ��]A4�Ŝۛ�mh!�tf�e:��?����)}
z�0���4�rR�^�/W�� ?]Z�boA�.B�H�!S���%�焚�54e~_���:-�����E��l=�
�&�Q{���������"jb;�7�~�3?╾�.���|�f�)9=2�3�Ϗ��#B�l�_3Z�6Q{V�ps�xIH6�$��>@�Ӽ2 ��3|vbk&�Yݦ"�bk��н�a��yG��
����Kh������q=j_Da]�����z�,���0�/	wq����B��=9٫Ě7yF�6~ \e�e��cVwp�w9T�Y'�F�&�	6�VY����Z����[#��@�o_ܤ8mM`B��C<��{��.�1�@0��4���}y$���؊(g������W"��%���5+�($�}(zݷ�\8[ ���[�9���,0�B��k�L�O(4�9�E���s;��J�����bp��	����u��qtD77��+��Vi*,t{˧�\z�?z�C�N�����`��|?�ӗ�jR�#�i^"uc�R^��M1���^�(uz��Ŵu�N(�+H��Ϥ�Jk��
�ߤs:�wUn�z:b���<��T�Z�;=������Р���W�5䀻"�&�~���5V*�sx>)���L,]���I.��O2��6g�9,�n�G�%�*������Ehҡ�K���颐<�̿@E�F�Sf��ݓi�W@:M�
�5!�k$j�7�O�t�G�v6r��ĩn����=1	���>��O�h$� �0���3��t��k���V��B�ei��hm(Ǒ��S�bRA���!����"<�zN��	3�o�����&f��S{����>�/�6�l�̞�R%d[eZ��6�z�p7|y {N����9qi��c���}Q��F�� 
y�x�A��>9��+�I��gٞ��ğ?����)�~�6��x���D���*{��kxu~?� \�Y�Kx�'�F��X|�3���C�����mf�ˀ�sΘ&��G�3��S�g�tH�����H��l�P՞,��|�̱�vl�wtwي�<8"by�3Hb'�Q��J�(��=��=X�����<mʖ��i����t<�����p�VZ���LB��ґ{�9(�`�e�y���� :�9s�����u�c�8P)2�����rc������ѵ�%ʧ!�Gʭj=;�	�yOR!�eV4��w&�6Q��5���u^���]��Q)���l!��&f�enE�f�����"vI��d�{/�t���E��3�ž��|�g�2b�.e�\p������GPQ�z���'��h���G]�=n>h��%:�^�l��9�Ǉ7�^j�K�,u����YZr�$�D�`�'Dp��#%S[T.1��WL~\,_?������D2C�r�"ӌ})�,t�=~���;�L����U7?,���v�|x�9�<}ʵ2�B�U@O*�#ʕ��+�t4��=�T�kc�Sc���$'o�p�b�z��<cK�/9j�vK��U3�SAfK2*�tI��Z=��@֩_�P�As-YĚj��0��Wq�U�+��F�IYI�|��}�������izg�Ѿ�VI�vx���c¬'U�3kr3""d͏�.�zp��MIf1�O�'y�+
[�᚟�(����'���$������1�8�r��C9��-�4��n��q���Hm�!���������c��`�6�#l���TK$5��C4��,oa������O��i�_DݚM"9��[4�� M��[ZK�mG,����������^%^�/5�!��i?-&Gq[�Z��S� }�����p!Y�U˃�/��� �DS��f}�#�̶x�C,V���r�r�j�jz�z��&�[�(�6���-�o�Se�S���!��w�*��v��K�xid�y�.�`��A2��CgT@���b�ό愇�)��W�퀒'2s��.���q���Vy$-�p�R���;?ٖ˵.�d?��ޢ����i�n��E)���˛	񡧁���^`�ߴ/~Lo/�G�����g���Y1���Օ������*9@�FZ��,8�)q7�?��ֶt���H�~�#Roj= ����{�ǯ�7X�j�^-�-O�0�G�KȤ�4��J���4Q�nv��̳�X:����֑��EN� �O7�r�v�k���|.N�Lm&��oq���u[�qᗾ��Aȳiwz�U�G��3=!+���(8E�z3c�����fC�r@����m��������"�ս��#�Ga���,XU�����ҷ�'���"�j�~漭�h�O��1C�P���(�cLv� �ꆱ�
�0�M��Eҵ|��x�PwYȵn��� �1u�
jj.���	N���P�έ`\����1�k`)�5-`�y����#W�\\�I����ݎ 뎗�M#�~~���*C��b���Z\����Q��jW��rka���O�i
[���>���{�� 6p���0�Vm��(FA�-N0X֮��tI��t7ǡL����~Y��=b[�RD^B����`V�ra����X�4`�"��k
"��\
��J�v*���9nj�d�Z���a;[�۾q�(Xi`ޗ z@��D�ӂ���[�"��8q�\x~X���,��z\�&�3��p!t��=,>8X��Б��&�s����O��n�Zg��M��F�ZpcI5@�e4�˶?�y��h�';�,�^�8,u��3�x�a�dL�דG/�Ff����KsP�C�	�^��5��:Ϯr��J�_�P@��p|��͘k��ƻ(�;�"f=��8���?��@����/�Fe��񙮩�K�wn��D��Y��8C�T�>�]��6BuZdZ�H����J����鏨���w"h�r��%:�3q�0�%�㴸��0�w)̶��'���Z�}�7�ZK�o��
��˓���:c�n�(b�~������t(�@�w�����ڴ�٬��׳��=�Z�2���Ɉsi�y\E�Y�7L:���N���@
�2xE���V,��PY��Bf�#���Y����.��C�Q��������QXg�=>��~�t@1����g�� �����(O'�D5=��	��J��>���]XƧ��,ó�߇��8W���|i��VFi�)�W��ܓZ�����g�\ �>;Q׊<x�#�3�F��W�u�dx[�i��͍Hɒ�O�w$������$�m%de�*�+m=dfE���Q����]�X��F���,�y&����a,�̢��wy$8��l����?F@��4SK˭���%��x ����t���A������6��V�QC�{6�k�N�?��� 飚PQL�)���l����U ���.v�\��R�t� ����f�h��V�,m��M9J/��l!g�s�RT������G�z	K؛��fA�����]���=TI,�vH>A2\C��ǘY��Ǹ�i��#�E����hӐaU�㴎bV�P�m"��Z+���!��`{u֑��(r��+9lo��{}Z�û�R^^D�Vz�!$O@J�du�HAQ�����Y�����P$��r�5�Hp^D�o�g�2��JR�W3�Q@��Cje*�LWG���m��^ ��I� ����%�5�X=拲�o~�E��1p/3d�2����� ���r&��6}����0�pf)x���������0;]KH~s��>n.�N����Lr6�"�	q��fF�ȁv��_՘�O)��f4������i����i����J\K�8t�Еa���@�QRe�	RU\��~9|C�F@���w{:��	� ���`{%0[���ED��d�J��獪�o�@~��]�9v}v�LLs%D�;�ϱ��-�q�'��*ñ��!��~��V�s��ݓĵ!@����3�Sɜ�֋��Hҥ�d��L8h1X3�{sN�N��i�x��T�󬕹���t���lW���������HM�V��"%]o=fC,v�X@K����_o`�`���%�����+�@4���M���E�	�1�MM�o�,��e�UUji����0#A����kvM�?��0�F&�R�C����d\z��B�8��+�|j���*F>�8�w��.�|������$Q�3*!�_�6&Fso^^AA���x/������j[KD�7��b��_�1fa���@z��Jo�dׁ�rX�t�~����Ls9r?_ؾ�����EN�05��e�&L�IQ�����Uǂ���N�Lo��sM���������_ִ����(:�ɷ�+�{p�ti;G؉���e�jBJ*����$�҂������]���/8¯l��܏����.�]@����N��*���;0�6��1j2�� �a�g>�1��ؙ͢�h�T�A��P:�����P����DnX}WOCq*�7X�Y�'���z�
�q\�/x� 6�;�+|;iv�M@�Ȑ��H08b��	u��NƨKݐ�a�1� ��X~tTxWr����:��c�6���jL��k�B�$�ϊ�G"��q�$��qm����ǭ ���n9"�^� R�g�+��fyt�'�x`�Ā�*"�`�[%�Ps�
�l��M���C^���t�^����i���'�2.zSc6���ff�/�an�T���������L���ϝ:�l�{���pu�U�n���3��\�o��7���)g�c�K��Kn��d���� p�w�|�&'�k���-g�3E�%� հ��@�$24I%M�W>I7��r�_f�F�q$�㓎y����y=`d�%���︂ �;q��B�#6�LPw�:es�},��� c4x��6	�o��*��j|E	�Q����_��!9\t�s�r�J��M®���֝� E
j�yQ�G	�	��c�:�+���Z3�K��L�r�� UUb*=#k��U$�!;�wꈟ�ئ;w��9m��*��>�;����N�;��m>S���?8�_\C��|��i�rUb�쁐�p�퍮����x��=!�f]ϳ��*�o�!c���5�ن�2��/�E��������M�i��3�>�$֠F�2mexR������%�X&:WU9���;a�ՠ	@Eꟶ�y`+�G�&�ႺiE�%��T<8:ο�p܊',�8ɦ-�o'M���I��";�t��Fl$�/t8�h�Fn������1:�FL��(a�H���tN���V�Sw�l��l��Q>윣Y�~���^�0��2�N�!iɇ`r�PJ^����4)��@����Aʕ�i�V�7���� }V�*�'P�L9E�5�iD��*�� 7�&\�2��n�X�^-�M$O���aY/����C��*b� )mJ�F��7�;�۬����XCv܆��E)+��.�� |H���|��N��BG �qR\t����HQ�bсaj�@f���_��R����Ѳq�x�cY�򭤢[�F�[g�����%>��:�uS(�N\"��+�dtH�E?U���hf�)�%��f�e�/Q�ϠL�4 �zIe�Z�6^\�p��2�(�N�H���'�\������Y���;a�L�7�3Pn�����c�����>"�SW��|&��-�1���g5H�#y��<���)��t۲�o��Nq]��z^�ȋh~Q��v�U�P5U�]���/VA�`��g�I��>�|+�������<�c�ՠ��ִ����r��u���r,��u�f�,��_����ɜ����@]���9�(>��y#��t��L�`�糬[4C��2��:�3ʹ�5�?��U���萋������ ;��Mھ�8�����҉���i�S��Ncrpe�2K��ݽ&�j���;-�Ë]���a�]Ғ[�{�����(�z���;�廢��Kaw�����>��c���>���\|�zM��L���?��q<?#�H�I���m�N��]=
�i�G����⁒�����0���$�K�K$��~Ә��=���Ք,�v=��0��/�Lc�5S�:RF�29N9��}KE��Ť�9�z�!�ɳ>{�4�ǽQ��1d�в2Wv�lԜ"㳛�p:׳D��v�/�)&X�������^��rb�Hȶ(l�_i����x���Z���ry�@Ҁ�'���qWrޥR�!!���};�����0cE���_K��BX��u�����OX�@�m��܂WgFiq�H{7�٧��yM%��ŷO0�5�-
Y9�R��z��6���� W��=���21J���7��Ew���/7m��;�1$w��f���Bꮖ��m����Z�w�O�RJ�矓�̹I��k׾WPS\|R�9��9s|�{�_2W��"�>A�p�i,�'!\��"��,���RHh�Qu�(!~�)mm�����/ L�y�g�,��H*\s����p� ł��
0A����w�� p�,��� w���ɺ�Y�Ab�%ɤ�ڞ�;��C��?��ҟ����wu�nۢg��{0����}�Dm��q�Cq����rFnA��10.b,�sD�!��	�a�I�����W筃N�������@�1hi���V5T?���.��P����ޮ���%W3�zᯓH�
� <��>&�T��=�Wti�,����&d�P���g�՗p_Ƕi@��;W��Iw+X�;�H.�=�5U^�9�``}�`/�c��F�).�����}�m����H�������W��t����\�i���df��a#�$�l����+ �v�F�%S�B�9��JQa���=-@���9�k�ӿC�� ��/���N�푟I�v�I�^�#(�W~�ԗ�z�tܿ�� �����q`�W����9S���я	W@V��>Ҭ�l=Q��~�S������p{�d����쐟���p�4#pj[F���8a]�ۆ���%�����зm?C`�kB�ܲ��Vh���⩐2�5��`��M��Y1�������}I-^0�`'��)H����p�y�ܣh�:xk��[Ȩ�]1+���	+R����PK+����/��Ԧ�u猸���K�P�UH?��O(�����(�`U��ĝ��5�[2۹L���*o�����	aa��p.�2Q��dye����]Ry�|��g��4�"�n�+���8��^��{u�~VOU�O>��bR�ci��jb�z
�B��7;�&9k8[�7&{b��*=��ڇI��.�&d��o����� ��U�������):7�g�5ϻ��=Ys/��l�1`���xj�,>���+�duoF)($]�|�?�L��sN��H����w��K�NdM
�е��3�fR�18��h�_���5�A�����VG�k���5n�U_�^�0�Q6d�z5��+u�������2�ح{�r�?M�����}VM����C�SJ��}��*�!P3{'_y��/�!o�^��7�Uj�%`���&0q���$�UX	�L��i�q�\},<�w���I����z}7����Dv�
�o�7�R���{�����M׼�^����Ǹ��f�.�k�;c1SG�(�ȍ��&� mt" G�y@�;�����`w���E;;�r�=`��H�W�ִ�	��ih��{X���q~��q����Â��i{%4Urg߬�ȿ�0ե���5=�X���|Ɋ�j�p}&�q)�I����wW_�G�8�9~�ܬK�Ҫ�V��O����с乍M�/"������9Q&	b�%�w�� ?��8d�M�� ��;頁.Mg�G��*i��^V�����:����e@�Ѱ�H�i�M��%R�hf�&s�<W�-���۔� ��&Msz��(��ޝZ��5�{_��K.O��y���p ���w}mc��@N�9�C�=3f���vY�����AID����[:5B#��&��`M��f 0]����)��;0���R���d:��8!�Z`���&ݞ?b���'�[n\H���(����(�^����	�].c�����K��3-����n0�MڴZ���Ƅ������} I�! �YIſ�*�.��c�;��'
wQDp��W� ٹ�񠗗_p��>�~��'Xh�Z�u�R;2�G5VE������T�a/i��t`���y��WP��#���X@�C������S/�	���� ��ݏcTZ�۞���w1.�s�&"&[:Q� ���X��U=��g_���s���rO���Z� >�YK�v[,��& OS�|������Ǫ��[]E[����~������s�J��(ЬV[��|�}���1b�o<��%���I ��iج���Q��]���b<�S"��~B�zXH�n�L苓8Sv��|�@,3Z��ZS���O�[����{��P�0S�:�-q�b(�d��U"��ͦ��[D��ՅY��L�.\P]o���Wɸ}���-��j*b��@�Y�G�ܟ4�6��0��00o
���-���ETX�b�9��
f���\U��D~l6�x{H�g��y����D���)�&��E"C�U�l�0��6��yW��=$Q���-N�K�<$�mD�&;n���>�)���fŨ펚��ڿ�L�!K�.f��{o���ˏ��6"w�2��2�X@��פ]N�i|u��<b��������@8��W�R��0���]��%�#�ڄ���H!�|�As���>����R��_&��t ��Tְ�1a�L�5Î! v8Mj�Oȳ%�ۯ枡\3�Y��D� �'��H�	MĭU�q���|���$�b�;hyw~����8^}�u6<�X�vZ�9j=�׌vy�?F�6b���!|ee�v�J��m��p K]3t�j��^�D�����ŗ<���r�1"?�VF ��k��ͥ���k�K��OW]=XK�1l�	��_�uϔ�!����u?'b�FYG�(
k(����|�ϱ+bh�C<��k)Q�q3��*�n|�;ǅ/x�I���0��I?��AJ��/�"�X�d�RMˬ��m���@'/��=�E`�|O'@`z{T<�R�.|�"D�!����C��n��m8w.�T����	��(*�ʷ���j�7B������������{W*%��[�vao�x�-iq*�3& k�/��(j$�G=���V�i''�E���\ҥ|q���p..&Em�"��i"e(y2���1�oP�~��� X��V��|�����˴lE]O��N��(?~���p�d�P��M�&�{�����}4�.4+�R�@��f+,H4��B�3���<�O�qS��ˆNw�R�u����!�f:�چH�̡����Eti�	��W,X�0y;-s"J=��8K��B����%��kK�^���K�L���Р�Y�5�A��\V�e����Y��t�w���zUI�*7�-��)ΰ���1��Dv�'8]�3t���1�W���M��	���˦���"a��TL�o�$���
a���(���Y�_6W�H8��j4���AĄ|��Bq�\���������	 �C��Sm�yl�&�̇h� �G鶁��ib5������l�̚C�7`N�A�D�>K�df;�`�8	�s���1C�rK����������200����Z��C��V���*S[�m2<���h�/�J�@�������H;�Ŝs�r�}�*�E���`QR(~v(9��^�\�X�W�aG8
���B�kowN6�����T����P�*��|
Y�p-��[��}���m�j�U�Y �l*p���\T\S�'��F�=��!��B�^���C�#�Q�=�W��R��ܿ?c�o6E��u��9�ΧM���B��1�7��K���.A��Hێ�t���o��6�O�	IoS�02��{����b�ld����|Y��D������f����Fɝ,�p���W��;ڱ�*�/����e+*~�n��NV��N����"ٳ�K=�͟Xi��#W5u��lc�r�}��H�&���+���Vv�oA��!ä���y��j��c/g�L��
�����
+"��>G0MS�[v'&1)ú_����l�ݣ�1���Y(�	I��ک��U��؟}�/�^���
u�B�(��rv�{W���f�x�༱�n�w�@���ʞJ��h��q����1�
�]z iĎ�x��>���rR"����m�[Y���oa㯕x0�R�Q���OY�mLg�t���}O4X?��(#���a>D���-���6��i�0>�+hq���W�kE�2�̂�W�e�-2C/T!�yۗ[��F�T��	ir[X�)sX+^���FL�ȱ�Ou���Gu~�5�DNc��0��J?�����]�Ƚ� ����(.�ܟ��Th#�rXOp�>�y�j��۝vt�h'>I��U�:<����9bR���j�n�'�K]N��]J�3K�	Tȋ��r�,�?O;KSDz�b_8%*�CuV��������!���*��ګ���W>R��g���F���
���ȷ¬V4�"����R��x)"� �+I�]�f�ԭ�g�;M#F����7om�
��;s�-?�w���Ksr��@4'�,̕2�S�#���h�^�s{�<@����,sz�������r�$�@����I�7����-EDFZ�*�W���%V �h'G�'Ҁh��ct릌���V%��@.u`EY/`�\��ۋID1��)�5��:sQ�Y#�(V�|��{	k��r���W�r���k�KT+���ϊ|��䩽�t
�ps+�3��Ma���w$�$;���-S��C���({;��1���G�`����-v�=�s���r��m�q�s0n��ьt*r�Kӻ�^�T���C]���O��`�c�Y��YO����	�`�E����(�Ud�����^Q��埄�{5e���ʱEVAy� ���i2a��NeO����ujM��e�<�G�sX�gx4�6
t��ͯ�${u�bA\)�톣p"4E5�:�E��;eW,I �/e��K(��\o2�դ��� ���_i�V��R3��q�洊QӑC�?LC��]z�z0ӡ��\x�>�ҽ8`�`չ�}}ԋ��� V,��\��򮂹��t#~|T���6��:��"I��l ��E�n�u
}1WxT^DV�����Z�R��VA�`�Ձ<�a�G�Ab��'Bu99,�c~�rc&Je>�3�]y]�ƥ�F��`b�n����k���bn�5�"x*g%�g0 �Hd?C	�Rn�I�Ʈ��s�y�$Sȵ%��T�Z������N�����!���T��Q��:���}�!v��:5��-��4QWL��)���"���N�R����y8t@���,�{��{��<!*$���d�&�+�5[[�� �qtT��E�1��//'l��,����n�(<@�@��G��S�[�;��%����@�{Cl;�?*WFH���hr�0Y��%�;#��227:���J�>�;�Va�7րʐ�7�h��N��0�m{�KPJdf�o�.�6�g� @�#������)��b_���(Ba�䷏<kֲ2|Z�����Q�0���)���2)�Fs>���r�����of���"����cQ[��*�	k���A�4n,?l�?.���^=�q�����Y��2mv��������y���>�IZ�OaP�����>>Wl�0*��b��7#�," ��1�x,�0��i���K!�f-��<�G4\����d�l9x�iFn�QI��՟N�pw��M��|�0�I����>Z�"Rm�m*eZ3�Ĝo�JV�����YX���I���d�,����*�C��Α�&9��3��[�YW��a����L���LEd������Pt{E���>�qd�[Z޿���Ԯh�]?�>�������W����M�����C]�6,
��F-�>�t�c/�:�bE`��3��ꔁ�Ry3�Wm�!>�a6|����к:��x�>b8ˏ���}��?��k���?E~��;D���el�^"dP@i�!/i��9lW4#A��!HRxS%����|WJ�Q�G�$3� :јn����tU��{�\�k���2��.L���g�z�q�~�nTn'C���/B>\
yD7��4e<�7Vpǯ�p��0>�[jN��VA0��ٕ�}?�:*��x�gA���޳�Zl���6r���l�rZ(��~r�D��	̘�����	XE�AD�.>0���K��`�R'��F?k6�H�U�������2w?�5%t�o��-�����0�`��W�����k`��z]��~=��D�����倇�I|�L3�A�X��1�����e]�ա��HdU�'1NO�Ԉ���;��e��|Tk��������}o�&���!��քJ�Pe�cH+r�
~C}U��{��E��Enm3��Z������m�`�2Ѯ)&֋wmn��,�r�Ň�F�Q�C���!����|~�%��ĭ@���Y�CH.�e$l6����bM�����`�#& x*=��)(�̢d�	{& �-���N��������ȸ��T��cR��{� a�J�R�q�z(ȹw/�ȳ2���	��4���r�����~\^�c���Tԁ��Pw��4�|����G<+��9��L�%���A�k��<�R�F��7���]�:�,m��џ=��G���k����������u�?t��<����c�'8����֭)�I��(I����i�Ƽ��|W�1��7�{�)��ZJ��Da���.[j(YR1Ds|S�6/�8@蒧}���1��]og�(���g���h[:���:χ����{H�)rl.f��h���C�6�B[�
���7���j�k%���Z��ӶE�S��Z�dٻj��������S��Cͽoό�VX����t*��\���1����e���4�'q�|���\�i[�V���C5�#���&��?����(}����]5�<9�גi�A���<Z~E-U�Ѵe;$~��,��#Ȃ
�-�?$�n禹�:)��$@�3��j�^�NV��i^)�E�q0�Fq̅�s��G�4%"s!.��RS��ђ@-��B�I\��$hk֓p�Q|B�[;�%3��a�.Ѱ�p�;ޤ�(�|Jb/@�iH�*��Mcƫ��@�3K�W���fgj���&�'�Z4d�۝M��LT�b��^v��M"�y���Y;�u�9��.�}�H����>�ůE��V'�5�l��m'�����6�q�e ��D��b�W,w aԁ�ת"�-S�%;��[�j���b߆�8���k���Q;|��M&���F��U�'jmw�tqU�z�o�%�0��NB�$�����zι��AеM��������H՗����lāV�jc�]`���!�\�L��r����FO�OA��l�N��a{>8�Z�V9<����e/}� X����p݇f.m9J�pS8�0�̋ld��뷁�8S`hx����R4���"(�#ƞ���� PX��>��$�z*o>���6��9Є"��7��5%$�AbQ��jpԔ�a}Y������{F��إ�
��,�{�/�"�Ғ����ղՉ�ȳ���!fm�sz�n�.ߓTɮ�ㅽp0��ೌ@�'�/���<�faM�R&O�+!�)�3��IB6�U>�:_�v�������vH߶n��Fw?å,7��&�L �YN�3�T���W>	Bk�Tf|X��O�F͛���U=+��TKy����Z��-)�=JL/5�7H=S��J�;ƪ�>�j�qw-K[|3��P���@�٤�/�J�9^��|��/�JDj�NoϹ^���ڄ��%��� �c�z+�eC��D	������0%ш�����yE�O1O�%'
H(���ӄk�k�6|Y	;�aX�IK}({%"[kXAJ31�S�#9���[bՇW��+p<����'����q�y�D�c*��jOַ�'� >��A���@O�f �A��@hZ����]�㕫6�Z���6'�+W���Y����)a��3N)��k/B���y�ߦ�0��9��
G��T>�Li�^^���EJ�Kfe|�.���@g#{��]�W����$p:T�c����Z����ex�ȯX(>�5�T �e��m���y	�j)9Es6��[m��1�ְx������û���#m�|@n΋�P�[:��I�=�6dυ7���� ��/
��9-z��BAb� ��,�ԗɟHrZt�
�e=��#�+��5�㡏Ap�X:d@C9��N��"E�Hӛ����Pc� �w����r>���~��I$� W��M�3\�([�}C��
���U������7�on��S�8�9%���]{�o��\HQ%�{q��u;�K3����=����T��5+�V��Ԗt6��j�.!�(���*���^�p5L16��<�M���y�8K�z�?� W�.A
d5��� �-b���{��y��4��j}t<��a����B=�o����=-�dn�g��%�;�"6�"������ճ��E\K�`�ۙ"~�r#A�l������.��ֻ��˴����y2���(������o�F��g���~�+6�f^Be/W�c�7���@�c�<a����Lg*I5^V�C�2ؖ����5^��1y�n�d�c6�-j��YNЗy��Q���Y����������̟VQ�z�� ���W�$O�@b�Z��gW����i�%.
Oz��@�D,�x�H�\�6�	���M�B�����>KCG,��U�R'+��N�v�����m�,U��Ć����8{�J�_-|�-��Մ=7]6���
j��M�C-�)Q߸�Q�#�1��������|�V�& <��o6�J(����֜ku��C���
�B�X`�7�xŢh`�+��a2 ����:g}pU[�[�tv��6���;ʀ��Se�����	M�d���_o������H��BrB>��3L�t�ȍN�>ø���s���~�F��]�A����^\`]X�V���ie��K * I�N���%*}���AD�DtO-6L盾M��y-&�4�Y���#��:s��t�7�(�S��`�������9)^��}��À1.Ę�e���wx�Z|��.^�]@�b}�H��č=�,n+<ñ6���`5�4Ou�XK�m��"����\�pg�f�N5�咛v��ڜrkA>�e-���e��D>pD����(�I)F��+L�Ql����^}DYiB�zM�4<��#�?g�=�Żi��o����b�ҷ�����6V8�����N{���.�����\������+�%�\�����x�`��OH5��k`#n��ɖ�b���DB�ʶS��dɲo_{=*1�����~�U!{���,����Ȓ��}����!X��	Z^U��d]h$1����pu���A�o��\�M��әB��7&jy)�(�F�2����|0��rt��|v� 8|)�6��T>�E~$ .��k����o��Z4�+>R�A�My�o���X���臿���~�ƛ��d]'�]�b9w���hM��#��J���'f�ރۜkI�-�68ag���'�9�q�o4�p���/�ь>"�N(�Aϻ�0�it�W�Я�����)�0�/�]��$�^xw�"ɰ=&ve�U���7��o���,xǸ/��~~��vSp�����:�}���ǉZ�ב�����%lȼ���#/������oV�P@-Sw.S/S+�O���_�{*�_a�������#<'$�R7�K�z�Z����,V'Y!����o`N�<�SY���3JoR>��F��$��q�Ia��6_JB���:��o�2�AQ�7��9��c���߉8��ۈ�Ak�$T��T��l'p�}�p��;��� �ۤ���X���?��W&��7d��MK��<��H����AC���Z�z��q��c�k������B�
*F&��e���w�U��x��(%�G�3Ck����7}���ǵ�ا�_���K��\�5��<%�ѹc��c=3��.����h}o�{'9����,�k':;M�\�!�j���BG}��=����U	+$Wnxb��Bg-֓nn��u���]�����J���������Z���[��KK�����M��U�wq�h�W�͐ χ`W^��f����ф���OԿGDK�k&�h^oշ\a�6���D*��*�f���	��ͱR8;R����=�)��e�N��*Λg,[���@6�U.�+Ay?�G�
�Ţ�����|�(5�P��m��x�Ӑ_G�
a󽛕��-��?�W�sy;�� �0$O/�!��q�-+�H	|�IL�����^������e��_�*q=x�˧Q��v�n�1�c]:�}�@H��6'���0Ln�	� cd^�Ec��<�x_���噥+�XB"��g��ӺC� �O�_M��IV1Ӄ�ū�*��S1������5^r*@<u�=��]��4i��n�o9c؍�	�MF�k��Jei.�c��wʸ����Ѥ��2ÉU-BQ��⭑h�BC�S@��P�*.||��0TE�Ʌ)��b(��S����d((����dO��N�����+oS�/Zfuoܫ���s]3=��k���������[�\o}��pǞ)gl��J1(���H����d��Wm�3��K��r��X�I�>��	Nw-����Pt��6�#4-����hei+����4z�0c�_��qK ���7:��:���	��1)>�Ư��2,P�U�6���-*K�@\�?���`x�556��������cD���}܃��i�tN�L�R�P�"rU*��?����ų5�=m���5�E�[N��������f�����_�r{ܐj~�\�Rm� ���>��a�����U�)�~��I��S������c�	%��}�-eb,GץQ�<)*�k�$^��h�C�m�\�i
^���2��xz�{}C4����/�
�wʼ�͞!�]a���_Wi�-�x�wG�%Z77�+W��ĔxCʱ�'O�d�IW�N�� F�&lv/F��7�)���$}�u�gya}j�N��_�E�D ����n�q�?쨉��&=[*}�`��z ����!.`�6y]T�z�q"Q[����CI���2�`p�9$A�WÍGAK�΍X����G�
����H}	c��j��%��*���W�:%�vg�n��ز�����~b��W��#l�n�q�>����ݍ9�ƾDgI�_{"d�m0�xO�'��~���:�HV�FֶV�ٌ�<ѷy^�����L��+���*W'�)Ì%L�?1q��7���׽U���Ԑ�7�,��M��J������x��o�ʾ{si����7oxewe�:�n�#�V�E[���BĊ8DU�5M�&]Y�x"�3�%�t<��͐���
��^NK�3��6�������'����~�E�����R؂��H����JTz���!��{r��`,�~�
�W�q�/�����6o6��n��tMP<�������F�Z��F|=0��~r�F`�Y�ŀ�(��S�a�g�T�;��]��]V����e�6���`w���c���ܭ����+2\c��=3�u ;�k.�;�̥�\���<z&�b���O\+ӏƹ/q������C>�c�Ŕ�N"�����=m|^C��)�|���;H*.����F Q��lK� ���.Pn/%b�R�~%���L_tA
-�����nC��lz˟k{�hĒ�:4�
��<S��Nĕ��7��B����HD�Sp�� hCS��([��n�}�=GIGrDl�$�����;|��Ҭ��г�n�9���3Up��?SZ㽚�TŪA'�Y�6v�u�q���x�������飆�����^E{�C���C�RA���@��`���ӎA��2+���
�[&_�F�넞�A�����DR{)XV~x��h{�'7�����M����73���ZG�;�N�I��I�ֱ�D��!�[eA�tOY�ٚ�iu#�,�~���?��uFr�B������񱒔��ucI��嬎s�������,�E�х0m�2 �8�rȖ�6"�k��g=K	�2.��Ve���1�n?�O�Ư��!�^#�A˂zH������-�P��;k��a��w:?��≯�\-ß*G֬�<��DK�]C1!�\��qNR�/����)�P�U�ߘ��,��8�M_���gqI�O���pE��6E	�E�+�eFn��/r=JĴ=c& j��H�ő�lW��̡�^��E��5w�4���X���>�
(N�w�)���n:��ѭ�uG��b��������az7����n�خ�/��o`Ė��Z�f���!xv����cs�� 1�I��UTN�0�(�cV��+h�4���
���̶n)"��c�L��d��h��2.���J��fT���F�(����\�U\"���yP�3v����C�ٜ:ݶ`/UH~
�P�iIK�q ZA��я���+�V~�7ܞ��M���V�������4��F��~k@^:�Ϣd��'O�&;b<�
�+r�MQ,��eڡ�r܁�j^�XN����;aۀ��+���q��b��b���|�@P��`(�"�0ڝ��������[�ӈ'|f����� �־��Š���p%��ƌ���GJ�R�b���y������ UO��XC��tN�LO�@�q�"0�3��-x.��`��CQm��W�禹�~�f��ߺ.q�)}e0a��Q�$r�Q[�m˃G�k������|��vg�Uߏ�ca���]�kW�4e_�4���/M0_;k<���d;{��i�4�����N)��1U���v7=0֘Vq䉋�j�:���.u3ϖ7�t�/�jlG!;��PPL���{w���=��?5�֩�c��fwaB�vdҼ�A��G HH����e	��� �M�u$�y�;z�f�OB�KM{Hƨ�	��m�����_EI>TK'�r婋�N1U��d��`Y!Ğ,����B�m7��;:��H@�Vn%X�����+�OM��I=�:�A�X�>��<׍��+o�Ӏ�)��X-��W��*�d�Yr)�B�#~eK���Y�nsE��_���k��K�Kk�ޓB=R}Yg�G[:�Q}���/�I�~!���!eI0=>(��k�:F�rT�l�ϗK��n�v�,{֋ ��1K�-�˺Ed�|~�.%�:5.	�Et�����21
�af��^�����y��3�\>z���x*p��z�h;��Nz�L2o�w��H�Z��ǭ(����?V�RW�4 ��ݞ	�I�d������x,�t��X)��i,P+|$�m��l�b$*n��Xx_3/�j��S�LPN��~�@��������d�_8gX�A5� ��"H_�zِ�3``���7�k���N2�����p����x����jer\W��H֕��|n@�t���C�� �R�XY�H�2c�������S�&{q�k-�J�!�/�˖[E9)ԫS[����[oP��r[)x�u���R�7�������IQ`cQ��,���?�R���A�L�s�X�w_V�πm'MC��r�g�ν[8��#&S��`vպ-�0'�=���m����2_��с4P](�j�+�)�dYͺ<I�g��B2֢�o^��$�l���t|�8��9"@� ��.�]˺�F&�4��<'�?o9�)[]$��9Xۆ�ԡ��"Z~�#Eb. �����A*c��շ��T�h�M,A��G.�/"Ou-$���1�!��rk�a��-P�M(%����1�w��[ �z��LN��k�-�B��}1�:�m'"h=��i�M_K�خ�Z�a-���4].���dw�U<�n~�J������d�DOZ�s"��ODY��Eb0S��ǈ��b)
H}�s�/��7��mzB�5��jUE�� E���bk��v��O�3��Hݱ�	��4a���iY�B;9+�Ծ˪60�H�Q���A��'O���R\4ǌ�����U��*���3Q|�M�գ�s"Gٺ�"x+/
��ki�Z����c"e��/���a��{�Ň�'p0�?�'������:_���	������₊�a�������Ӯ�&~��*�32=��=u�̵�����i��/L֙����/<��e��F��p/0�I,�G�i*nW��',.W��f.�}��6��?p��r���ڝ��YI&��qta[H6���kt<w��_%�F�<~ �P�A���yB2�`B��Yz��wF����?�F����gę�zSR����B�|@�o:�6��W2O�1bd�;�M휃�k�A��|?R�M�}� ����Eo]Ry��}#5�x�����5�]��j�L�0�E��fSs��%w�d��B5]b�f�e�~��!i9�������J�j�Q�w��r��:��Sc�i�035hVN¼�	�}i��L�t��b>HNϽ����p��K�ĺ������iFV��쪑�-8� �MC��'؝��4����1��~E[$3��Փ7��˽S�H�[]*�/�oK\	��&�j��X)�b/���^'ٖ
�����lO�ƃԠT����]~�)��|�����Ds�+�	��@�лک��c�栵e�����#�:siW��H��y��/���[��u-Z>E!�ѐ��lh,!�U6~z�{��/hN��n;�����blK�E�̈́����7���P� ���@$4x���.������^�p�Dx��w��4�7�ѱ=�؛5.����2��� �Nᝡcv�G�`������{m0��;NW��w9Na������X���J�LPX�Dx/(_�fj��]��� �I�+s&�<�I��1�Rz2C}X_�ex�O��y��+�ڮ��L�r�l<�5)i&���	�����ɷ1}I��N��dA�V���,�a]��%�����Ct1��%
jn+/3]l�"w'_4p|d[ѣ�1\��M5��yHҐu,	�P�}'ܙ�u���L�Y��2�#��С#���G�@%�!�s�S�~���8S"E�{$
�=R\��Š��i̥M��6^xӮ�f�8��L����Q�U����W�$1���(��Tt���h�ѕ�����l�$[���ea�������p4���n�+�㎃���+MK-v���p[��j�/�~�E�!�:k�'	n5
��`<φ��Wk#�a��Ir_��f/H3aG�ؠ
��g;��a˼'v���{�w@X�ѓ{��譩pY�8Qe LŁ�8����(ߓ#:8������MJ X�bO�k���^�J+�H����)D����U�"�a�N��Ԩ�DMLD^Y�_�� �Ź���~򶦲9̏�1��������+��6��V�N'>�ݢ�/quk����D.�f٫��b������$�QNq�����#�
�3I{����Q	uٖ2Փ3���d���%��S#b;��������;p�X��w�y�P�I[і��}�&"ը����7�>e������Z�@������B<tT.c>�X�_;ʛ�-L{z��TG6�� -bu��ѨA��b���y���	�k&��6_}߂+\������a��۽ޗ߅o�Ȓ���%��NzB����i��g�	V6k��.�s��mS3fJ�G2�[�ؤ��<1`��86~�kM����.��*���1;��d0��T����"
�B��f�R��	�n�g��@"6L��U�a�I�����+��Om�V^ڮ�I�Z]�K% ��)�X����R��Z�u���:8��;��w��
�w�Ua=�3E�:���73�IU�S�;%��Dd�q�ŠXp&�g�%U�@] La����?�3�{�?C����c.Ʌ��3� ���B.�}�i��s������gFm,�>uL��V�lL�ѡw�'R�����d�� ������#?����L��zK�� m[��L�~�.%�c��-���3+[�\ⷵ��מ��:֣��,~��?!V(�^YЈ���� �%��K�>�v23��
���� nrF{�:�,*�]'���PH�����c�r1ﲩ,���-�j������7����h�����K��υt��Z^�e��&�^B�r{�a�a����28ȐG���jH�h �+FjC��U���}|��WQ	��f��r��NH�3����J�Gh�]f�}obس�-���R���x��ms����0r7N��"��p'�[5ƲG�간�Ag���@��:,��z�J�M�Z���;�� /��$�����!C*�iDK=�f�tl4�
Ӥ=�vCb�%��������yu��V�J�.��2v:�8�]��?��Y��/�bmg���ޣ�"y��y�s����퍿:���#˭�@;��߯h������������K�-\��dŵ#��7�&���S*��r%�K��R�ȵ�*�L-�KƵ��ر�����ѵyΩ{��~J�!��*�o���ä��!��d� g�b��>˂9�d�.�mȬ7��=Y���	A�E�l2��u$���Ёm���}2���������D�հ�t (T785+j��1�Ƈ�r��N�ީ�Y���x<Ɛع�0��,_�*owto%Q���$ ���Jt�s��F��;�@{5���|�4<Mh3���ҥ	f'��4iB3����G ͻL��`�C
{�U�����3�D�e���2t
�g��H"�[�51�6N-2IP��;��W�ÞP�;x�R��۝��/�Up��p�����Ӌ�OU�0��#Eo8��������+:�Q+�Ǉ�S�{7�c�-�|@ݽ��"��> p*�d~�(���}J�ݜ)E�����NI��+� `Qm��k������ѴMCb���g��.�ml�2�LA��=��˳1U^ŗR�KE#�\�Ճ��(c՛
��)?\Z��㿮��U��DHߥ}A�L��4)G/��7��6�D� �y�Ϩ���^kQ _���/�����;�t�K���E��.'�Z�"�n'Qb���F���~��^8�����:��7���R3��A�V�ڑ`��˰��R� ?1\/v�J�E?��;��w�w��+I�	�P�,x"�F�c�yT�O�p����-�ѵ�ϧ�֫��Ӵ�+������X$v� ��eM*��¯`��,yG獉<����q_8�9=tк�L�cHDA�� �f8Y7�Z�f1�܍Y�J�kCu�� ַ�]y��9s�
����vH��� ��I]HӔk*�0Ή�a��l��X���F&Ԍ1�|B:J�>*�g�/1b��}+N�Y�T4̩S����cLk�GRC��\,��x���Zk;G��iM�$/#.nqs8n�ǂ!�k%�,���B�������/N�K��퉄��ā���mfG��{�#_i�Ι�5��R��]h@��'f@n2��x	ܔ1J'�k�����"�	��L���g:��3@�یB����{�R�+��2�z���u��F������W�5�D���I�y�r�-�d���dЪ���Z��ӑYR:!�E��,@wX��ǹ��gQ:�\d���~c����O����C����*�])�	��n�-��}-�&H��K^�_��!>.�4wa�"�3ἂ^���t�\���HEc�Ҹq�
�ZW��;�N$߹�(�~�1���G�Ofb���$�p����~�GeA�_�硋����`�A�����v���ME�C�#�(W(��A�(��aw���W�h�wq��q+�Hy���ݶIE�St�:��s��|/�]��cr��=�>n(Ƭ��� wQ���G���Ek���u�82��)	$$���j[s��!rn��{�?f62� ����V7��ռ�3�����1-bg�k�L O2���S����m���[M�N`Pm��:��S�>�Y�N�_V�؞�	��q3�&T���e]�`&w��%I7|�)a��cjC����M��X�'���yx�C�;ܒ4�����0��7Ed�9�ߵ��M��Nx��OJ�;�>�vy h��H�_oڊ; C�X�P�*B�6R��/VO݅d�ܴa�Q�B�����\&�5����C�.]%�W��@�,�sPJ�l)i�OL'���_�ݧF|c�{��8���W��.�����FbLY���9`eCl��N�M��3ڢ���̄�������.�����m������*(J8�u\p��㨤��~��>��/b���iCv�q��9�)ɒ֯b�㤪3XլB�R�������_\�7tٵ>:�W[M���&Y�9VFPV��`�bp�.?�X�wuR+w������8%y�h�KJ�=��SA�����q/|W������Y{sQj�%lU�e)��8��y.?���zumcq�f�dm6����[Aȸ{�6�{ߛ��^D���ց�y���b	X�?~H?Ci9���@}wZL@�O(����.�����K:�|�_䡒j��U�$��6D���7	ϧ	���K~�!jARc��ͥ�#�y`��U�dmgݓ߻rP)� �#��ܨ�KIx鿕PnDk�Ӌ�'��ǿeήP
�1k�.�����?���n��V;$%��_�	?c�r�����V�q��� R�u�NW�h��hdD�j���d��C�/@�!�|vK����j��p���;�N�|_��:@ǖ�܉��\D}Z�Gw=��͈��j�Ppr_�w1�mv�Rq�_�k�Yu7�#��Z(���BJC�\�<?�W滈�'S:�'ǵT�~!�m�n��^��`�,�a�V ���1�tU��n�aPK�X�z�e_jEO�ǱnT2�x���Ĩ�D��v$��1�g�� �9�W"h>F��]��W�>�.���x���(;���R�;\s�J��d�{U��u�zn�iz]����5_�M�m�⡟�L2g�u�\�k��e�3�p����](��i�߂��Ӆ70LՒ�wA^����P<�&�K��DBj�R8�b����5���T�S��䖛VT�?���*
F�we�C����Z[))ˆg��5�*Y���4��Q|�����Z�{w%���Z(�����'
b�U�\�]!e��*I�\��y����[U*��A"%���z] �� lwq=N���'o���F�hQ��R�Ah ����u���<5����`b�HT����j��u�@�*��U�r���*9|��#.z�	����s�>�rp�I����b!pH��%4[A�GF$�� ���1�~j~fy������v�H���K$.'5%G�49F�>"�)eFJ�X΂}O���֒k/"A������y/S�j5f�6�CƬ���w9��t��!��&	T$&gD�� ��1��m C����~����OAl��/��4��ѽ�g`Y|F@���9�J���	%��^��*��K=��Z"_
�_A�&d2沃N)E�N<��'sA]4��,���,�7������l��>Mi���� Ɩ���*�g� �:�y٘6s��I��g2�b�c�x:D���yax�z�'VX&#���`l)O�aw^g)�s/�^ܾh6f�[@�Z�:wOI��iI՘���@�©\Rh�		��ݟ��fpL���V,G����`0 �BL�4�IoSM�C,�"-��Ώ���Nx7Z�<�����AF�?��#)�]�S�i��b�kPQ����߽�˄P���+q'�'?�`�ƱǶ��0����dxS�-�f����ҡ����az�y���W��9���o⥯éN;���Ev((*���Ɵ^�G{c;?�`�q�s1��]r̳n"�h�ɩyoQ��O�S88EM�h��i!~�N�,��D�i?9o=p��TI��^�4��n�^]��:���02|��Ԣ'�$�s^,�ilO#�o{�\�]�bs �kL��T�s��{u�\����3�Gu��}�g�*d������,j��Ą������|t�3DU�"��K�~�թ;T"@�֟'��\��W��9a.�{ ȳR�� �ȍ��q��lH�v8vLoh�wQ;�)�w���ô4�9����XEB�j�vJ�RtC��],&��Lx,�	)��3����8�vsJ��B���fi�@@���d���DM��k�iP���������zɩ�'�6;���h�C/���a��Q�Il��V���Hxv�$b�����o��:��ml�	H��k���<�+Ci�z+9F+υ�NF���$��+�f{�&���ܰ����ܣ���x�,q�;�m�͊Ɗ�_���I^V����>Ә�E��z:�Z[�g5E�M����`��:A�rﴬ5�J"��?y��L���x��o7����D'+I�JS��(Qy/�5=�B������"(H8�(�C�2'B.�'^��n��+�	���EL�,(�q͵sZ����T��.�Ւ�W��Q��<�J^<54��:M.ɟ�GN�˻h�)}����f㶘�V�z-���s�Jy`�i=�ƥ* �f{%d�e�=����,
G*�ݻ�p�������_���@}_]�����,0:�0�aЌ3T��S�*CVj'�uoV��b
�v���\T��۸!' ��&��W.��$d����+F�� 
���I�˗�I���r�������ʇi�~�]�T���_��$!ʽ�}$��"���<`n�\{�"s��0=��|�4P`�үFl�]|�%?�c�d_��>���E�����:���#}?��1Շw�MU��8-0u��ZC�+���#Sap�!��[�iÅ��Sg���B,��(
�G[i�t�]�G��djJ��`�P�֌�,0#�_fq�.�����
(�v���*�\�O�����+e����ӆ1��q���Tor7�����h��,�&�F�ǧ5%v�
~�S������}���IQ��DC^�c���2&�V�l���C��Z�X]O`�����nˁ���/�1y�f��A�o$��G�X�z�c�=��я9�_S�%27�2��&r�
k�<G�z����\�[�^8:c�?�{��>��!���W��r���N[���ͦ?���wD2���x��gK�1	e��H٩F�#g9���X.@���0s�g^��=h�v$�M+�0�Wb����?��
�P8�c�VI??������^�q��M[]�����h�N"r%��Էqj�F�]�d��1!�����,֟R�Ң@xQ8�4��eT[2�ݱPg&aO?-ZY�|1����{�����8��?:MV�����ac��iI:{a��b�ڿYշ�Ť�EI��B&67S��PPF�+��ԭ[�ƟrM���c�+@$��[����Q�*м���?�-�%������3"�|Ҿau��U��5N-O�`�EE���Y�N���܌ѽFR����GY�#Jvcl���h2�h��Og��o�o�
�E�d��E��A4=`��5��6ؿqgN�NR*�oAP���_��<�bP��h�	pKD4� ��-L�*�{�l�\/FO��� �I/ڜb��koi�����sG��
Qp)?�޴P����.}���|�&u'd�>������
��Y���K��e$�̟\��\�����#j��U����e�h;�IH�e��� ܣ_8yBfH/�I��E���+��eV��f���~J����U����p�	!�³��e"��O�N����ʟ��Ə��yP�"�6�םU��
�_஗��۔�-���*g����P�8pn�� b�rt�<�L�3ϼ�,����-8�&r=���/�s+����Eਯ 2:��C�C�:�,P(�I�Pܸ����	yB=��[�,���Pf}�@�	�R��������<�@��-�Z�Q��* �����8���^ �`��`�o���X�+�=
�}�z�p���k�R��#���m��6�|b^`T��JM'�4�eU���ު��:GXCKJZ��?�O�s�;, �y-O7(u�X��Os����/�T)�׵�2v o���}PCQQ����'e�}�:�4��o�y�	l�#8�
�
�rR�S�$�k�|�(��|��Y�k�,G�'v1�ƿ�sF�W�S[P۪Y�����/`u~�/|~�S������f�@ivhe97w�>��ǯ�Y����7����h�/Y唹��~�'�1��Qf����<��d�M銚�9�*��J��_�}$�(�Y� ������A<��Z��g��e�л��&�	����i���"Hߩ�G�+`��|Cg�!� ��IO�U���31-$?V$���6*6�%�L�E�_$Џ���`g�o�4kE�*�!x�dF~�E��֧��Z�*�������D6<��=l�በ�1M&�F����3K۰���p��y��~�(�:�uHKPv�b�H�A���Wߕ��\p�ߚ�i���Z���|�����R�P�C��[Mh�@1~<�����*�U �Nl?w�Y�Ӱ�Rb��*��9W��&�*�X�b6bC`���b6`6�a�vځ���?�߶BY̊
��K$|�4����Q�.�?�? rFy"�Q#_�-@��g���
��]��\Cx9#�lM�x_X���wV�jL$�y�=���0��\j�v����kr�O����8Ȃ7!�oB�fG���'*ٍ��ېVK(骐3m��6���1Fr%�x�l_�hŰ��J���l��.��Dn|7����X�>����s5���2���f��!Bv6EE�O���A̡��ْ]§ַ[=�m���&���K~��2�>[��}S��O� q��E4䥔Z`I�.b3�S�����q���z��n���>R�*��~�ִq��A�Hb��z&�j>�#��O���s�;"�≔yXX�����9��M�7�<���4�p=��Kt<qP��։�Ӑ�h�>L��p�_�%����t_=�Pޤ��$��
�ndH�4���� �s�8�5,ꪌ'�{`=�2�3���8�^�fFNkV�'w0$�a��	��_�\0���/�P�{����W2�$9+���iX��ҫ�����Z\;�Ւ��#yY��Ž���2{��ӡY�V �|;*0���h�`�����Ir��}N�<�b ya��땭��mJ���鎌uce�x�P(���9p�ߍ�󾋜���*��ئS5��?��I9/�#�w1;x�
����,$�:*^#�U��6589^�~Q�z��f{�1�5�)g������	��4)XŌ�Mm�<x]�³�Z��Jl��@��q�_P��b�DkSTA@NQd���'���o��m�7����@�ĝ��8&4M�6J4�)��z%Yw���ǭ����\ �e.�����iF�xJ���2�S9�lS������_��phB+�f}��[�N��.t�O�8��p3Ѡ�+rB�z.�k�T�
baV��c�����Qf)�e��/vX���9c�˳���u��΀P&�p���-�!6��ʴ��'��h�9&.��"�����X �N䧊gp�����.����3��{!k�����BN���꿁[5��x�+Y�R�� W[#�9���k�Ӏ?)�<�GVh��C�l̉ZC��r@��P��/R޶)�v;����c���g�Ĺ֒5��%�ĉ���uI�L�K~������,= �k�HM��wyǹ#h�F�-ǧ�M�}Ƽ�kӄ���zڴ݅B��BmE}� �n?�c�c�͍�p��+C��)�u+��/����E����9zEY����I)�l����f �Ӝ��%��h��!R��t�2谽:+z,���d����eHR�Pԋg�p�n����X$�5�O�4aw��H&�!��nH�!/�o� ��4[f�L��N3v�Q���f��q�)�<L�))G�e'Z�xF���F���-�7����Ґ�Xz�i٤��V�k9QC�`ՅARѧ)�8�>��hV��e-)��"��/i�����#~�L��� ��e�HF?������:���9�P�w
Tk|��ahbK��ɚ0�C���Q��;���4Vԥ|� ~�����r��e",����*����/~Ի{פÒ��Q�4Vx~�P�r�g� 1���޼��-O,y��,w���K�,f	
JXT���_�W�+������4ҵ�JG�r�{�))L��K�:�U��goυ�t�8��F��w%���y�'akwHy\����C.~�q.֟��6f1kA����\�jފA��o���P��{+ENVnFQ]�ZsSmp2i��G!و@��۪�{g�?���i�k�t���%:ظ4��C��c³�"Up�r�y!\�Q����Դ�~�IXW��1�4N�SX륵������b3-ˮ�J�Z�HJ	v��>��i$*�����x���B�i$�:���'�$ʫ��F!i"C���� 8�K[XU�7M��7��f/��	��X�aπ�\�=`��ꝼ�������M^w�ׯ�:�h�l�1�F�zzk� �%4�Sf��j�m�x��aO����u������v�)H�|�9w|�R-|���!�2�V``�_���7M$��&�U�(#��	���(�AW	��u��-��z��*1"+��Bq�xa�X� ��	۶��&�z�`��K*^���3�;j���D���ȷ�qÙ�J��N��N��k���׹3�.�Щ!2����?�f>���xK�HY�}P��t��[���J���!����ڪx\ƤX�گ�j& C!ͤ��0�"�R�Y�	��lt؉�8�D�m�c�#o���Y����+Vjɀ�w�a�]d��l��%>��c�,�W�{L+�Cg4
����aC.�@�v(�{t�l|��(�T�o+O3�������ƍ6�g���f���9=v�6 �
J��ڭbj�YQ<�E*1&�F�����)�\��檱���l]1{"�(�0Q��½8w�Ho�qª��F'�O��dG}̞u���������[�-KB)���K{	�J���d�g�Pc��`@#�t��I+]5��7�N���u�Ʒ�5T�^Zz��mmF���9f3�O��Z��� ��������{B�(�Y�Fr%��_�+�M�n�1zN��6���|Wd���oY�Kd��+�A��>�L�o���v#H�o�ڂ�ru��ŬJ
���a���uwgi�e��@��R5���U���8�9AM'2�a��z��x�w�谡���F�"e��y���w8`�`cU;U��z�����ǭU�}�����?��g�E�Ϭ�[#�2�J6}Q���Q�\�]�7�*��}��5�f�&�Տ�H=X��F)�	���Ae�ӥR�r����x��[��b��3=�j���2W�����(Ϩ ��˵�{�����J�'����V��dȎ�f~�g�2PGZW$�/���������،G�W=�+�^0ae���hm{R�B� �YD���ɱe@�[��U��5GJ���'����)h�)%�ѭ��O�����Ş���hm<fz�u&d/�"�)��2D��"�>�p���i�".]��ϸm`�|�Kq��{�k[<+k���+4'T%C��N�k"/��li%#K���~���ǵ��N"擆�շ�F�S����
���u=�`zJS�p}L/-�h+�g�"$���$��=i��0�qq���syI�O;T���X�/K�~�^�R ��jk��_���$�-��"��F6��9��Sq.���?o7(�=}�4s�s�X�|̥���	�!�c�	{���>x���%t*�PI�CR����?�BSg^���c�������D���,�p
�q%Qu�&�<n=�R�~�6�1���g�-C�p��֌,��1��F[�׫R�ߺ�64��������L���7�&� ���M�J�mf+�ģ������R�w�_;bI�%;�Y���Z{��n<�c�k<߬�F]*�a&��0��dc9Þַ|�*D��� �S1�C�8;A)��S�F{��֓q��[�. ��"�/>Y���rèX���	�[�x���b���7��W�K9؍!��O�Ok��� x��͉�E#-+��&0��E�*p�iP���������>�����F|�M�n�A�.V�3�b[��5��PY���0�ӻ������tLQ���)�de���@fދ�\��;`xm�Vi�|�����pf���1�G�!ވ�t:5Grr:z�����j��u�d��ƈQq����2ՒPJk)%���~���ċq��-	���&�v�9�&�c��L�z��*we�G�(��Ұ���o�4M������i<�`�̅4Q���S��@pl[B�V�l�Szwp{C_ϡ}��5��
�������P(����y�̰��G�#�h5�F��7�>`R�(�Hh���=���xq'���\b���X��0(���Ƀ�(�o��CZ2R��u^�Y��T n_�bn;��W��.��Y�~��RS�ypI�0��(��ۺ��\�{aU��OU�yߑU��Xhy�g�䨵j�#�ȵw�_tT�$����>C���?�Y��[��+XD�H����X�˅CmV�.���>M�U�>�R�ۻ�#j��ʹ`��`���`��ws�G8/VP�#=�IN����)��9!~&�[�i��hq~m�떎��8�x������4�2΋���8^b����ߩY%�YFa�Y1�z�w��X�}|{#x�%�F^��ѱI��S綗�6�X?y�r��Ƕ/�M��X�7�l0�
By��o��<���6>�TD$�)�������:/�}�|A�i��_�VZ��2&ݩ���M�bp�eyIm=(r�BrȊC�%9����X+I�s(*@HQ��@�9t�\t���Jޥ�ېKf#5�}+#Šn���
r�ilPD��}p���:7�,)�t��cU,��aF>����
����"�&R���Rp�)�j~3���M!o��?�b�p�Fi�t_�P��N���w�.,+Q��bk�zp㽠�j�^����E�A?�i��L�������G8�O+�6�a�^4�,z�a͏�, ܂�$v.�d&����������@�`�C�J�l�OM԰�i>b����0�zj<iy�c���d@�Ϧ�,C�#�	�ZI�'O�(o����/�5���������Rf��Pp٥�����-݁��W�^�R���;�&�Ҥ"�3s��IZ�b���,�"P��.9�8�A����_Y�'��^55���g6���μ���HYD9l�vh��n�� .��QZc����%�_E �덜�7k���>�n;�'��1�|Z��BȤ�FV>j�����,>�h l���7��~�y{�|�,�h�����V<de�K&��M�JU��{��V)��V�,���/r��	ĝ�dp#���w|܏9��.MK凩�ņ)�@"'�#:� X�"Ќ`�;�榾�d�;<+2���G�/̽�%gģ�����,b��|kR��Y�o���Ň��q�����+�_?���:��&$�w-΂��B����E���?b�J}�xPI��qGF���.��O��H{��|�X�$��/B�*���&N�S�v�)��% �V��W	9ZQ1L��ZJ"�|辈���3��Z�l,�4�I��+c�*h�>ў�R�zW;�7�j!F��ˀe���z���P�D� V	\�Êf������is�/�sN�ȶɺb?�Ҵ" ��M��iWg6�����{�/S���W��9�d���#��;U�Ţ^,�n���8�_��� �(k�H`�(jek���tcs�8�[@4E$�����X|z��JF%p���k,6�PGx.s��:R�����ɧ�멼�v�K�[5���+��L�Ϗ���(zY���zP�㛕vr7G{6���������@R��flÆ��䞛�I.\D�q*UB-�c ~�>t�V@8C���:k(�����P���{��ɻ6���v��r��0��"O�k�)���ɠ��+ƌG)�Ţ�����(�W+3�� �(F���>�;2��M�ZU�7����-�xٸ�g�J��!\�W�e9]��J)����Obg�V(�!��r�/��j )��m�%S1�XG���������4�B�;N���LYf�ǉ�z�P
3r�;����-���0��� ��ѹ��R�TPV3���uZw��f�W�Z'�~ױCGΓ.���v��#�/�~/�3(��	߅#R���y�>�kkUb���ϗ@���}w멣�b���ye(��-�w�<ט��p�_�x~�Wel�
�WK���"G�S����\9�߈��J��{4��n9t���"�׵nXUxAǢڏ��|������AiS���X��sc  Bz(Ǚr�:N ÏY���$2�&{�(P�	3�Ҙ��SK�B�1�j������\��q���E�ex_cX�R����)?�?�r9�� w�-��n���O~���<�F�\4u�n-�3�7 ��!$X�w�<k���:1���
.�F�D@�Qs#��6ki��rop����+F�s)�n�F?�H�W�&�t~{H�{��
1	�Ū�LY�YF+0��^!EC��)x���$�����
����K�1~Y�����7��_z+��#���|�����i�)QB���6���|�W�K3��|�>rᗫNM-�=N;���]�8!N��Ą)��dA������9�5e�4�D���ǎVe��7��pw�X����-��7DP����4���e��Y��])�siy>1�����P8��цZ�J�z �6 ��qŗ�����4"��h�&c�-����v��Kn?�ԇ:���k2��{Դ�MY����&�m��@�j�2ARY��+��<��NP�D�`�5���{��1[�#��$/��(F½�?I��`�m�f��ǭ����Ԁ�`����F'�2T�O�}|�/�=��b�ex׃�u
�Q�k��R��k���������;��PnQ��]��݄a��	��	� ��y��4��W5@L���f_�G�8-�`4we�{�z^y���yY�cȿ�d3��Zd�ts�0�����l=�b O�Z%����� M+�����ѧ}� �V2�U����q��r,?�ܶ�L�7���ȣ"9cxpCY�����v2���8�$�����@��N_Q��H�� ����]Ƴ�
�{�42`�.��d⠟�t�q=}'�1K�ٿ�JP7���P� l��P?�@�Gȅ��F|E�SCe���?�BV;�h���G�"I�b˨݈��D���j�4���%����IbD�%`��jb�\iz���x�+��^<���Ƣ�wau���6f�M�>3R%O�^���<����%|V�H;�����t�Q�Dq�ٙ���g�M,�g@~��p1�/Q]�%�՝Q��d?��x>^�U5�@j�9z/�����E9j9����γJ�� ���{�Us�V&����� /C��K��M
+/��9q����7E�d7oK��� �64\6�g%˄�y��o�l�-'�_���/!�?a�ER�g�	C!� ��j|�o��N8zL���?�]i\=���ɾ~�~�ĵ�R-�&��D7��S��[���\|�&��3�g��9���*˘�**�z�S"����'D��6��� ����B�5�*c@�ܾ]���u�d�2Y�64�w7��C�5/[�U�)����#`?*a.ڦ�e0��:��W&�� \��U`rp��u�z8x(�nԬL������E��E���d`ʊOCb�tAP�(�B�V{`���|��wIʨ�G"a��M���#�"�$��Q3*_{P�}��?�4� $Xb~�I��Ԝ,��ʬČ=�」}����#�#�v��)���]�t:�+�k:������5��J���#�up�PI�q-�i��؎�*�J�eV���B��N�Y�7�Ӯ�B&)۠N�>��_�nS�����9AELK,�tB1G��)S�j1��2�C���e#�Wɒ����a��E�x���iD�GG��:T�2�V���LƂ2w�V�4E��ӇX�8_CI/��E��iݿ-�0&�StO	Ά���̝�&�4Ʌ�J�'�n�������e�acrK^b��:w# ڀ���F��a=&EW`��[�YJ/�*V�w1�d�l4�r������C�s��F�߃�a`|}D+e{��̑d	ε/09��Yx0I�{>��g�Myj*K��ʹ���G�O��،a��� �����Y�Ԉ�����݊�' ���ɞ������Zir��c0�+������Cj��Z1y�~q;��?�yv/��I�9��F���F�R�{f�>DǗ�ڰ�@ӟ��aި�G�y֋�d�[A�X��EY��/���R'?('O[�}��4gy�u���$�����O�� V<f�
��-��єT	ۡ���s\.�3__��y>`�9�dsp�̮�Y��Y;��e�72<
��l����M�w��C���#~�G|�s�vV��P����6�[3w:O9��`��Ǭ�7$"��1�e�e&��9P�j2F|Q�aVlVף1Y�
�i��9���|ԡ�Й�����~m�q�4�Ҧ4��-Q�i�(j��u�sͮ�$Ăv�ц�W�}��	+�0YYdZ4�и�6�{���5�-$�G�I�����܄��	~ЉQ���J�P16
4�����v\���$��9�; �Z�l�(:m��H���d��rK���	��A�E�!?W4A���Ҥ��z
�)*�K�;�`B\��,�B2���[��?Q��ʽ:d�i�w�����܆��ˋ�Kͤc�����H�l���b��J��?�����y�	]H�xT=ٳ��r��_�ش�E���7�z�K�Ν�W� ���+�01,*㏀�ƀ|5}�zWW
�z���"�<	?z�t����b��>����	O)t���1���͐pz�蓪�V�+��Y���쑀l�Kx�xQ���� ��4���r5��TC"��}��E�vw�΋CasO�݆r�
R�Fq�JM/`�Jm�[ ud$p�%aKY�.&j�oQv��xP�5�g�5��4U}�S��#�M���q�1�B�\{>#�`⛂R͕Q�l�������i���jj�&p/;�����۶�4��WB�)�G�9�-�f�O�z�d�W\���g�W����p����kGm�"��c�18[�xc�}AUǙ�Jy[hR�H�3-�n���'t�c����>��8�Իx{b\��hy���q�\鐲#�H�$�6��<��JʲD��j�����m�%�E
IC��KW'���m ��Ոf��2<1܋��g��~�!��n����Y�#�� ���t��״�)�j�Jׄ�6���%F)�[[�%���YdcC~��W���u��iL�t��ī��3��+7��"*XEQ��hF�n�iUk��Z���k�~�11v�+4圶89@�����^*cii��c�
�[G���M��ָ�cS`��?�_����Z�d���5��lv���W�!�U*Դ��Ȅx�Yy���Mlf�����}�ƅ�,�]=P�R��W'K�n�YH� �� �����z��]����n�K`�=�
DQ�,��s�B��V�~3�y� �dR{����� M8��;����Y*�ux�We#�B�'mei�e�	GS�0��f�L`�0��j1T�L�nj0��~�5{�����7�yR���Aa�����5�ڿ��2��L�;�2��-�t=́x�Z�����0\zԪ�8zFY�/��4�}N�k�pA��'/���eT,No;��~��m��
�X%L�
u���b5����(!��o�v�I<9����p����'v�B{fk�ȡwK�����NB���8Cy�w�֦
��p��7�!Q*3^AQ^c�v^�[A}��J,͢YǸ5�I��"w��K�$B*h`%w�t������A��I���!s���Kd�A)��ÍE�uA牏�ˑ=`��`�wK��h5At'����@��u�dY�s�h��eP��:���O��LU�}b��9(��Y�!����Y=�4�F�D���AL�j��Xz��c\��r%����oL�C�'�4���ĜŃR�O��a
�?y\���NϠ��Q��캎-�@Q,rg	Z���"�t%������߃��7��<�=� �pe�~y ����g۟�/�����Ev��e������UV_���IvT)�Ii k|}�Е1���YԄ0r���&`��N���A`�] �۫�_��@Ǥ�	��|��8�_���J$���Lܼ��oxl�����g�45~O�DH�jQ��2���.�z|�*�Ku���ƕK]U`���Q�@�ށ�<�+"9	$1{%&�Ћr ��I 
����1��VrkKoO��O�}�[����C�~�۞�l<k<�9�)p-�B�D�P<�U�Q�A�o���a#_��0��Ƶ�1P�OG��yC�t��z7c%��iʙ}y���/`hJ�e<��&��|:Km��	%Ι�2>����81�����U4~�_1���_���6�\=%���n=5ɗEs��OhL��fD%���8��˳-�寬��04�|�B�-{P�v��8C�3�x���.l��������n���\����ژ�3�	�������������V7&�S��5gU ��-%��N��������.϶�Q33�Y�e����6���A��d+��A�0�N@�ʠ�r�]�"7`����ȩͶ>EZ��{7bP!#��=:&"?I���!�l�B|x��Y�L3��W��uX��7�.�)
+Ѝ����V��˽�"���Nl��[���73C�lX�︛-����a�}μ6��C�m�@�Pypو�����4�g�.��jFL;����w�iTp}̹0��1�g�m�S�6��_�Zg��"�IɆi�4I�k&��K��x�_X#�1�UN�D�>����F,}$|֘G��F���XW�q�H��c�K_�|�E[�%:�F�l�=���7�����X;���$��T�@�g>�;%{߁�nKM�ה���;�y����i ��e. \40s�����b��\S4(�;�_JC\:w(���&sR\��09��J�5Fc����rR�9/,�L�$��_���e�6�D%���r�BtƉ=�xF.��Ի��g�&~�����Q���u��i�T�[��1q�I�fkW�&�d�������՝]ld����0
�Fϟ�����p�ϼ�5w�<�&ZhM�=jǖё׬Y�v�_��:���=���a�!�].�m�y�6%T�(�.���5�x/���1Dc!-=��{Yk�^����K�..i��=�ͩ��y	����V��ڊ�'��J���,IQ���r��wv��m +@,v&�
�;��B����N�4��{ �ϟ���M�=�o�Q ��7%N��d������H�������y�RM����_��p^�
�k��(��F��ö�V,7�7���E��N�Pi`���Oo��Tc-k����pr��K78z/�(���gi���9�h_��+�kw<�*ՙ�g$%���cc7���;@'6�����쪈i_�4Z.y(=�-�k���>�2�����0=V�G�5a<8�&k`	�A 
81��i�Ǎ����,[ -\���J��9D��FKn�1�ݫq�����0}��mv�uY�F`u=�v%.�3�ʓ6�w�������.Y�WA�>��Q9[��jeY6���G��=:w�7��������%��/6P=�8���U���)��-T�Q4l�M�e%��x�&ʎljk3g�{r�; �b��g�Rn�Ğ�Ӻ=�)�FJ�u��u�����8�b}�M4s�E�#�%��}�vot���G�>����x���Z�Џ���S�	��%�����/t�MW����v��/�594���i�p�3F��9�n�`�W��Vp��ua����=-H4�c�o�ň�T�H$Ў��>d\��6	�֢a'�ȾK=9�'���'���#,���a9�ZB}����)�I�UZݭ�K!<�ʵK,�k��ė S����>����#��q�]Si�� _Rx��)v�`��U��k�Z�	�_f��/ƿ���� �g�=�\/U�&e�X�C�ڋp��p2��r@?�����a�Yȏ�*��*��ơ�ų���xd��7E=�qI�����8v���ĝMmB��kʇ�T!� �r���x�ǧB��^�Ø�<r���9��#���Ϫ*X}G���ϔ�#���	��0#r`����r�n� ��<g�9켈J@
�C��"3���5�j��Ze���Da�UC՛(8¶��f=��|V��3�'�G��'kK���	
퐟^�q�tP7���!5Żx p�W��T;�L��1	!J������K/<F��>�b��F�}�lH��l7�R&k��V�5�[�����랃��(�PF~V(��{z�h���D� ��5�P��D�؄�V�pa��]�xr�W�Ֆ�8��M�nF�	M�4�	����B��Wd���y$Q��.d�?��z�TQ/L�9($�<�	g{;tW)?��uf5�i@��gۏ0o�5���kCe�s�,6pW�/w?�-H8-�����g���8�Kx``y��Y�S�BE�� w��.�J��ÄX+�y���=ka�&՛��ޛ&��Zg,)�������0�$ŋ�?PN#\>�9�U(0W��񏉫�*�v�uS��<�j�^~n8&�����N�\z�7&b��b�~d���#nm!=QC�9ҿ���r�j+. ��'�J����|�H�G����W�O ^�)�������ڎ�!`�-<�QVUl���8�zv��F����=���Q58Nv���d��`]"�oL=p9f�"<�\.n�;��2���n������X��Qk�Oƥ��8N'����?�;j�E�� ��� �@�h�ӯZ
D���	雡Z)������~�Q�h���3>kB�Q�IX%C� 	EP�X�.Tw�t�]R[$^�ű<���q���Tv�Xq~uL��tg�Rl�/�G�	3Z��^���bIU 1�L�(�y�1(Y�V�@���K���.o���lJهZ4J���C&�+E�>�M^A��W�7���O�#��״dO�?C>�M���1���镳�Df��(Y�*j=ۏK��OK� -�bB�Q:�lO��ސ��CX�%-q������@�,ѽ1d��.��+��ӎ���Ƈ�V)� ��J�GD���@W��""A&(�!�%��>&@���@�K.���|�\C�āS�%L̡t�VH��{:rQ��#��%6�53����M�њ��r��֘�	���o>�vʴhlG���u�x�0��:[CjYв���?�l����ճ��r^�b��11���8���r#���e��J����s�� Z��!��m�\$/�����SBbϡ!d>���݋>m�+8b��BKj��w9F�p���fI�7O�cLTc|�i�e�,�v@�*�u/��.V���d����}�ӕ,��8ۼ�.��bt+����sa޶�L�m���c�Pq�P��c`3�����W����&*��Z�#M�;��<�(hp�@�������L!v+{�=�X,����H��k�t�+Ί�җ�k�
 6��
��*-Ŵ{s%�O��׉���i��~l���j�g��'�1N`>ez�ڌkW�qĨ@U�ٍ���W�0_i�=�Ow@���QW������ݵ�`�����7e�Y��ΐ�5,�;�:��w�΋Aj���$�/m��pm_<��fL��Abhw�ܤ�d��9j��v^�dⵙ9������H��l���ss��6�ۤrl��2l��?{�B~�|ܝ�@Y4�s�qo���:Ȓv\,E*�"����0����N� ֙�'��+��7��TA�b�����t�747�jl�֨��t�w���BZ�kF���W��uDEV�
��x����[y�#5��/�7���Y�{Ş�����7��UIW���]9\�n)58��ʅM//O�+�P�":�g�Hu��`����n�=���SM>�TvaՇ
��9��s"\�D,�pu��J���9uRM���������zS� k�5ZL�t7>��Qd���̅�~B�:�9B�YZ�U�;��p���K�з�X�kj���'�^Z[�����K�Ulon3�axz�cסd�!���i�it���i%�#�`ܟ�uF��5����4�Y�qf��WV��%hwzI��wymC���/�A�5��!��}����w3�6���-H��m��KLL��������C7B]��߉6�X��6�(�lȦaC�Y�]�2�2�:Ŋ��C2��0_�����92���m򰘍��Zʥ� ?b9�Q�%��J�r�ṳ�M�C���zoI#�Bی��*⓲�l�1ڑJWMhl�iЉ��洐#������_�ٖ����7r'���N�!�̀t���J(�]�����v<��wP_�Ќ���n���ח7<���4({��4{�������t4>��c�Y���a�3�l�:zM��S�}�(Oa��Wo���5�_�wJ_��j�֏�#� l7\�j����{2$�6x�j^�l�����)�q�{%��RB8ξ߂�L����y���}
(p���I��˖2���t��h�=c�䂘tk��G�<�oe�V�!졅�^�5��"��w��T�o F1�a�4GL�e��@h*IX��1ְ��cV���)V<н W�Q���C��\-���j5�4��$tƹ��L�&�-y��U֫�����zj$��F����MQ��栟�.WV�L�d㬆��ۍ*�
~�EG�<]H��h��m=�$;
^�f������?5�A�tnML����
�Mȩs��״g�S����.R.]`�y�|u%3����<�"ִl��ބ�U�6��%��l�UgK��3�_	FK7���ޔ�f�$E��]+��+�0�d�DVG�����#����3���t�0&C�e����j�ƺFЀ&�L���	�f��i�ErK��П�����M` ��İ��É�pX&�Ɗ�ASؗ
u��ɐ���z�U��Km�Q������<��'��|��~��&�챉J 7�n����,�IJ�UV>�;bn|��j�SV��D�D�ύ�PV�rg�장�f��;ю^�~~*��h�]1��%%X����^�Ͽ��Z���&�EW a�Y�^����4QY��nq�}@��r�c�<�ɒ�e���(�r�ő��=�$?��>��X����`L�-�r�j~A��+a��6}����;Z�`O_+%>F<�(\��b�s_ݱ��������I� �r��H��2Rdm��k(m� �w�3hW�&�S�\�X8|u�Lf����@�%�3�I6�*@%4�5i�.��U�@Rp�Eܢ-x����`G�!}{���lJ���	��������l���c��Sz�
�C��#P|/�Xi��k_f�'8_mJ	��'7
��7��$R��qA����_�dc2�B���I�-O�$��c=h�(�ɪ%#-�N|�#�$i6�lK����&ȦxI���HvL�ɬ�"�
���?FO7{���Y�3�:���hT�V�<3�0�+'e��׋��~gv�4aFzP�� o�/�[����J]\���/�#������y�j�6k�~m�VQ��?���/g�6�E̗am쥷ve5K�⯲0P ���@�����0��A�h%WM*y{���1��#�4Q�Eb:�X��/��z,��zǾ�v
�(�?�� oB k�p����)��{����:6��X�'f5��jq�)� �T��""}���qn�e�����X�Pv��
�X�Eg�띠�=� lmVM鋤�5��=�Y���TXlZ�c�
*"U�ʻ	��х�.��
x��`�_��u	�I��;�B�pt��2p����6�Ӗ��2T%Nٷ&����|r�`������œ-.�Q��-fHIl0;��zϗ�L¥$Ce�Ix���?]}gu~���=U`�k�%�$�c������6��7�9�>9�iWQB�����
R�_�яV"2�u��0�։����φr���2�"�tY7 ���U5�|���]C�g�Z1k7�9gY��D��J��:���O۸Z����Vvȼ��D�D�Y�37m�L­J7C�Y���=�����%2�T��@C�H4�o�R���|�ٓ�NP��Z�D�u��)�?���!{rLV:�K���s �ڤ��~B�9���v�?G/�0���ے�:�?��6�e{h�;���8�(Z���o�ĈN��� qU3���\��i{}��o�J�-��G�|�/A%�i'w��wĔf��T�smT�ɢ^W$`5o�O�M�����»��$���;rϺ�߄��S��𐷊ϛ�XV[awRB|�;���3+��=����+F�v!��P�3�/���ޱԙ��׷��20�ӵ�[�
���M纻�f8�S����q��Q��'VfZ�#����۫H����lc �iI�P�S�I䣊Pz��^����r#[aZq��mv�!(r�4@����/�=�0t�H������ca��=:�VxLR`��ć�=�	Al,��[�	R��c���v�S|L������U�Fj�� �v��0g ���~,�p�Y|�ذ)��Pޠ��竔�if��PҚ��5Ka��`GBo�cᆎ�	�����k��W&�=}��!�0!	V	8]$}:����?Z�!��h���������F׺���Ѐp�7=v�����|�����i?#B�I5�6(KS�3�js�MXX��S2q����7W�4��	x3��� �:Z|��0������N=d�%HL�X�5s��1��l�����'n��C�_���m����m&�S�C���<����H�]�1��a��ɗ�}g�ny�h��(A&˅pV����%)��ҰL�~4$f���f�/�>v�9�^�Z0�0n�r:�XF^����b���#����q��m�[J����`�{0<-��%i.�=+��'h/%���Ñ��l��׽��3�Q��p5��f�5��:��ˡD�3̟f~�rk"Yj��5�R��׀�.�:�o�7���$}^�}Ԣ�^�ߜ��MÓ�9�F8"kLP��-,�
W�
^]��T����#���]�ɤl�>+�{��J��py�]���[Q�Q���>ة������}��A��(�tE4 � ���yG#/5w��?�&1*P�rSl�K���v�Z�В`̶D���������v@�XY�(4�u>>ml[,YkH��Ό�Xg�	��{�r���W�hR 4v�s���7��0�wI?p&\:�e��4�6"�}k�V�j#7�8Z.��u��vG�����g���h�;W�R��*��pk;�)8S;ƾ~��'��B���P;�'�z��Wvڦ������X�(MSV�\_!�����,���Pkg:�W�x,��
\S<h4<x��;�f���8]KiM��9�g8:�	��*ִy}���M�5�y�=q� 4��s�	�(��G�ʒ�}��Ɡ���?J�Z���W*��CWِy�!S������>��(�%r=+N����`���Y*��1Ιᐍ+���uE��-F��#�k'�Q�q�	�N��D��������?i#؁W;/-(~��5j�]��n�H���i�x��G�5�S6���@�|�`�%� gI�F��ܯ9�8@<&4�Yd�κ�Yٟ=�#U\���_�tvM`gX�#�Z>	�+:���)�㿒����_�k�ױ=���F������䛟(R\]�s�1�����jcc�^�s�������C,S/c��0s��QBWq��8��|Q<���2~�lC�Cv��R@\�N!����?#͵�1���#:0Z�9��D� �������<�zGx�,[m�Vk��Ub�Bc���z�QR���s9膢� h�$��o�L�#�8Nu	Q�`�n�|$N�9�dz���}�΢��Y&S�<)�3��a�ϟk������`�N�<�	��,�r*�Z(�G��	���p�J�#O����˲Ed[E_���a�p�$ Ǹ'���v:aZ��\3��p�1д�'�
���6�	�ל��Jox�����O�B��흢b_��<g�g%��G�#F�A�?������NG�@jF@=�{馕��֗����:�9��X��M�I�⋟m4��˻L��n'��I�g�.��Й�������Ĉ')�x��՝2�I M�d��mٜ�Y2����j���C.���TB�.~#�p�� �R��)}0]Y�}���{\��2�y�};O�9I�*t�`;ny�Kn�Af����E��!�Ex	A_ה<�;[���4a�1a�ZF��R����I�X���޾ �$�<fT���q��ߋ9�u�"�n��O�#g� �˅w�:��Č<ݪf�"k�g#����>�&�L��J�:��YD�*fP6'��/�p���oh�d�KQe�<�RD����o����Hx�S�~dĪ(���C�&�JVh�g�>���i4z���ߝq�ShȯZӯ[H�q�h��)��JJ�H�1�I=e�;%�d99���/�#G�1���Լ3���	L%�\�s��(`�n��a���w�A�O�dA��X�G!�p�GE�T��V|2��|��`�\�P�d)�ظ�(H�����\ABO�`�9Wl �`�s��pR�����Ԇv����=0	�G�m%��aG���Q)4XFַ�>H�${���}#l�&xc��k��Ͼ&eͲ��b���J|���0v��6Zz���2�EX^ :Y�+�p��,�m�KtSnrp
;��p����HnJѣWu�y �P��Fx��̿,쐍���6��uJ��*�DO�SV�H�.E���sC�pō�%�0#eE|��0�I8Djw�u٠��fK�?�Lx����˧���2M��g�(iK5ol��Z��w��;x6ٵ�W�����Q�x[a�񤎎���?��L��?Z�c��V�w���⣸N�����-堭#'eϽx�! 5_m/x���j?n��m�����@}�񝋬-9 ��l����t/b��ކ��Kd8��/Qd�6&����|x7����mAS�kKt������@�(,j=�Л��ɕ�ץb���g�=�j��-	�nz�=�q�X��/��<l�xF�_6�'K��m��Wgۚ`U�[�0c�:��l�7����g+���['�ԋ>
�aѴ� 3K��-,�MIu.?�wؿ�h��fj���ag��%M͗o<��ki#9�pU�p�m�h :�q�t{YZ:x�Ȧm����fr��ss���
��<��8F�l��^sﻜ�=}@�l23��{ܕZ�X,�5�|"�>V���Ϧ�˶	�a=�k,�@��,�ivLN�B%*�3�����$�����yW���]��'���Q}��ϼ743n~6��ݑ��YiG5ߡ�36)�Ƣ�/���l�´��Ń�v�;�hmDƾ���Y��t�g�f��N!���j��Y4,���{��H]�Z�l����X������z�4f
��X�^����A�҆��n��G�8�%�t	��
q%#��(@-����������{�x�:A��-j���]���b�-H`�]X.�^JT�~�ρݘ���Pz3ס/��7�ʌ	���ֽe�&HX�N�#X�O�\�k�<�jD�=&�ڼ��I=ƈJ,��vά Amc�z�A��uw4�
M8��TO ����� �^�z��+��(y(c
���4ǽ�?A���ϊ����
���2|԰�J(8N0���ϧ�/��ʆѪ�Ɩ��,3B@��/�ġ���h�O��ko�N'�<�hvM�`L�*�E���<���M<-�y1 ��ҢL�ل��9�aL�}cAh�o��:�[VI�����@F���ʬ�`PD��HíV�c�ܸ�>��8i��S������c&��}t����ȑ�n�G}���E���Sv��t��)����f���>�(�Г�Eː�C4��C��q������ҐpW���������7*M:}t-):���|.�Ө�<��L�!�a{=tb
��>EAR"юpA�I�gv.�x-Pl�3�k{(i��q��N޵c3��qr����hO���rq8K]M�D�N�9�"��x��?m���Z�ñ�S2��J��0Ѯx�K'���E=�yz8��p!a�����.�!A��b�^�"�4�֟B��x#7$9'*�x�rd܆�ש)�x�}�6�C�.刿&��;:��-)�G�z�x7F�C���	A/�X6����ߣ�A�j��\J�ɿ��_�!���Q�[P��d�
 ��R��|"+�o)o6�)����V����y�Yv��Ԧ��~k��I�Q(E�t)'�i�xN -�C�k.E�2����buV�����0c+K5Lݰ�&���
ײ��Y<2�G�a�ܱ��%���Y�)K�D3�j��i�%�����I����b�<�^�$�hݡbk�+���ߴ`��4�o�Iy�[(��Y��dr�1+�I=_��݂��_�뛈���[u6���u�^�� ��)媋�ѥ��:�3<���]�I�Te�@���^��ퟨ/|&��8��0:ŊQ��t���m�:m+j]��1��_��=��O*�n�9�~�(��;��m�pv^,l�|k�q7��C��$%��[j4]�La b���(@Ms��*`0��Y��3E�	>ڰ�bP(���@���gn%s�Ѯ)5���<�Ќ����f�����d���o�>D�3��U[���P�]*��I{H�~F:�_j����������YIz�d������9�'D*�N�[C������	�����o�l���O�����4)m��p^X<sM0�ձM%�5��"�4�?�����1;���~J,����xר���m��m�:N6���}�b��[�$ #���pP"��BO���8�s�*̏N?�J���d.F���z��~�e!� c�/�,
|x�נʨy��u~�w���&�%���]���<��Y�Jt~�������	��e<ƞ4�i��C����j/}�`(�x���<�+q�*z�r�I�/�.�c��O$����q!��WLm(}G�
�P{�9�TQN=���'�@zW��^�}��P�԰����w�Ѭ<�=4dZ][�;�n%�����˼Z�uR��h��Ĩ��˒f��*��4ӕb_�y$R$���a~�h]�� ļԔ<��� ��zz9+A�n�>� h�<�J�ŭLaPM t05�s���zs�l�����S�AJ��������9Zɥ_�g�Ik�Q寵����͍�X��/QD%��-� �?�w�86��zYѻ��~��~5�lԌ�d��3#'�f�X��T�AcT3i�3f�D����݉�,� -.m��TyqVTr�;v>Թ��7<@@:m��d���⽢@���gT��y�{�����gϖ<��&$�î�l;��0����a"�Xv_�*s� ��8�tnA7!�����5��g����\\����o�����\/�bQ���v9��xdDa��pTm��LDZ0�N��tw�x�`�_��U���Ϣ��Y|����X�˻��
0Ԁ��u��|�d�ǖ��&E�f�P���X�W뉃 ��L2��O��.k|��i�P$��7<̀�h��P����[4N>���k�@�ؕN�k���~*�+�4,WV����o�Y����q�p3�Y-�Zh��}*.G��W�@�[o&�z��Bm�����|xW�Oh�D5�\��G6̔�}�]�|0jZ�Z=�j��ХB�S�B@X|9X��~�e�4���/�%wf��ќD2B,IH�U����z���Z��js��Օ�(�}�x�]'U��%|�9����;�Z�កl��J09��I<'��]06�����.Pfq�|AP]!c(���}�L
����g�B�;���&�G�z�W�B��p�mG/��2�ITa�Zgw�%���-�J��X���D�0��qR��'r.WZ���|A���J'�߁?���0m�a�Ne�T�Ə��;r
§��ضΞ��P����=����⬌d���:��A��Z�{�S���9���0��5Na�(ʕ�fNwx�n_��5�H7���=oq�3��������-�齅ڜ������7_� H��֊\"	�6A�.5 �85l��΢�]gcgn��Hmm�',�6ַ�{����$��-�'���Y][�ϥ=~72�
~���(��u��lF�<[	]#!U�j)yBP�����a�q5��T9*_�ew����˄T����'T2�:|�Հyjm_Q��)w���_9W����/.�P&D֕���s[���$x���J�1I]�rw5�����k����':��"esoW�6~&4b����PGͺ�Vk��/�����.�pHOt㊛dm;=Q�ں��)�D�5�
?M���ꈾ\��Y�����U��'N�B6������g���9{-}�G����4yX@&�r�D1(��V��VI�f�zB�?"����1�8�,)�u[% ��!��v!jԉ��|�B�Za-�4xg��S��
�o������Z�����O߄�͚]ue
3���B�Wm�I7r��@5�u��,��M��i�Ӧe��,�1��� �,��K��$��1��D`9�n�Z7��g�;+�%b5��)���d�G�9�5ڮ��io4˽����4�6�gi�{�hg6���j�׈�l	%N4��/[Edd����lHK�V{Y�q���xe��$�ì�,���5���syg��S�C��)M�����x�x�Q��+^{�m��_�'���� ���1�oO~k�}��FK��07n�e(mH�Kh��6�>^�v9�T��T��:�\ 
������w������'Ч������f3�@�(Q;Y5V�:��\%5��M2���A��f$�  u�iȨ�/�q�	z0�e�o� ��0襕�wD��!��h
�$�c��7w�.4Kx��}Y����p�vt3�r�d��F#]��M�U�'{O�I�;�;~�ȠTz_�����0�UV��<�g������F�n�^�����.aQ��ݳ�"9|��o|G�v ����u<��F�K�ϨĆ�$�&	a�M���(-S��w�Jp�8�a�,U���,wN��=hŸ3�o��*>$1Vn��٭�_�.�$ػ����kP
	�*������S���C�Z(iȊI�8J.��9Cqִ�~hT���v�Qo���ϱ�s��V	;�pC�3���ɮ Y�{�݁�u�1x\� ��)��?�Օ�!�2 �� ��1W,�/	eTN��M.6;9��kI@?��$b��E�4�OKՒJ}3���N�T+G���w*Ē7�0+���u�J�F��0��(J�:cz���ٗ�*�#�}4aԉ b��:��'��4&+BMtY�N�YW��1���@.��OTm߾5�v]�AҒ�12��u`{1���K1�D�����JkٓHa��.&��bd�ڇ;��AH39 �����cb��M�dR��4��j��{²��J�"v�.R��:�c�;�곴+��ɐG::�c��ܯP(�My�Ϥ��R��}�ЊZQ6z:���pD�d��W/w�
5�n���h��V�If�&3�Xj�Ґ.8t�ÈGW��	�I�aKԩ.���p�M��L2��p�=M����=��BS�R�^C�����y�ɫ2X�5�TYr�,fd�s�_�=�����73d�C��iU���O�Z�qGg|�e�W��
<㝤�sy�oC�Ù0��K�b���6{ӒC�Ǫ� �Z%<k�3�Zi�.E�a{Z��2u�WJ�]^^�Z��p\��:X�L�'XG�qjq!����!p'�s�B������99��[a���j
�����bk�Ϋbf�4��a�4$E*ݍ8�5���7Tq�v��E���7�9p�M:���T5L��1�����)�o��/�����ܔf�'���l��Ý��oj\Ur�s�O�y���p& �ȁ�nX,H��.%/����(��쵲ϳ�f'+��4�u�[���L�NónA�Q(Y'Bc��+Z�s2m�d'2�V�R��:�6��$�Y#
=$��p�F��O��,O-�8�w>&���=��m)lf-�q��,+�A���`�Ϩ2�+�ed�)G�Ζ�p�H\�J������f��}�M������I[-�z\B�O�AA�ۍ��P犜B�I�&�e��]AH����+}C'����^��
��"���4��E��`�]����
l��f��"�����Ʀ}���kOڙ:��yS�Q�V�$����Y%8`�i6��T�$tuZ�]%�@4ƃ���!T���5�ũǥ{�Z�p\�kZ��q39�k���U�`��٨����\"J9�a�7Ϋh�zh��U��4���s�)t�X�����mN�_���f�� Hw����Ew��D�&u ͱ���䘳S�3� ��[Y�H��p�!�Ə�K���'� e�[/��o.)k�X��bw��2�t�}里6CZ&8�u6�=}�#�Z�k���g��ׂo�kΐ�!�����|��-g��I���<�������5|�h��/h�iʹ���,�
Tu�ۚ|,��cEX~���Υb.rc�h|���&�x��U?���ߩF�C��Sэo4���4�	�$��ι��V�7B��4/1���>,��F��[��D�C.u�6,� ~��H<?[������`s*Cr�8�B�.�f��؆RbR�li�f|��0=���pJ�;�yY�`��^O@1�]�X��:�N�>z�/5{��(�J}W!W<�W��0���̑E,�P�,	Vsfq�Ӕ���A��.U�d�g|O~��&�z%��ߋ1�4��������m.�"ɽ���Ո��Q�mH�TA�/���o�I��	"uYWD�^��7����h-+Q^$�ז�C�{	*"���g�-��A&�Ar!����F*w¡;�>�K��!�י�9Q���B�Z7���Y�Sm,<�J�>pF��(&?�y��(��q�mG�>Ý�BY�L�ǓE�#cT��~���H֚�����\�M<t�ShpG��0��Avp��g�Ղ�	�r� ^�t9��Eݼa������q����8��5�䭌�f[�;iNU��څ�]����2����Ƽn]7RɃo�r|炒���Q��S@�b^P�  	�^�Y��cM)�.���+=fx'e�7�7|�uw^�x�Q��&��L�اΞ�,�-�"��� �?���}p"q^RP��
AP"	��b��b?F���N���p��G�M��6�7]�q8R5��~�JjY H!��Q�z�ͮ<���P���]���1}��|��S�ò�E䟧���l��g�?�a��X��gr�����L��y&��:RߔL�L����q�&Y8EQ
0d<d�z�#*���IDQ�+�'���6@�����/�wn�I�m�JGub�(���Ρ�i�x,�Y2��OM�B���].B{E���6���ڸŐTDUm�E�͙x:��"�Q.��?��؁�0l��'��=2+�����Ө���n��5Uc!= \�(�B�m�zA��ڨN�{ݙ���@s+���E�}�xP.F��r��;}XK]��e�5����l^ ;�:�?�-@M�h;���CB+��J��<+�}~�z��O��~�D��=��Ha�M�,�̦iēĬ5�"���`��;�(���b���6IM����H
� u�p z�.?�)P5[�vJK�'8B?�^��a��ݿ����J��I�����\���:�`%0���K;���hR��c�0%�`/�8��'P��п�9�l���W�q*����W!0ѯ�ŏ��V����'zgo�}+��e���B�/��y��k�d���Y�I�&�9�xW{�i���?M�z���z��I^��L���F��!r��$C9X��02�J{�
��s����\�n@�`qLF�,6���Oi�r�;AK�Ӥ���ia�!��!"f���6&J9U����C�� t%T4I9;f���lU�潸jA
3��E�B'�VU\����Nd�PҺ{�A}7�{Q�G>W������w��Lٛ$:�J��>+w�`YZ=<=�#�k7�l�!�X�vO�.���x�H���`^��1���v�w�Q�n���J����,GD>�Y�㴲^f1Aa8"Ӳu�:s��	����W{��Y���I��It����T!�mZǼ5Ha8w�>�M5���a�R� �VW��4�6��`�$�k�[�s� �/��l�"l!��!E��Fk�����6 ���٘�?6��'�Xɫ8�4a�=�'�-��[�Rz�C����g��Ux@lм�+T6]�����;�Ɋ����Z9:%����m�T�Q\,��[_ߜ��y+Һ�l��i�5u�ӈ�`a��*IA��l�I���i�k��BS���}��?e���]�-G
�bS�����]�{���ڶ �XSH�k���ggɖ��+�ȅ�KJu�����5��m5/ǖ���5z�9��ZnP1��f�}�fB�@�UL�n?�׀��ů��H���Y��q=�<7�i_iqա��1O�_M�o�yJ}"�����
Qƻ���q9FQH:vӫ����5{9���(p��ޝ�!w��t�H�7qd��1s�uGrk�2���O��o]�/���{�1�Fu�ؾ~*L	����6hV%G}�Ҧ-º+ss���������Zf� �X+���G\<��G��#��Mc��Cu��Ia-N���l9e�F�ȝp�.شSD��=��Y���y%dak#����x &K�=��ez-Y��N-d�6㗲�������A�*h�u p��o=":t������a�����y�=d��~��jN�'�}1S���@L7i0����ߐ4o��x[��y���%��C�v�+���k�������C	:�l+b�����1ǋ�Y�=u��M��p�.�<�������q��Zt��$��K��L�Y�>�<5El�>��b�'��%��3i�Y��$�(H8X�~Gon���/e*��a�:�$q�!��QR��S����U�2n���O�>kx�A3�fs�7X�B	��*�(LfC����t��L_�0K�xV�}��F��R?�����<��`jI:$�M��A�z�n��F�P�A����/ں��g�"���N火=��������!�
�9�Wb+��:�^�m�XkI���(���I��)F�H��&�aW����{M�y�H0ݾ��9�J<�pjc�5g�0��6�z�]�un���]#���P�?:>���oB4�?�5���(��`>��64���ȹ����K؇��$�$0/j�sB�$�-_� J��;��nO*4�>{w����0"��y����P�S��p7"����텓t����S����vE�s3��m�ՓY�}���z%�c̢F$*C������ty���<k]����c��]�VCh�'!+�֟z*%T,e}�EG~�ʹMun
�4P[ų��Z�`�z|m�j�Ւ�f��Y��]���m��u��}�}\���Q�q6�SV?Y�������O‹<�Y�ۉ����hc��,G<!d� wK���:����V^���E$��ꌭB�˶�H��D07����ʄk��A���ko�\����x�����~]� �=�v"�XNz��>���d���k��F
ƏL˳V����/��ۃ�sp��3���0���"*�&����'�e�j�z�]A�;�])����#��P�e�m��l���,u'2ɗ*M��ټ����"��ȊA�OF<�fil����w{�,�9}1J��!V+G��F��^©)�4!�#���oL2�/����|z���z��a5�L��&݌˟%�u1��.�2c�K��p:�*��'ڷ^���n�&�U%�\~L��h�ݗ�ˎ�ۉ$B�j|�(��\����SS- �����vGi�ߥ��)M�U�������m���=��S�<r�=���L��o�z��ͥ��ơ�D�?����&K��O���)��F��>g"j��t�����h�Gj��O.��xiT)��n$<m��#~�g���m~�?h��V�HT?��� =ĢFG��'���Ww= 7+& 3�3��@�~�~z*��s���1[-�1h�z��
����a^pL.5�yvA5��3�BP���9f��2$��^H0N�=�3���p7�1����&��2�p���+E���̡��#R:�R�Wn�O�ǹ��r~"��w/o��*3�GZ�
���#��x�:<���,,��4~2���V:Z��o��4��엪��p<4�pi����Uf�|;/��-6���T��8��5<,]z� y6�#l'wh�[��cUpͽƞ��U�J5Ӣ�AH�+o
2v���'�DY3o[�cNo�
J�F�gCg�o�؏��w�<�.�ڎZ�9Lv�����⠹!v`��ڈ$�
���)���>aLզ�[K:'�˴7DA"�H!X�Dpn%�A� �]���t_��~��B�#(kM&'72�o�4���TT,Q`�N�(����4�ݥ`E�H,f�G4aF�ʪJiYķ�
'��W�cb2�<!�Tۅ �q�\�q��pz���Ln04K�3��K8q�({+~{�er��+5w"�* C�G�8��Q٠x�_:�u`��o���I@bG��ܲ��/�62����>ߜ��ʛ�f�n{����r��?2��N4����*�!�ۼ����c�a
G��fÝě���+$8�c)�L���,�����ɭ�u�|��g^��-@.�^���5�����]�	#k��ě.G+��^�ܝ�e%����Ϻν�����Y@9�ט	��b��3^�dyw�P$a���m�ͣ]Oe��x�{�Θ��/�]j�����BHvWrJGi-q;']W;a���"��`m������x+,�S���NYQ^Ha�Ԛzm6�-���V6��._��5�n�_��Q&����IyS�9z"�����J;��.K�ܺ�0�����6U�?�%��GDᎹ����ڈ�:=fK�6�=��j��0�����)���C��4 �����p�xZ_�J��U?���g'��O�,��ӊ��?��E�B=H�j1�e��Y��h�+�?����U8�V4'�5o�d��R��u8��r/@����%ͱ��rC+~Y����Oa�����
/�׽2��'�5���)5r=JT�s��ʼ��ዔF�eui:���J���*�v5���D��ʰ�AK�u�*p����7��ȡ��G(�k9��%���D�ꮋ[��@1�M�_&�+���y`'�j8�� 7��@�dG��~�jU.��w�cq+Ө�NΒFʾ0|��������!T�]�'�<�d�B�����i?m�6/p{����˕��͋���m�y��2��pl� �Ğk^�a}����F��׶���t[/��@�DafY������uթ�d�l`S4����-�&�ᗥ���A<7Z�3���z���CV0�g��pYem���y&�X�Y�'Q�{i)f���}�����B+��veݲ�qg��ב)<���Y	D� *,(��ѳ��".�[�~��Iܐ�t��!#��S��f5퓧k��ϊs	� �r�i)��j[�H��H����$��� �^F��)�N.E)�����g I���w���Pv1��"�-�:�A�s!����56"��T	����$�M(�"���_Zɓ!ʨp��oيy	���{y��(ȡ�Rf9��;�_"B��"��|	�K5B��g`��m-�B/>n���L~��Ȼc�0C�Ww�v���`�s��Xs�xΝ��W5d�Q	^�b�ϧ��(�r��(	K��
A`.�@�Ԣ#F�� ��!{�8�- �|�#YNᒗ=$����B0����W;Պb 6��I�O9�uKx�nQ;>�3`��Py�
abT�I
�U�1Ú��W�[8��"�!�I���oؽ��]Bq��U�[T�L�1���2 �;f��,�j�O�����.x����frg�XYw<�:��`#b� �휝�ivڰ�C�\�(��{F#5F��q�����鴟�DzX��K��%�h^�~M�A-�W��{̸��]�P�g8QO"�k�x:�j��A���X�1�3���4L8��Nc�5���#��>3�E��e"������N��S�M���_3�>;�U�-��{��l��UZz[|ú�ቊ%.�Wc E;w������v�������'��G��&U<�0)g���@�g^�/���)V�;����J+���بO���֤��I�p�=��o�mX2�;)Ah�����	t���<�A���$*ˌ�5�F���Rr���]�_\���W��iU"9����Ie'M��N6�0�_���.��9J��C>r�H!��ѱ+��}y5�z�������K�1g����P�:��k�@��`�|���($� �)�X\,g,�,7�҄$	2 ~�|菓��M�Hvz�q.�`�8�so0+E9E�kƵE՚[�k,M��E�uqa�!"�afu��,ᇊ��b	p2�5E��S���jS�=$&��,��_�+M_YD�×A	�d^�H@����"v|��u�?���ZUg�b.�f����ͮ;�}*��!Б�M��)��DG+[q�Ј��K��<�:����4`��җݺ�-�n�lѥ	n�˻/|~`�`�z]����Zo��(��1X�+$��c������3��^�A��H�q�(�Z�)C��u�Ͻ�LP _�dڨ9��|@���y�i��^���-���x۟�����/v$=�m���u����Ep��1��?���C���6�{&� `�J�W �ﷲ2�c��C��&z��R�� ��@j2!��8���I�AM�<��F��eҜ��k�h0���a(�����i癨�Gݤآ�w���"i���?��7ԭ�U�������,���b�X�-ܤ���(��=��xnL���0GE<}���ǫ��ǈ6�v�-�:b3��p�5��M@xC?R?m�ڊ�m��·mI.屏���,����W��q�P
� �V����2����%�Bb0�I����L�p�g�7q�l������aD�b����Hχ2�ٜ�ыV������z�� R  ����x�>y�+�b��L��E���6f��L������&�hG�5Z�����up���K�9���kA��6�g��ľ��}V��X%a$U��A�Y�v_���Y8�"�F9'u��p��M_�{hg�
:�3�Ǥ�W�S��0�3DݓeT�"v�~k�a���|9�z)aa��^=�1/�C��uA��ѹ+���W������J,������Љ��Q��G����aiN��"����cw8U�;��$��GC�`�=��t}��ZA��dP���,��1�B���P'���A����"�Jڞ�Di��LV���ס�3<U�������P�k����cEK�	��W��-��TBw�?_y����Bqj�	MB�EDՅﻝ��#}_#��$)di)��ʃ���G*��'r�^�g��<�ស�A�*��y��,��u.�e��C�f��9xz��'��I�L}0�A9���g�K�[d	�:� �T�g./-CF����9g�� u�0զ��A�G�'�
�j�7~��K��m��*>�oP��Y�ml_\���b�͍�pQ6:~�>%o�(�:OK����'�\�ek8#d(kN�	��$�����Y$�2iw�K�C�Hf;��$�R⢏�^3�"��¬��=�!�>��Q�|*��(� �__�d�H�x���=��I��u.R�Tl�~ɟ���Շm�} 2��cw{�\�9�j�� Q�H�6ˌ����]-8~(�A�����nΞ�'��Y��1���tƥ�S4���ME����`���-�9�Hqܮ����l���%���W������:��v%�W��.�y��+�֖��UP���M\�d��"�Ɣ���^=�l�Z�?i�g�484���Rk�V�C"�� �>��O*3���u�^T�?Oτk���!�Ҏ��x�ڐu�q�>���~��� }���}񬩱
o�I�V)��E��:��]�4�Y�O*G�7���.����kd��`������#�6�4%
�"���_��9h�*5�/���ؚ��?��b���w�&��u�HK9c-ԙ�3y�QX0�����d0�*N�#��T/�F�p��˃���sl��t�G�qˌwz1@P����ʔDc��w&��Z*�ZC����Ds�'l~��O�Ir@��O�6�@Z��
�t���n(���V�b�z+ ��i��5k.���ZVd��,�1N��c��ݑ��`�xF��|t��e��S��X�Ȳ�6�h���-(Z��+��\q`f�.��B�[Q/���^�I�
&6-Qq��m��8H.���k�5�,��)ˍO�'2d��W�	��0��~"��[�;"�@H�@�%�SY!�_UqH=��/艸�&�#�M��#�~�A-GH��8�sq>�E	,������'�^��	o��:�-07ٵ}�����'|���"*�]�]!q��+h,c��RG�p�͚<7.�i��";V�ĸ�3�:��N��j���>��(� �����}�ܝʶ��f^�t���fчU�߬���f,*�T>�M�)ϣ��IF?j�F�Nw<t;j���i���YW���٢�����ٻ�	r�eÒ!��[gt�cS"�YN��k�"KʷP�
尃�����ym"^��{��R7ɨ�L+Lj���9"�TM�.3��ja���@��H�Y�饃HT�#(�G�4�2�E�ll��	�յ�&LvWk��M���&��&����s?3��FN�lY�b��X��3g%Q�U%> �w'���:֏ZJ�������{�sb[�}b�Dm��I?e��۔�F��77����diT=��o�5!�*3�&�&/!�On��4��<��d�:��]����O��p���.��$͌�ݱ�!|!���5��Nb�CC�!�ˀ�2��;�A���KZY��>=Lj�e��5�'F��yf��.�,c+FU:�i�{�a�� 6
Ի`�+���"�4�񼡰�6����Ғo�זs�k�����#���4Z�1�%/<���V��vכ
��${��/�۟|I� ��Ye�NcG����iZ�?���I����&ʈ�[C}ݕ"�Y�	�3�>�xI7������ϱ;��)Z~�1���J~�4�۽�J��ճE9���=��7�����x���A﫼P�9YF0C�YH�=��P\r�	�>�n�%��ߓW���{��z�	j��Ȫ�8�\j�����Y�_�Yk�z>7�}�Yb�b}��cm��gȯ*����-����^U���ڨ�=l�E�򓷪~j��oJ�r��Y���vFy�л�ڔ�g� �b�恹7y�e�>J������E~�Τ�Pi� ���/�d{���ǂ�֐�u�T��_�O��t_��������ު����J��m��� ���K������a�*y�hf�qR�aa��ND1�ֱ|ǱL�Wt�9�VS���3�ʣ�]�Ԫ��-:�(�4gJ��D�K�h�_��3S�t�hN=.���r�;(�'���Ӫ�Yv ���T�^�.�I~|ҼҸQ3<d�di��x'�c8ND�o[��RL~�������`��o�r*v���Ͳ�:Fa� �B�}c"�d�͔to��{��4.�>9��lWHS]ǩ�
:�����JP1�����~s�����5�E�A4��܌�UOo�Y�)�]��w_�k"����RҺF�����>WxD�`����lb������u�,W��4%p��H-{�E<ՆL�STG�0�,D��wu��Ν�&��0u���n��`*+>%��T��W�ly�:����	�a����Xh>����i�쫍y����ڤ+":�/0>|�A��y�4q��SI�Q���>�W�M�E�@A��<L�3�K(4��ײ>#ltHԸ������ɲ�N5oO`9J��}�������ڵ 9�A�ʙ��~e�wr��`�!N�m���b@�$6�s��/�h�t^H� �cY#$HTm A������H�e�q��ƨF�f��c+���]�2�����/�{�׮�1���͘}Q⟥u�j�����c���/�ZÏ��E�w���N5��?w9Bh���큢���S��3Oש)?6�br[���?�6^iլ���S�)4fǯ�ܺ�����sKy��ҍ��G�����͒A?Rǥ0� �}'UcXC,]U�����ݦ�W �XdQ�f1�P�1�Y�O��]�e�ב�o>7XA�b���+�E^��W/��cT�P�h)t�>�VP����i`o��%o��Ds�A�+p���o�ȇ��	�/^�~JRh�i�ܢ���Wߠ2@�ÿ�˕�£rnz�@1&Sb�J�*�3�&���a��D���Y����m��Z���#1����罱|������x�O�}(�I`������jB�9��,���l�uZŹ�J����#®~��1�װj�9z���v�[<�p�M_��Y���Ĩ���[	��[�<ٱ�"�C��M�sK�G�W��tˡG����q�,���ƀSЁ>��II�RXmVu�k?H��-dY]d�ܿ����Q�z��SJ�eL�)�a+��3�:��$��i(Yڸ���*��9��r x]��s��&	_.��W1�
e.��3W'c�	����f8�Oc|*}�����čL�����
��7��-QX[T���J����[:�qW%M��=w�JUA~�[����{μ�4��g��m��	��,�Z������!�7_���tR�f�!�{�c����)u�Tq�hWha69oY�K$Cz�l���s>���z��I=�� �1�Gկ�mEiV1�H�Ɵ�噱��u�v1�S�c[�!��(m܌\�>#�fB��G~a�e�x�i/{��ۀ�A3(�B2��ձEm�:��s��	��6\`x�߉�?RjMd%�|��.�zg��S�:�T�����}��U�=>��&�ݕ]��m�uk6w�T��$+�'��$���wf_��P%���@b*�����m,$�ʢ3u~�JR��o��Db�ڜ�71�z-}�I8��J���~� �VE�J�9�󤒩$ȑ����oa?�~mHyPv�L݇��fO�o��Ң�������W�7Q~���k��k@�Z��'�њ�	h����ON�-��SN����z�.tO"�5�s܋.�eq�����D��AhE�ܹ�)�j%_�`��-�ns�}̡ߘ4@�N�e@���q@Nt
7�d?���O���
��H�2t;��Y|2����tT�F�?�����5��=0����{�KLi�e��{[�3��xr�q��g.Hq ���������F���F$�))<PQό�����q&�T�}��["�P\�{���\0)S�b�.O5-#p?D���:������Q�4`s��w��6|W���Y��1���<�H���m�3U%5��h)e
r,xB�����q�JA�M�(@�iEi���':Ϥ\�n�N$����2B"����V��|��Z�^)��&�fv"}S�Ǥ���1o�B/��A�*wS��p�}ِ?u% �Į��;J�kW�m�����-�f;5|쨛l��"f��g���2@����s�L���
ymYW�8�y�Y��h�g����!w�>NVӷ�2�R�����!��W�p{4CN#��cGzI4�'4�Nj�����3�A��@sy1��n)Eԓ'"��b{�gUt�=�5~>��D����,��x�9�)���% ��iqy����+^������X]G�N�������OF���7�sBw�F�m"(�WX;�C@_T�f2?��YY�*��@�).�XZjs�ɓu�h�gA�����hyN�p��F(�`U��������۽w6�b �3X+��\�x��quFQ�����8a��d$�������Dj�Tlߕ�y<����?D�F��'��������ʇ4�i>��T\���������_�2F��j����ǅ�Z $$o�G�D��B9ken�aD��~���^cX dR��?������c{\k��=a��'�X��ÄgES�4i�����fc.������ێ� M�XqFs923B ��N�_���H�55-���h͞�sM4s����@����Tņ'0�E�3�ͦ�^_8�M�^���GҐ����V�9+�y>��h2�[ĥ�|צ� tv�q"�<MM�%��cP�����C4��EMBE&���J�6��@�5U�>��K~��%�i�*Vj��`+uk�R����>f�H�b;��6��JG|ֲ��@W���*\��t��5�����y+i��^0/O���8�r�^�?&iVQ����R��o��"�0v������7$V�S~O��8�t%����k�5ً������1�&��|���L4�ƫ>)k[���Q�g"�m��btO]��k�B��:�Z�hΐ���X����lf�g?>�^׸�4/ኅ:q���¡5ML�ۛ�\�-��1�cY�   px��
&/A���z����FB�g��hYxR���9DK?+~�d0�5�n���V���p�d�Q
�O6���^�-̫ �a3��{L��*C���F|�`�M`=����+�|�r;�ѧȅ{�����
��T��iaW�:����CŴ�n��e"�il���aެb4�J��C��!{Q�.xĈ,�:��,����7�0�z�lå*���eU!���!<e@g���(q�&��%WzQG���V�����z���i�.�ƹ���{�B�n��7���X���G�A	�D ��H��,��mԏ7|qO*%�^xQ�<�-c�8�k�y�z����[士i���y|N��?��1!uQ���>mK�Yճ�e�� TL�]!�m}���2ݩ-i��C�s�1��ao1������!������^[�Hu��G��.���8��y_R���&_9|� Ia���K֬���d���ТP?z~o��A���>�yOhs8��<���4c���Z(��F4.O�ؠ���lp,��BA�q"�c
���25��iy�{a出�JJ�g�̌Gh��8�s�q?���(�{.L�s���[W�W���.�den��he.'z�Ԇ�9~�� �!�)���'�/�,v����[��(3ðL��8�p��� �'j���k�&Գ/���K�AN�/B�lϪԁ�a���t�f�k	��-������6��'ý*v'ȋf�B��aѹ�ǥV�.��<m^�pt"'�����&�zP._s(�u���{����̙j-�*Il�şcf���Ϧ�b,^�@-F�)�7!W8�`�����^��R'Yj��� �,��{��!�f�8qA��oG<�?ie�ԚslB����?�RQ�\���b#4�NQ{-�AJ�sC�0oO���΂>8�-�����KῙ�أ�֔ ��v�
�<q
{�o�->{`�w�.��f�=�t�{V���ͨ�/i:}�� 	���ԏS��=5�"��D��`���{$�ag�>�Z;��Of���" k�6
��J7�ucM�f��{���]g�+�K�������:g�2H��!�t��R{cQ��mZ�ā�:�<�`��W��uݎ`˃�(	�B�L�\��ϐ���ꩧ}A�x�TMGό/�0aku������R������^�~�}����H�r�O� ����fmU�`(��F���J3b���R\��7�Ʉ2uv����.��GN��U���xXG��$@�1k���3�d�_�K>�(��N�'�[5�
�|������z�u�e4,�
X�'�p6`�c�@�mn9�.��X5���ނK�q9#nKwma#����%��go�Jл�4u��q��H�����i�b{\?@�)�����SC�p�5�q	(՛o�����ǁ�����]�y�D`�;xhQ�\�ً�c5f2b�YZn�Av��1�,�˨H������@�y1���zb����ڰz�peE�L-䲗�8�ӠO��V4,���$z|v[��N�A��\/8R�L�	s�}^?��ƅ� ��X^�����g?�P�\���>y�>�}Rg��N�pz�_�j�UY�Bߕ�W�i����ߞ"�ED����b���-}��vj���NyכZ��v���ʛ���wE�SU`�Q\�:槜��w���}7~�y�Ckt!S�sj�k�$ p�S���f~��po����:<f��`�0��%�o�Jqjb[AZ�̙��ԫ�­q�9���!x�R�O*�G���RS�����~���eߎ��d���YMm���8�0��z��[?��^/�ƀ��^z�w)�t�a�S� $���չۭÖ�4G��
}8��f3'tG֓B���8�AcI��(c��N8�/�vg���[�L�,�k�B��8��O��xK�c�|�ѹ���,�b��u(��f���P���hK?'o)��,D8t��}��WY�T����N�/��ǊP��q���3y���h�0g�WN�O}��%D�N�@QC$�u���ˍq���O����2 _H{���<D�H�Vn���S�-$K�u�RT"0}� ~�r�m�쌒N~���ڃ]C�4$���X�l�
�q�P	M؀^;[ ͅ\�Y
qsJ;.-I0{�����0�����ÊWZ4,�Պ����f Q֡S鬷)�F�%z1xu���G��I���5�8��f��c@&�n3�Ġcx��V� 2�K>�e�TR-��,���(~����j�`EP�@G뽄&�oۖ�ܷ|W��?P��;9�"�ȃ�G�^��jZ/�*y�q�(�/���V��w�aM:����
8� �
���9&��^��B;b��Ŀq\d��}ph�*�%I��3;�wi1��]]K*+#Z�d�d�����4@��%��l��ꢵ��%D��Tm0#?�7�n͸�!Ѣsd�̐��H(_��������e�]�xS�}���������Nbo]�s��M���W53�j���J��Eۇ�Ad��`P��_���ў 
�^�D(�;�hZ�f��OK��E����:����Ǚ}10�W_	(��eqP�����o����qʆ#s��CI�c���+����
)�7�qn.K\s���͡9�<��NHt��Ɣ��eP3z��r��q�s���d0J�f�ݰ{���*H �������D��j^�I?�G*�?^�O�E�L�A;{4��AG�/�+&�rw�@.�gel�%0H��0�r��O�>�x�V�އ����fD�|A���I��E��6lI�'��A���P�Ý�����+K���g�K;�l��� �dx� #���ӕU:���yD��2N�{B?kF���&D�յ��6�o�`�0��_"8d���N�����6����R���<r8���Dsk���YV�J��O'��hUl���U3���#yNv�q�Ui�T�`�V!3<J5��
)��03�2�R���Yf�yU��_�i!��
���8%�Y�T����RL�h��Y��n��U|��ޞ'�U�-@_��C���N����U5}��sJ���_��x����
;`-~<��&�g� ��=�}��V��5����+�>��!�Sr�,1 
g4��X��-�1L���V��/���&�L2�ԪA�8զ�>y3��证�0�Eѵ�_���=��Ј�n�8��}�!Z�u�S��Ye�F�,�aO��?�h���N:*��o�?*cѽD8&��}��T Jh���6����@]�H��&+RȌV��!�?b+(����5q�!v�ҜBv�0��;����~m:q��c�԰�C/9�_�-Z�{�J�Cv�A9�����&�_��e�j�G;��H�!�1��q&KVI_�L<`DW�z�gm޵�d_w�5�b��3��G`���ŃB�k���CL�;)ޏ��W�:ٰ����N�cm�_�X%��;�_��,�?�=�
�{�w�dn�,%���c��{yR퍷�[��&Z|I�
w �/^rg�I2�i��x�>@�&�2��?������b��C7��S���DB�Tf:�{E�Ka��}ێN�u��vB�NvEf���26�=4+���J���g�h�ڋ{��.1�})�M�,?"��2�k ~�U� ^��ڧ,L5s��IA�(|�T�EZ7��L�k�?�á⢨`���	������t�5�		� ��ɻ�|����Aˏb0?����&��￈�7Rv��S��.����MP�wX��z�BEJ%y�(�~�o�JJ�Gr���+�Z��&гs��r4Ɨ�ٮb�F&"?�M18'�QG�{:dXLq?K����ME(��4x�o��6\*�YF�_F���B=�V��e�Z����*��F��!0���Wo�c�)AoC<M^��T4�eM��9���D�2&΃J�]���4	^�RCRV��R�P����M,H�̣�j;�d���	CFJO���	�^�7��\���5 ��6�3�M��FJ�_�W�3��ҿ)W��Y����L�����u�f��a �r��W��t�C9�h� &N�����%�^����-6��pĢE�#���΅7�﨨\�DW���PU�W��1,���ک��I���^C���42������P��*~\��8�6O�5�����ㅧ>�	E����	�)Ȯ��:߻8!.�WE�t����D�L����d�)`�zu���;���8���A�H(h�4�#��E�^�;�8:��d�9��>�jM����|��N.ӹt�;��(�[Tk�j솿�3���=���d����lE*�ܰl{,!�����*�d�`�ȰdF�<��t�׌�2g4�<[���|W�� �A��9����X(y5%{eA���փ�Rq3#?6�wY�P;�ꁝ����t:�$�#bk����pc5?l�}\y�Űs������*���%�î��̵BX�����Ji*�7����x@�ah$����p�*����ZB��kDV�[���WQ�=Ex�������:�dQ������1l��J*�P���TsV����7�)Go9R�v��(�^B�ܩ>�/�"�m�DWj�Wɼ�\i���L�����2�AK܇{n�ʘ�/)0}�]�����Y����f���x��4җ��t��2�t�f��͗
;[�0�b �B<T��H����0ȣC��]ET�S����S�}l�/ �����m]/�I1Ѐ&��Œoj#��^w�ː8�ZY����۲���H\5�"�"���f���4�f�j�� ���˶��m�V����i����i�^�Q5`�)x}ak��۪�s4�g0���O0�\`N�G]�;�~��wy��xl��d{b�P��ԧ���ͬ������y���p�Ptn� ��%B������c�J��SK0B}��i2�bD<S"��ѩv<~���W������\�����>~���D_�Y�F;����A�@��J�>.��F+$g)�����)�߬w�I%$0�����{�2>�1�QnD�}��@$H���~�*4�EhR���� �E���Ҝ�h\�"O����T���ן�np˝�-׎����S!���%\�2�+����� ���C����e�@��%��-Bg�@��?���$0��7C����IS�"g��u�rV7���
���¿,$?l ����m9��G܌�ep��ٮY\�T@`['�p�R����٢nn,�}T�y Ð6֘�Ր+�����QˁQ���h5�T[M�������O8�����S]�.2�LQ�@�!��8x�d���ۭT@rM����Q���������t����/��m�hZ�3�����}�q�y�o�.Y�Q�(E���i�ԥM��-�k��K�A��&��E��D�'����l��G�)�l��pԃ3�G,����X�Ku�.+����+������+������Pm,�Y�"�W�KS�lq���<������<���tg�VYNM|}qD\��uBV�m�kd���,k���SOc����n����lZ�?vB��=���ˤ����z�)�,�W�qXw�+�9u�E���d�P���VEa�d�i����}~h�x��9���{����!��t���=1����Ӥ�Ӊ܏4�0Դ�?^��'H;)�9�w̖�9z�O�_p�<��r���{���Pu�#!(~f���(&a��w��iP V�E��.�-���}Ұz��lr�cW8r���Q�[��l�4+�;�J������ѵ�/a?}l	��r��yPA���@6�g4���x�Ξ�v��Q������
|�J5=L��(���u%c{a��ˬV���y}�ix��Ҽ�ȓ��Lo۵}{�Yd�I���3�t <�1�;F�jW����1U|�m�9�<�����Z"�̕�}Ld֠��G�{6߲O�'��;�a�<����]��l���H*���. _U��7c0�s_��ce�;3' j+8��N�7_����DoJ��==������ξ[-�[%K_��U���h���尻z�n/��t��K�#���s�ㆭs�����V²,v 4�U6ނ�e�8��ㇴ_�_���
�2դ_���\g�'/N��:Y�2����T�k�ۛ���r��������8?Q��������!�}`���.E�'UTk�oW��+��#�wܐ����1A��ۀ �?'g;k���vv.#��������>ƺ[�$h�Q�����G~�����#��dZ��I6BS&�	�hRS� ��q�u�y	>����[	r�|,��j9��$q?�H�hC��E����-�\m�C$��ʘ��9�[�U�..��
��3���Dpg+lx-���;��32��)�}vf�O�]{Pf�9uaq�ah k>a0
�m�y^�h�rr��3M������eP(�+����ybĈb=���b�/x  ��bp,qfJ���H��Ln=�b��O"\��YCl���'���++Iۅ��I/G���m�l��J'C&���(�TAU��h��m��5�N�T��k�EF�-G,����� Ǽwp,��M�"P��0��Օ�l>��7�Y���7~��֑���Q�E3�A'�����K�i����u���D�;y�?9XO��eO'��X�
��U�m�.���jp,I�Zp���"���Kki6�P�;�R9+�3�8�MFѤ��N�ȏݑ��D��W���a��i����_��镁���4��yJ~�)2�ܷ�U&7C���P|�j$���-���Lb����G��2M���~	���Sr�A�}n��u�B��y@h-4U�Y��	�Tg�\���Zu�S��f�X��G;��-1�Ҭ*����N��,vC��T� d�ol�#� �3�#�/jg41�m�!�2��׻�3����><��|Xn�v�,p'�Ϛ�KN �m�q�C!�z7�,���Լ�qU�D�].�_��Z���!q���""_�K]�����2�����5	jq�D�o�8�A'F..%G7����y���RzF 
�����n�7�t^9�����������ͪ�5�ҵ��,g���)��=�"+�Z����v��.�u��`{j�A(�?P��T"oUv$xo����)u�_���i�T�4�\A�θ༆�,�8��k+dh��LBi�X�h��nd�t�½t[�\��YEs���I`[X �{��g\����<-��x�~���l�?�s6�*��|��5���y`����w��h��V�sd�!T�d �'%j	=M��Y�l	�ćV����k���Ù�6`��ȸߗ����n���P~��Y�ukr)Y
�,K�����2�hh�྅�k�.�k�oFD�j�_�cie+�\���Ƭ3e616�[mOvs�HF��������O� Z�J�y�e��L�����&�֪�մ��"�v�W����V8�	T���:r��Aj�^)�G��r�ǣ��d���N]�P��6���ڡ��v�����8���2;tJqK+Y�1��<���?7�&<��0YB�S�i8[o��や�p�CC����-�Jx���Yu��pr�I�o�qF�bYdZ�}�!Me�n?#��3K�z�bd���X���9�G��z��	��&��{]������!M�9#�7n�	l�+q�~q�SW�9����\CJ6�^�hE�����2�﾿��W��[�=�N�[.��Y�U�{*�{Z�߉(<�%M#����-3�]Ս���@E,;-�5�5BsfH/�ꜧ��-�Ai���܄���9��'m��p7�t5ccJE�2�b�y޳��p�8��*����k��_�R��J����M"����l,���gBt��'���~���}ūO�=�! Wɫ��E3R�m2�X�"�
���>��`�9PݠK�]�r�`��ː��Q�s'4%�NYݙ�T��������[�g�u���nN^�p�J����rs��c�P�=���Z忻xiP�<�^[h5|�)�1�����SE�����"f�K��HI�[&�"�}�j�[��&�y�����4/��]�J����Ǣ��Ԭ�(�V�!��Ͽ<�2�w���9WG�	��8.PV�D@����V�=_{���u�s����"�!O�9m�t5J�kݧ�]����G%�~�{B2�I&����vΒ}�����%�x���#i��L���qZpw��	l���I�$�L��� P�q���zG��y�Qc#��ӥ�g���\�}3��vPSwu�m��L�ɇD>]���҈T��"�T_�Y8����짹����3�����a\�'x?,�����*"�+�-�J�EM�᱔�ǭ����U���<z�1�J7eGը�j��L�[��N�/i/@QJ3_����kB��]�e
�Җ��)���g��R�)y9W!����Ͳ"f��jF�n�pV.6�H7��e�
#C��Sm���UL�LJ:�p">Z���}O$� 3�|��K]��ڗF�?��x�#w�	Bt���B��_��C�l�6:�O�x3�,1�|١}�=�Ijh�*j�\Z|-�����u��"Qv������Ԑw�؅!p�[}��<��g^ѡ�3Կ ���b����8kW��P+�������'1�1�!��W��E[%v(s)���d#+�}���U�����p�|�5����%K��w�Fx�^�����W�s�_Y��yRG��I�X��_�B�T��%�I���:SPg�[�
v�u@Z,v�V�ot��ky^����\��!6k�F��o���l[2�<�-�7�iBT��q"	�PA��(�|��Jf=�.�b��%���?Tz:�\������}m	�/�8_x�F�� �W"�'�r���k#�A����
�c�*輒-���&+�q��2�Q*����=�Hm��9�{�C}�(1�0l`�T�x��rܔ�0���e� o��Q�x��]sXkadpQ��G\Y�9O1<��6Ώ��SÍ�(��U�R���E�+��<�!�k}U�9�G6��`�d��0�>����"�m����T�D���P��p>)��S�� ��~�BF�т-�o�L^�hJ�M|�N���@�k;�w��T�?d a�(�����/��t:\�S�ϵT�;�Y�����D�p⮷�|������<ϞD^d���0JZx/1'�
˪�	�*��^,�l���� ����Xy��5����VE�~ٌ=`�T��ax�a�x2�π�%��"ă�!e����#�;�Yv��z�X!�ܕԴ�woj3�Rc��	�$��,U,��%{�O'�}E 7i�Ԗ�Jʟb�*,��{�_K>ln�#X��R�a��󹌑_b Toy�G@�ƈ8�|{J@<ߌ'̒!c/K�f�5n�+��:�8{e�c�7+��'���%��]�]����eH��$V�l���el*�T�����aRdD������L�� ��@a��/�c�n#��"6b_;�`�f*�b�u�q�L�^?�z5�',	����AZoo?��$����(@��>���q�sde4��ux�U��*G��;A�̥V��7��Sfe�������܁Ol�xgWY.��Zw��d�cL
}nrs	��E��?_��=*�g	y�>���z|�W��'*�\�x�K�_���o�{�#i��(0���{��qB��sF��T�8�U"N�H��D�C�����{�3!��A��^!Z�o�y�q[�u9��|N*`�C"+�%o
����p�ξj!�,}V�U���9�A����N&u�V��R��ntW=K%,&��P�P����$U��IIxF� ��ͨ��~d�>��&|�쓤�#@��\1+�p���?�s�_����o�n���������{~;�pr`�ӠUZT���C2ٖ��\4!]=��ׄ=����
t�R\�4�n���� � 1;&�4�Ï3_zY�;�9%�3;��ц��-?"�5f����g̅ߢf��f���*��$P�{�n$�CȷI�b)�NG��s��$��vd@�n����2���������[첝7�Ma�=��n5���/�g�.�fR��j��4�(�3���_�"LG�� 4��ɿNxbXptJAK6���0��br����U�I���-�Q^�⌻h��7���];���^�� 0����2�5'�r��À���`��^�v�]ōzb���e}��ep7�SL�hѮ�#��Gn�e��ѣ��U���f4��R!۟kus�~�ƃ;q�|�]+�ld�Sdz�ƣ��40�E�؄�j�$��b24���@2�R?��%�M�.u2�`�̓�R��O]G���"���Gɞ�T�,;�g����I�>B	�)������ �A�ޞ��20���W�F;VB)P XZ	��t�w�aA����h��~~`,�T=��؍Ǩ͝�/�D0s���]vB��1Y���6
�]�����76b������!k��YF�Q���'�Z����"��.����98�̓*��.�uc�-�&�o���|��c㢄4�ཫ�o-\}5�Wh땠3� �@}s�v	Ҡ ��}�T87;Ϭ�$�n��m8�ם��</�⥩P���Kga7�ݤ}Y��˄>��H˦(s��bY�T�b����\*AM��I��ul܌����6��Q\�R�$��6�?C��A`J��Q�/dR�N�{�=��%�)��4M.���s ��)��'S{��M.o� �ن�~�h��o	�k��<�ӥ���D���Enf<{�z���G�X��v!�=:Е�Zl�4d��]o�-T�d�� T��j�6���Fo��v��4��3�[c��H�=��1$�K�J>Rm����+P��E�H�����=�3�?s��o�@w�Bx��a�NV��*)W
\��Due@
��%���v�Pm7d�u���}_A���+�BF����Y�Q��Q�Z��� �fi;�)�gաQo�I��ws��*������D(��̫$8)%�?�vyC��z++4=Np��4e����sʵ�ܘ���YKSzQQ1+�v5���	�r�� 3}��qNU�\��)f���l����Z�J�������P�����Z�Ԗl�)����oO�@_@;��y�iS���i�nrr�����v�� Y�E��$�A�[��u�ڕ&u.<(�"���A����*�������?�	�/�r$�
Ֆ�[�N /�}�� ����嬦�`2W�hD����"�j���H�WB�g��G��tn�BU��� ]Pj��\�M��������j�0�"B���(�ˀ3���_<E���q���T�	�l�,rQ�LJ�$)p��wpS���l��;�G�k[Z��>�'m��FX��������֓bK�
�\�D{n8�A7G>o�"��7](�۞ϙ$�:�J���@ʪ9v�Ms/���8�)���D�)�p�C���}�m1N�;���s'����W2TF�8�z�`�a+�6a�2���吪��+}<���枕q�R�!��u�_�<�t�`ً[y姟IP��6���%��߬X�Bk}!��ȸ�j���<=X�5��+��t�j.���V�ѨI	���n޳X���j������k���ztL:� h5��=�Y�C�Gаv�R����h�����G\�vn�s��)TpxJX��f��.�*�l�M�7zG�{��jgJz�P�Ӆ� U���cZ���!��r̠:��8����1h�z�ܰ��5���p<�,�;�¤9��bM�H!�J�*O�C���t��E��Կ�DӮ����UP���9'��X"Q�a)e2M֡ ��� ��h�#�)� ���$+V:� ��l�S�8�ADO�ݚO���
�U����Fu�w=�x���+���N���(&4=h�-����E�&Vl��x��$����Hd
BR�GK�j-}�ؚ��&�����E�5!��3�)��Ȓ?mu�x3m�ㅂ�F���9�ϐ�M6�h����v�����K��V���b6����bUr��@� ������ C��FPh�x���d�Mr��Cb�Y�~�B��]��<�1�`�fc��g��ъ���L����bq����g�4����(�~�rM��>�J���wB�rB��V����R�ʿ�����N`B9T&~;�f��B:������L�} ��s�]�E���bY��U�nJ�^4�� `h�8`.ns癗��i��o��M̥�ը6� /��$��՛��Z����.kd�&��I�Áub9҇j��*_fg�;jE�d�*R"y L+O����2S�uu���ݐ8��?�r^�\v�)��<yճ�bU>���deo�I,,������������TP6[�v�~�#�8v���S��^<�EN]�O$��9?̏�c暈��b��|*A����1�y6I �U6��]�v�H$��3���T�[{����piu_7yj�ү���"���T�{:���b�N�k�{=ˎ�a�����hdO$eZ��!c�.!Eu�y�G"�g�eSqڌ'|��+�=f~�jAe$ u�5|��x��]()g!m�K�u�5����x�������iDi��K��8��y?PQOC���!��}RJ��Zō���Z�!����K�T��L[cV;99�S: �3А�pR�AZL}�\�b��/��a��9�\��u��ꌪ�cb�]c����g'�ͭ0v���s�ؔB�$RY�dYE�g�W�kh�s�H���է]�؁�|�O�N�m�8�bjx��tm|��N|CO$�$�Lʤ�a�BZ�
�Ij�2{z��cE<H-��V}8����׎��A�\/ֲgU|~�ֳ���|LP���{x��٪X��+ �~� � ��E��-2Q�Ou
=�Z����*��gU�X��4~Zaa�)�B��L2���!�^VP;�3� W3ϙ�t��ѳ���?����?q�jH��}SVs��T�O,���7��m�X�Li|.`��Y6�t)5>���.��5��Q��~J��1��2�(�5A����7Ig�A=
��r�)uP'��p#l2c����/��Q%�x�-߶|C���ﺋmL^�6lF��GG�`��.��1 c�������Kq����(p;CB.�̤�xN1�,���	�sV��`d�X�=�լ�:j�&5wd=���usKL�q%@�����%�� �E�J'�����"i.1֒��o����������P��j��E�ZfKF2=�hɢ����.(Jf+�RN��?g�Fct4�Y�G#ay��"�ܑ��~����hs�g����	Fv�/����20���p�U���Jbr�_��H�b�{��G��P�j�;�e�^��^}?�͌K>d�?�]фv"�R^��`q�����A�/�u��Z�'�^�E-	=v:�dI��MD���k��!e�����u��K�t�/��+wF��6���4������q�SH�)z�?.l�Ia3�^t��9���;�#���DЪ�n��S���������K���l`ңHH��$��
G�����,��؅y����Ϝ��ˋ��T*��yҋݠ<X!��h����Ⱥ!���(�ƲǫUȄ����I�YW�!�����Cq���-Y�[s�laC?#������@r�y���d!�6�v�m��]"�n���� 2������i�&:�D
���:+j ��\���2Ҵ'@s�zH��^M^�OO`H7�Ӕ���Ƙ�Cۏ�:�(#=�ea��>tXPDքP@���u?]���!
���.�a��a��z0��j�Q��^`m��:x�ϊ��t���A�C��zb�'�Ȅċ��e\Oֿm\;O�/f@�C,yo����j���*��o��" f�Сn 2�b���� s�gQ��o�"��+*��=��y[��H�_H���cE��9��E>����Ђ��Cx�pH
W��ݮ���}�v'1�Vh{.x�� �<�|E�}���}��FK��/)�6ZpnU+�H�������!fRq�?A}���B	.��+4�:�S�fѻ
�أ��.�2V:��{	Y���=�z!l]�Cϔ~�Y��Ca��q�bM� 2�F5�xV�o�ͭ�~VirxI�6[��z�&���)[77�/�q��h����:����lŧ���' �r��TU��$�=���FPk��B1����DՑX�WǞ��~4X�I��S��:�u��y䤲;����t�^�?���7a b3�]ٰ[�͸$6����2�G��}6ѨTLR�-��%5��Zi�H�rN���}S�u�a�t#�mϻZ����p�j޹�R9+�#s�u(���E !,wC7�L�^uԵ��b;����\�ԑ�8��Tˈk8��>�ɢt��ɷ��M�IW�Fr�W+��K�ϩEۙ�������
PS�ė?9���7����C������7q��a�9�C!�x&��|�N&m���2��u�b}���W*�y�Z�<�zD����G~��?,$����߀t��R�,��Y�v����E� �bC>�7/��ݮ�͔`�d/�?�� K)�����迓}��5.���#,�g�����!ָm���r��K^%�=vR���g�BR��Y`��T	����f�T�wciL��W�\N7UPl�����e�T)�.p?<Scl��>�%K��&��Y������1�F��\��[��PǍ��B�"
8���6�x�P�,����dF�����3�q���W���.� ��}=;���:P*ޯ�	� �� r����植��ѭ�
ކ�箛�Fkq���	-m�f�����F��[�"���)��r��}�x�W�htO���{A����>\���2v-XS�D���air�vT����a�􋋺����i^���� +�*�q�-}&�j������P�PBݸ�n8��6�~��5�	T�vK��Cx	N�C�6n{D�֓]���^ΌY���U��d��{ �a��h��IS���:�b�.���D�xt�<"�*.��x[��!�[����'���d|�Aaw�y��,.-<��Fs�R�>A�g�П����ɺgu�A� �\�2�/�;��xrO��E��|:�f�p����D����/�=�1��)����`^po��˳' ��������
�N���\u�{窶˛�*yP���<7�EZK��2�@k����bMJ�`��x����"N}��7�Q]��H+?�7C���0�-���H�����_�It�,��D5Oj�7V�8���1%Ck�J/��S���'����o�2���I��M���/
~M�A�ra�<*��9'�i�z:���z	�4�C���C�Lxh�vB4�� [��
�H���	��+#+��}=���c�<��Z&h�O��0ۢ�U�x>C��d��o�������e�P�ʣk9���h���qD8��)���+��M�zY��*^��z4��lY-���Z!(dFhD�RC%&���3F�d�� o����m�;�c�%�G���jv2�#��,DfK�}��;H��4-��6m���iN��#��R��q������њ�YKR��M�	u4T#��Yl] "��4�k�p��ص�(*v?�CߚL��oY;9'�[G�{�W�51 +����W�p��G��oo29�:\m|s��eecm��؁c0�i'� �5�8���n<_�
2���R,1�8���_�Z���������ɖ���K	W�P逻�%į���x^
�@D:�����b�(➫�U����s��a�[~Zwg���F[W�+ဨz4�w4��3�JH��56M�	F\#%'����Z�Xo[6ko��,��̾\t��ÍG��4����A	�tF�����ɘAA�U#�\F<�#ln����&�؊Î��(�%�Iy��R�c��H�6�F&�70m׆�/���Y���κJ��cP��.ܿ�f	jv�S��F۶c�ѩ���J�0o,� i|R3;���X`_yf
w��}��
>��0~[���Yɪ��������$��&��2�������Z�����1kR���Pϗ�t�i�J�q|�{��̈/f��Da�ߝ�֮�����E�ݟ:������VӖ��bpȐ�$���_[���'u�ؙ/����yc�1�)΁����������5r��c�@,����#�-����݅H{�8&"~Õ)�j� �&�f�f0$��"�H�rE��ٸn���=���s,����`l�!��cf[������ȓ���|����X+�yG`C�����| ���zH�ڮ;͹M�<��ᄹE8m!�7��}g�|��z&�O\����[M,�59,��7`��}}s� �U[:����M�F1Mi�����5��P��)�(])
š�4۬����7�1T�����߼�m(U����HŐ��[�I��00B�f�ҩt�k:���8|f?Hr���a��9H��>�w�"����$J�J¯8:@���+�FG�o�"�Iܜ��IM,D��l�k���ک��v���\��c/�vF��u�\��������9�/N��q�VL	ͽ����S�r*w�o�|�Ziז�j=�⪔s:�Ƥ!�����I�T�W���t�"d����
��ގ��#4��Ⱦ~��xi�u�����>����[�9"Y58W>�k�Zo� u���-�KME��D̠[�H��s�毧L=��d/N�
ѥ߹
�� (��a�N�h��`�X�&�#�\&wc���>�3�{[^�M~�rC�?� ��ɑWGO�.G�M��C+�4��:�.�V�������|a��t��&d}c��c��Z�}��(uh���y�O�F�Z��l���ɦ��@R֒i�6Y[M�Ӡ�cr�b�W����pj&���.��o�:�y1��gV���cBi���9-6"Z���\��Q�hlS��%u��-o��5�8+���z�E`0������f��Q�ð*T��B�g�2�-%���w�i�����A8۰ۗ���n$0��rCx7�EC+�Ӓ�V\Xy��hl�W��H-u'�����9�R��}H�e>�u])�v��P.�(#b:��5Y5�ɭ�{�B��?3�X�n=�v:u�S&�i�Tvs9��껤�i��=Ȫ��ظ}��^*�Y��W4�-�2�:��g
��Z��tT��As,���j[����Vv{:����j�����j=?`�Zu�%1:%�כ���;kzg�үX`�R�[��E#2���Pſ�����a��`���&@	��oA;O�Y^�!�8��J�h[��ME�`�u��2�z���+P�J�ޛ)��@ �("A�j�,
�_%���xF��b��9|�� �(��"���}��^��t���	�qJ"��+����D�	�ؓ�L#�g:F�%H7F���}}�?p��*��Jyi����5��ϻ]3�3�8�ch��y \uh;xq;�lYK�5n��I`?�xiVO�H�D`�| ���-5��	�'E��LF�N��v?��ݖ�=�
��=�7�:�>д��Tl�>o�e�C`�w>%�Li���m���+���AI��y:gC�0A*�۵�*���=\��o4 (`g��"�j��pΧ��	�Jt��sM"���M��!3vΝ�M�̰-)&���w���l�� ?�}��^��XV[�BbSӱ�/�Y�H7c��ݧ��-[_�WQ�dңO))-��i���'��v�-�A�2�12� d;��t�陋G�D�#\�;�C�C�!~0[b����	n+=_���`���Q�Ƿd_<���¬nv- ����T��nU��W0��z�yĈQB�UG� ��`�:�'�f��m<�db�4[~e����;���R��``t�X#7�(���ȉ#�a�A}HaE�2����ev�)�
��g�G��� u50�S���m��u[c3t���[)e t
;^�_ߦ:[l�W���ޛP;�ܾsg�GG���Ӫ����<��� V�c�&�z-��WG��f���0���$�l�^/R3m<��~��C2�f�&D\�yM�~)�*�2J��6�_g��3�1-w�>�8Q&)�����g�ѹpO>_$mqE�~&�Au�=���f���NM�v�����@�[/�mk�{�t���/��=`��zL8�(�B3�iy�H_����fx^�{�Plś�SP�|�,��n!��k�G���Em6�-�h%����n�͂�RD)Q��!���TI���]V�Izg�,D�Y��������j�Ͱ�ua�Mu�Hj�l٤���ꬕl�<t�ڹ����f���ޱ���m����Ul��b����|ރ�[����h�u��pL�ͪ-k>#���i����CZ@�"8�l+�GU��X+�}:-���K�>��C�>O�:�m���(��S�b�0y܀o��Ӄ�����?Ozr>�h&���7��].jUH2��a*�G��^���Us���dp��r飷��e�2
P�$�vȐ�ZN��^��r��]�l�f"�ٸ�
m���v��y0 #fu�'��˰��X�o�V� 4(��h�x��
o��c=ү2[�H2�n#�뿞H�LF�F�Dd�W��k'���5N�"m.K��HM�ar��#����GW��o86�ԝH��ű�l�&ʶ���&x%�QhEG���p���� �=4�R��R��%ȉ�C� �"�i�=U����x
C�B���Gij�d{s%�O�|p��h��xܫz-v�f1Bm���'�qP7o�w�I�j�豌�h!Gϋۣ̚H��\,1F����E���.��1���mH���$��|A%^�����d�y�(�'(�I���5s�/��N��[%�_�jI�Ҿ��@(0�e�U����{:@x��/�cg�A*�����Ts�<�x`�囊��A���ג�ÌrR����,&�u��Ö���T6ޡo�T=w��S��t�my�����D@�*_���Tr]+;��&#t��m�1g�m�0�Lݵp s`�z���;Fn�,3$��\�~n�H�K����Q�}O�Q^�5�~��� Z[Įmp)݇�1[w_nh&oU�l�7�J�/[4����y���[���%Sf�4m�!����>� C�5��d0���X1�"*�@d�_w'�q���R\��7�cUiLL�>K���aަV̅��(;,��Y�H���sEK1[bf�`��Ef���Lօ@<��J��Φں9�^�sPn/]p	�	����*҄7�v �@3���2���ۙ�zh6�.�"'f�:��F���㇗���{��8���&Vy_9�M,�k�?�����3R;l���Ԣ�,���@̦Y�� Nz]�h���̟CJpX]��{h�Ƿ�O��%}�y�A<#e@�0�*��J�']��[�\9�G{��qx�y`����	�����}~�-);`�̅@�7U�:�ֈ=��V}ȼ*{��2�?d����8�z�{�k
�@���3
��mAz��+7	���<��â���+YS�ܜ�tM�m�9��^}��M@�:���� �t�N��m"�c)�w�����i�b�!�KF�&+������A�3�`��`L��Q��W���
�e市�z�pG��Д����͆`hE���ae 5�03E�zD<��~p��ऍ�+J�)�E�3�z6%�6(t�ݺ�_�<�д54�"p���d��U��Wު��
�o��E�>ѽf��q�=j�4ꭝ�/d�hV}���H�F4�ωض>��ȃvNv�n���XK�����q�;�ڽ��&��k?�L�/�R��;�i�(���y\��[�rU�˾"4�J�>�&!sȺ�f��[�v�~O���0���&I(�5�A�J�����<� �����������4��[�q�	��ʚT�&]������yE�sSrg%L܃�����ju���9$�ȹ/�qGm��`�=���ΐQ�����>M=�0�@��S�%��|���{��^��Y��xVu�Ѕ#��*�����uoXե�����GR�iG@B�j�"r� �i�DUxy'���u�|��:��	Z<<�5�x�&���d?~8��ب6����=�͑8���&*��h42����So�K;6w�5;��>X�o+�E8m"B5z��w�CF~��'��|���VI\�~k�2���=���������/wU�/��0�j��3x!�WQZ~�@�v�#�FŐ�]x�JZ�Զ;�F����F��!ve�I�bWx�́ty���R�}!������/b��ZF f��v�Dce �๯��h�v�	�/��Uܼ=���3ET��Ӽc4ǋ�?��V]"�^c��@�{�#	y�F��dp�o���i������A�_�@�Zh��n�>�k
�X�;>��+˩T-\��""n�����L�̏
�+���& �*���Xnѧ�x�uuz��;$�j�{z)1tȚ�sҾH���S�F/�!m�}1}3����s@Y�隟�Hu־���9E]�t��/�@�)*����u�t��b72���7L���ȇ���M���ˠ��1�U�%?�FI��j�X{�`��t�?*��_/@�C�HT�J>3kDB�|��!��]KzL%��3e��Kn%f8�
A��|�Y�5�_: �������vx������ (s�T�(:EG�`�$��R=���B_�cs�Y�,�,�.[p��u�=	j����Ȉ3هP\�]�&��c	J*}v���ôBz�`�J<�
 3vLw�h�:M-璆\L�\�9י������ڰ���,X�����6>�>0����4��Ԅ�h㈲0�Y��ҡ��ԟo�{�=�O:ٚ���y`Pj��t��#�ث��]���D0�5oM�x�t�Ĥ6��e��`%�}���wn��o߉j��P�R�@�a�ۻ	�@�M�tt�h�9ۏ�[3@\�i�U�J���D�gRԴᰝ��Ys�0�ڂI��V��Dɱ6=z���a��3�r�f|��_��X<����9�	���!A{���Ԏ��������c�6$��	�'�K���@����Í%�!CTW�H����~�6"сIN�P���*a�<�������Qr��z}N�?��J%�{�N�22v(NUU�H�g��ot4��R�I�-��o���-sֈ7I�~�X�����߭o}�E���v�9�-V�Z
}���'����⛵��_Ch�M��y���M������O-�VR�`�_�r�לE�1�D�G۝��P���L"��4g�l�yN�jfKR���\��Ugxd�t0[*��o6��\�(�.5����dX>-�Qk]	���Z/��x3�jic�ٲ�̡94�Y����e,-��o�D�4�|Q�Ǎc;ց@�����i�V ���s�j�G� @Ӊ:���:�h�R9�B�������:����Eb���h,PH�#�Xc|�Y�,2+_Z���$?�Yߟ$��d� 8��(��f�o-���w�	rw���&XL�D���k�;��(�ۃ�>��4�hOE�@s��E"�$��x�~��'SW�����"J��~�$r�7;���2;�H7��9�h� ��԰�\�U0<I���ʴ�-OD��C�bs�����$�Ñ^郲���G�}�Y�-"�)�{�D�F�406p˩�TÜk�*gc�y(=`
����KTlQ@?wR }��T/.�$�������o��n�!d����!Ù��t4>c�����W�5)�҂�3�����Q�ӆ�i��ϫ���a'i�׀�:O,�ϸ���6����p۔���'E&���-U ��������F��ֽ'�
�3B&S[���PG
`�{��9?�@�t`�aX�S]4�.�e���`D�ܴ��f���${k2�P�ƥ��1
��]��Oi���˰ʶ` ���)ߚ�/��w�9�ه����?M�Q�s�a&"SJ�%DK��O�TK����Ƙ8��>����FBF��+���+�\�K;\k�E{���P��9-��GRmXo���7
R{.S4!)����1�a'�>lv��e�L��~U��c�cU��%@&�i(���t�U!�E�-F���5l���_v��jM��ţɓ�q��dr؃��h��m����EP���{_��W[F�&~x��ʡ�L��}
�"O�;^�}�y�a����N@��z'Q���91#�\��V-pG�c��ѩ�"B�?��:.��{����6uΙ΂��eI��$�mvX(ݟ8]g�|j^�6���9G�ҀvA�R�tp�A�����*Af|�ꏖX՟!�A]�љ>9�V,��}h�=��A�MF�d}6�XLa93u:5��
��ʣ����C�W�W�D��¬��_1al�s����UK� <�"��+��Ɓ���v2u0�q��T�����J��}�Q �+����mW$�Z����<�ς�n�J�fΌڥ��H��O>y�ڗF0r����:&��'|_�LjJ|㈇�*��ܜ�ʝ8��%{_-��*A�W6�I�Iiv ��MD����Î2I_�Z�W6r:5n��`vʜ�83t<n�IS�&o��P0+N���CL���_�n_�(�}�Y-}�,L�B��������=$�@hXN�b�xx�-�`U��М�B�^Ȯ�(��Tu�j���P�Ǖ������oHG����y��.�</�C�r�c�w���:  59T�2�K�;�K��S�[E��⺹d������%<��������%����c��n�%a�b{��Q�&��D<_��,�h�R9KZ��%W�b������Ӌ q����^�Mg��lT�,�y,ǁ�iD!���3Ĭ��[cc��X�KŸן��l{�v��M ���Wf ��<�M%07��n�Iax���/�˗[OӪ��̷�ކ,7�����vަ� |U�3T�UR�:��i���+Q��2} ��i��\��b���D���	RC�ޱ�&�h��ek��J�uie=ߘVq��.�c�dq	b�W�C�Y��x����1���DRH���S��Q�iC�흺�LL��'�ࠂ����ǳA���m���<�mzg)���&yI��
#٢��E��Mپh%L�w���[`s	�%��i�{�CV�,MdcQ��{�c�XքY#�_�ID
߰��ȝ�"��lD��\��4�0[0S�� ����i�B��lJ����(��
b�3 V!�c�	�[Pwv1�v���^�Ox+��睫�ck�^�����A�mr�O.�O�+�	�����O�����'wpq���U�>������뀁@a�or��WJ�Է��w�:4����\��lVj2Ŏ���
��z'�^���fn�^���^��&G�5�"���~�2��b%Ͽ%T�t~���pb��Zv`$h=�l
�' �h��{����$e�q,��ݏ�����%b?O�(߲B?O�>���/(��G��I�⟺�i�u2gx��nƘ���*(�~^mƿ)��S&L#p0MȐD�,o���#=���2֏�L^RRn-ބ!���ޯp����}�u�/���GWXܚ������L5'jod�!��Y���Z M��m����-a�d�V�������Qs��f1�A%���a�C;L�H7�2'��	��	3��1�h�UO��zÔ�w�<Z=j�*�sT��
N�cɄ�aU_��A�U;��9�F�L�;���<�&w�Ϊ�d�zp�W�nbO��$�܍JI��P��'�T�IL���T��W��%yO��[�	��^G�`��`q�]����jc[�@A�A�	�'M�1,T�s��i ����$A��!�L#����c�����d��s^N��;����m��O}�g��}~�u�L"e���H�j=�9b[R�t���xO���ɋ�|j���-���E%Á����b%�<�gZy�s`�r�d�����>���gZ�;r8�T��Q	X
�Uw��l��݅���d\��8B��1�0a��#�� w�T��]��@G���6#P��'�ڿ�R�].D��l���-
�)��G��Φ�Ն=G�X��ǿ��w� �$[�0��1����:L�!�˪��`��ֱr�CKs�{���A�P:�ZG�F6��oB~��%��&�E���I�ܬZJ~���'R,�(�(�m��(����|��̻�� ����͢&cs�8({�V�� S^I����@2��,}�����%W�}�erO_.Av�<2�{��i�ll���e{�r)h�o�P�Ӭ�`��>[33������� ��b���!k^�A�'���wr�
r/��aEg��Yi��j�z��4�B�G��U�I�
$���[�"�$�
��m�a��O�Q���$&�r��y �^θ��Ϸ�Ԧ���A�m$��193Bs�6�"��E�n0;���y��_0�Hw[��E���_���6�c�/����lj��<Z�u��U�X�FTβ�ը/ڜK��@T��Ŷ�WD ;)�GԴ���J�L/ͧ�ZG�0�G�m����[;;�b���YY�>�^���'�6y�3�{�n���Q;BT!�V�l�Y�
�h���G��_�*n%�F.z�F��eLݺ�O�a����u�\���s_M-q��:ח��en���-�0��b^`,��5J�;�V��c�rU��3�ze�J���֠���~�*�p0��t\I���Բ3�=����#��=��<l��x���5�`q�
ᣤy�<奏�Z"av~�hi��C�Ü����tf!+į�]B���&7q8HK(˼��	����E��5s���|rM{�� �Z���aC.�X99�L��ҷ��7�����*�bD�h�7~�<"D���j��(��ZJ5"W�&T�T�C��o�J�o4/��,�6���,�M����Ă�=t,ۙ��0S�UT�� �y���-r��2�5�&��c$���]��(e�J���q8)�E`.w�]��2;����_���@%��m_��b��8�{f��wNp�!�"���Tk�6������!�wi>�H���zN?��}�����1���PA|�Λ���K�Z����o���B��1/S�G©-i���T�������s�@�y����+n�"\@tp�f!a����E�%x�[?\ٓ#�	�|*�<���d��u�i����/�z��t����6# �F���@��:q�`�!�Q9-�k7Z`�=<)�%������]ꌷ|��x���}����]ҥt�¯�\R��_�[.�`��#����jX`�Fv*}o}�/ښ�'
��� �?�˒|r@�P�ŵ6(H����I���v��(0C�׊�k������|cYJS���$�Hͽ��:��#\�M��L�]H�T[�R �5*�q�z]��R�?<�=l��^�)\�&��,=��#�#�	G��]��6�)T�	�{TgC�V졜�1v��ǎ�U���Y�$�âY������n&\�ӞA�F�x�o-�6�[_�*��.���g�ѕ��Xj�U	|m���l۸𑲘�?�z<F��0]e�ֿW�_��?v�H�[=�8�E55�ޮ~�T>�4��aQ��@�u�j��}筡���C����U��FU�,l�|�1� s˷�.c����5B��u��D�Ag�E�Bj��ә��U���&�mB�%|��@�3�XE��s6��o�}��y��{��Å� �B6�8)z��4"���*q.:������2��*�Ç�[i�����;P�;�ݾ*��L������� �ȍ􉡌;�JK�Tp�ş1`B=�D/糭~���H?k ��r'|�%�@���(�~!��6�d��FJ��\w��$4��kDStc�g7�C�	��+P[pv[t���/y�w}���̚��j�6�CG^R��"�-*�ߢ�N�U�cD��h�����x���6-"���c"x���r*2��.(U��Ӫ$I�W��&��?>�Hr���8mC��!%��L�~���f�d���2���$����S�'`ȉ}L�D���Jw�i_M�]��a�/��
Yҭm
ӂ;� �LCui�ډ�2��V���b\�:��J]�k�n��J�%���->�#��#��ۨ��w �d`�2=N`e�obW�?�4S�V�O��o:~�n����t��Q�	1��EW�ks,t|�Sa���G�@�$g���俵�'sVY��m�U��o�g�ӜM=hl�u��0���]�{.�d���q� ���'4- �����9ĺ��>���5�8��25�U�p�)�+��D�0'&�.q�qe����v9�HR�U���xa �/i�
w���86鑾x�y�vD��~���Ӭػ�5�y�$o�Zh��Z��7�/�lhƙ"�Q6��� 0��bÆ�t;U�;��
�5v���3�	7;��Q�<{S*b�%��_ W9i���˼��6@�B�
���8��������%�Ը���|׋��a�X3\�}s���>6
�9�^���#���{B����@�V:��g���ܢV�>!1�� �fqݬH<�l�
��=/�\X�0�T�l��������6޿n
�w�ǧ5f�ٖ��ľ�y�c�ى�&�ed!v_!��t���K8&!����O�dp�HO P�ԝ`�L�΂�T����ޭ��Eఀ�oI�<���rb �C�.$\��Pf5��n�7�Y�kd����U�(�a]Nkl^�ݢ���c����@��X�w����N�G=/�d�Ce�yH�.��&�dN� A����4#������#k�۩�T���EV;��'���!8#�B�e��Ch�B�AS̈́ ��/.k�BE8�F_�CD���w��e���P��|����U�?��@u�!o�ߞs�}��pCz���{b���Xf�L�&2��ί_z�Ȭ&:f�$��X�G(���<B��״��!\�UŁ�f�^�k-TGE,ю��3K]���=GcT*"�?S�ʭ�h=J-%��%���+[�I ��F۔ر�����Y���ge����1�Ec�}g���5@�-�n�F$i�)#�x���뼠[��mz�׼�:[�:�[�u�R��4��U��|R���nq������l�b+$T�Q+���h=h��xf� |W��S�-�ܧh/,��o�L��3��?K(F ��\ (��P�ȳ�Z����u�z�"���!U+�!e�*F�����B���
����;�r^����c!�p����$�(NbDr�/[r��P
���HΗ� �qǱq3��za������#��r��Q��0�o�IX1B	7���0��N�c�u���e #
۾�~�n�	q�~a&C�1�T4B.��Y]ˇJ���:j
m6��;�`]��ރ����HZ�!��������K>=4f�P��J�$��}�!դf��I�|�3�	o������o�zTlp����&5^n�DS�%���;��و�/� I�x4�[ud��h�,7 2�ь�H���w�f�Ë��	Wh6��8]��R'<��BY�#��d�!��� d�l�R]���>B�F$T���9/v��)'�JEm� ����g����c�n�_��W���nlY��k�">�u܈8Y�ǡp X3�1�cj�k�cȈ+xy��Y�S >=d]�伦�0#G����T]#���(�DH�2�+O#"�@L��a�zh!Eξ�4H�k��Z�0�kQ��#b���גi��W���Vt�e��]=�Q]A'�vrU��U�dh��ՍNh�r���i��W]r{��>�g�n��mU�Oj6��? 7��q[�tE]���c˓2�[�Փe��a�F�Ѓ��~�X%��~;��Jۖen�@�m�jp6Am+�v�>��$��T<"% �9�7��n��á�
��%�R���S��尀����}n=��^�gЬr�K�ު��tw�]*֤/sV#M��C�v@jbe�Rf����8-3�m�.�r�x��{��7`�U�,)�.1
y"�Ta%���!�Y���	���f�LX��X/�FԶ�ݕ���h�3����C�	�������yH��P��`QJ���������6�H�t:�!�_���M���ں���9��j�H���Qa@��O5F�jU
���-��H��Vca�����}ho�?OYG�vjgyn׎�򅪋�6��&5�D�t]e�¢ϟ%rEK�B���ȑ�AſFLa��$���k�,+Ƣ}�2��T-2@&��D^�,�����="'�y �M�ygcF�$��WT&	�V@���_�0��}Ы������.��`��}��`�J �����v���Vl����(� �-����7�ϘR�`���+���=�bظ�h��������4'{싏`��j'Uwߓm���ˮYJ�ų�`�x�,�4��z*y��6A���QoH���"�@��
�豣}l��+��X�{��I�E��w����!�N)���͙oY��ٻ�d�ұ�n� ���፰�ن*Yl��+`�f"G Q���Yy��)G�hg�~���r�8h�.�SJHN05�7�{�I�oG�C� ������m�[����ao����o�R?߶|w.�(^���'���rB�k�QZ��]	��°o��O~�ޘ'�A��X��e�x���m�����#��۝T!�Ƀ���ؖXTB0��a�dNz��*�de@�b��m�W-�?���4/��x)�,J�nʱ�&�Џļx��#�Q�^M>�ɽ�|9R	�Tu�w'd�A�a�V��w�J�j�&������31k���g�i���X��1�"!FZ~B�(�����td��?T�qX������T5{��堪�o���A���QϬ]2L���V�m��o�;�WO��* ������d�d��i�h��?�O7P5_�Qt
@�Z�j�d��Ig���"z��n	*�����ooĲ!��������0c��<�RUv�f�K!��Z�ۚ�,�S\��DH���Z���#�Ӫ3��f��z2z&p��=�Jl6=M�}�s�/�S��u�=:x���d���`����C��{�zO�m��EV} �@�L}�t��'�G��K�+;zp`�{&��F?>�޿S
U;�#�5���
,#��ey���R���R=���^���>�Y��J������t%_˙�������1�?��c�Q ~�7KS��h��?f�FI���E~F"7�)g�R��>+z<��p���<Sھk�4'��8ȵ�R���o�}���@���Aߠ�NTR�\D�Q�m�6�T����[�TX�c��Pe43t��yZ��	T�)��H�r!:�%I�1�g?K-�^�j��ؒF����-�;�\���S$%�c}�_w�����˯�b�n�È�/7�{6�;1Ż���,��'(d�	} 8C=fO[�e�Xen D�,u�ɋf=���	�r?92��}Ii:�`<���%Ia�8j�b�8('K��?�;.�2 A�`�|�2WP��S�tz��-�-u�m�����Y6��Z�12��UM'0�����#=f@�Ŀ*��Ȕ��U��$��32����dV?�UPU���J�eã�c��b�{�m��S]Uea}���=T�;H�R^Q'y�Y�<�����-��� �:*3��涥�aD޳Y��m����]�>����T�o�HǛ��Y�E�����h	~�\��r�^�-H@ޫS,�9�/k�bLA�����2]��T���R²��E��"((֣r>�DN��3b�L����Z�:����	��B*�X�1O=+��-��C`y�|}N`�:ab5l|+�͉�R��F���D�m�P)2�Z��>N�:�qQ~�/�j���0�[Y~�
1�~_Z���Ee�&��Q��Ҿ��7;�bv.� cC�m$#�qe�.f��|��c��lA��nޠd���oK��{T�wq+�/c��<���O����s��}b�c�#Ð�|}�~�n�Ʈ��@�BJ�c=-��v"��[$p>7�CU�{��l� K���I���l���Qm�r�o�nf�j~_P��E�l#*�
�H�($�퇝��ap��Dl�i��!�m��F�hܐ���~)X44�w�T{���?�:�<%����d��=!�;��k"�D�@�dj��6�=X7<ٟn�͗�����C��e*��	��C?���V�h��>~�2ۨ���*k�BаQ6/$´�
�zP��76��G2ɣ�Ev�
o꾆�b������m���Jd���� ۹�(����(cŇ�6gɢN _ߔ��!4Ą���7-���
 ?ZO�9�����0J:�Nٱ�:e_��P���c�W��'�����_����;�LQ)
�sZ=�-D�w�.DX����G���H�u��D~wJ��6h�n[2���V��������%�%�o_:����8�)������}FuN�q�����Vlr�S�K�X#D���|	ǎk�Q��wO�tY�N��JlsG���X�740ާ2��W��>��Z�1���\[6��w�ϵK���0l�ul�E��)}7��'R�\o��Fj���`�LЍ����$�z�aRf���w
!J�4^g�9nF1�s=ۜ,�_8���5v*���gl�D�~�S��3��!n����Ǿ��s*�����H��k�Àׇ&ibt^=�����5� ��o@�-��.���c���|��w��o^�V��U�-�<�S���5ojF.:��`�bvpx�
�h�"c+��0����Z��P�,9�r�Z/����qT�{�Z�aZ��-��>t��I�$��(<_V���&l8HU}nJ�Yp��h �iv��q�<#�i�Tv���p�)��b�u��l�{���L��F��B�J���.���½�3;�ɪ��(����j��E6���U�n�F�����/ y�Ĕ�T��KO(cE�ԙ-���x�b�J��gr�ɹb��|���Ҫ�soC����~ȟE'�h)|h"����S00���o�z���OaF�%���I�^\�2.B�0KP>�>��͉2١L��l�1k�faR��DH�lH���G���6��
헰�^o�x�^�� S���[%�Uj�ީqr�d?�~��5�q����_ ���i�Pm
 �U]\���z?��[M=�J��n,.ٶ~w7P"*Z
'�+RJY�c�V��V8*s��'VS��f��%���=��\˾���}�=�)�k��gM#!ă���;E�z�]���K�8L�Wn�m~����b�G����,��y����f����@g���s�&���D�����U&Ja�8�s@I���X���y!��-x9�@P7W�A��*�-�0��l�V)�&E:F�e��T�{�q��6?�x�m�s�\�=�o�Jo�g�Ű�E��l��[��Bՠ�\�)����a���G+�_��
I�H��帪|�[q���"fjj9skH0�b�Ħm��D ��y��ްg j%9�r�ǈ �F��1�п���4��H��/4���X�#XP� �΂��/}�'���$���g�Zx�iu��W�AD��Q���j�����n4!Y<5�,��8R�`����&�,,[������ 4cL#d_DS	�n[m&2�Ŭ��)Y���go	p�����*ns�r[��=& J��5\GU�[3��.*3[y�!y���;ݯ������Ċb}+\��OE�'�C�9�h����r�%>��&�3�����gtXIΧ�:�'����WӮ�Iw_a���Mح"��"���Q�U~TSB)��4kv�W������H��m���%ϻ���.�Xt��Sm�B��w$�(�;����1��*ʈ��O��v�K���5 kF����,�鏾J�����'%�%e�P����w]D(o����72p���d
���x��,]e��~�yg�8"�ie�&փI�'	�^�F����P���}�8����u�AA�C����=��5Z�����z�0������]��s�$�_Ix�.1>2���}Cd5fV�X��ЯU�7�
���wA����<�7:�'��E���mf�dx�P��`i���8�-�� �@��0x������P'_b��J����w`��cvp���~��V#0��X^�o�C��8�d�͒��ܛ,qym?]̖?����·rL����N�ۦ� wZ�����῵ռ���	E2?�G��~�t�\�(���p�u/����s�����Ϊ�<KJ��<Zpt�5"�3o$4$�gCXس��^�Gz�D��۞�}����Ń]W�1��6���Y�Ihm|����dZ#F>�,}��fZt:�[i⭣�����!e᭔w��mN�a��R�Q�~R�G��^��4;�h���b�KzFy"�5;��P��ՠ����eI��Qj�݃V6�k�9&,�D8���HfX{�}^ج�¾g:��P�=��د_+��b��L�N)���z��EZ�?+�e*�,�Ӵ8Tב_F��c �#Ԉ�%4B\G��t�����,6l�"�e��d&�Fv2��oX�����CS(]CL��)�r�Z3Z��S�hH0W��H �=w�z�����`)þ��Q���~� Dw�0�}L����dT\��U���l���ƹ����j���������!������b��!V�D׺�ݾ��{��@�2��0�'��M*�qS$����]��%�K�+���������L����ת��oWD;�A@'%s��8�Y68���C��������/Q0��׈eȠ�c��%���Շ5�0Î���Z�ԕ��u��|��:M��P-Y�3G$+����G���'�8����g߁/�@z/SU�-j�e[U��w�P,���k0��ɣh������^Ã.9����O}3,�6a�:@�´&���Oq��ɘ̕���R��o������%5��F�g�A�sZe\,�;�E9�-�L�Dj����A�,1ֹ.�,��c��hg[�"�Ҷ\�vp-�ʨ3:�6���h��{�L�CPsc��'69�}��Jp�GtZ��H2[�Zf�W~��V׀�ݦ]�ۘ�������吓!}��=���B�� s����I/j���2�ܐ�;7ƳhN�	`;����,�A��}�v�,��̍�´t�y�����"�p���MT�H��?w ���u~����]㜈N��<���;��9��Ӊ�&I�������*�Q��[]�m��aY�i��k���,$�r*1��s
/�n%��L�����[`[�]�]�*�5�2���=\��WlEI($�<��R3����n]�'���F�d�؞�\��4dC�3UģXf�U�����䍌�cQȯ|���ܭ
tU\?��$6+܄i@���lh�0���V���]����#�T�����f�V���K���T�B!���zʛ���(���@۷x�������� +ڡ�*�L��nӪM���'��|��Q.'a�ƉE��M��X��l�-*���%TV�GV6��s�5лQd@�k%^C����1�P�@�v�k�Q�>c�3ʍ��W�j=1�&�����$�=��h�?��Ef��*�f C6wmv��T����K���)�Z�^��3��\z��LΫN��]�|@�����ȯ[���}���Mk��Gپǉ%�#��J<�H	��+�b`�L�-b2��x�r�1$��C���L��:qp����d�H��M@�"�*�n�R	���M�2jZ���u�+A��[$okA�\��`_�ޅ���z~D��~ݰO
id��!�>{��=H(�;��8!<�bTMbc��V�dT�[BՂ�	�%�?�3���Z�+�j�[��h�)I��u���'D����3P>����@�o����R��&F��aγ6�3��J�G�F�=�`SFʎ%�3�"�mN��$���_�ߒ�=%��RKN���k��s��Q&ۛU�ȴ��j>`�E%�Uf��1܃�Z_`�.��id���3t�Vܳ�Ac���k�R�c�F�#a�0Ć�%z]��/�j�w���~:&=ᤧ�d�A��q%���>.�h���X�J�HHo�V�v�����?�1�*ʞ4��жf#gE������k�r����6���;9c��l"�?@A�W��?��l.��������讁�=i��N��O�s�S�PΏԯ�5@���Ds3�6� �g0���B���5���`�	��IK� �h���
����D5�z?���?8��s�&�z	�J�g�7�Q�I+ԑR���L��.��9�~�4���|����\�xq{.����Βq��P_�0��v��ތ�ުz�9?BZ�gn��J�ܖxڱxa��|��G̱��&Wk����f�4_��#Kl�B�!�UX?�1�vݺ��X��W�F*�|%?�D�t�� ����^R
c|��s������;8����L������QP�C/�Q�`��)WĄ�F[�����<��T��Ԁ�$8N�(�ECR|��@n�m�+7��6�B�����@�� 5�*	>��ur:�JB���nx������杽@=��i⾗|����K��>.h����Iu[bY�P��-dx��l�N��
R@}���WU��N'𧞷
��ژd�ғܷɂR��~&Xt�늯Ӵs��#��	�'��5<P���M'�Ù6�y�i!�!g�(�|�J��> 1O3�k=���
3	�66rǛwS:4��Ydj	�u�;�YZ���K�(|H�G���<lv�°y����m�+g~r��W�6>�<������9B�_�e���7�J{(���}wk<Q l��o�6�}�5e�تwũ)7��u�M$�V]tg�1A�=�(F�����Q�6�ns1���gLG�%��;l��IQS��z�8U�ې�(�_�>e6(�i]|�n-��w�>@�$b��	���4cOs'�`��?�X.9�r}y�pn{^�ߝ�J�8������
���$s�Yh7t	��Y>_M	�P��Q��rd�9z���B9���6:.������c�:]e:��i��+�+rf��o{o&cZQ7D1�
*��}����m�l����h^O0�0�}bt�hb�z2��X��-�C5�b1��T�85�A�����o!!��'5I�X�q˽�H�B�I�?�$�f�uq�n,!�	���]��]3um2�>��(tf�R�\y�65ej��9Wr�F���኷���h8)�B�$?\�=��U��,&�ڗ�-���T@�RT6>���Qy).���5@�x�H>n4�ՍN�ڄ����/*n�`��?w{I�ٺR��G'��9�ɪ$��D��N���d=_]�|���U�
;��mI��s�'h-�^��8۠q�H���e��h�;��vG:��r�b��`B��zyEt�C�4٢�Ʌ��3��Z��O�g�qO ��q?t�{yxR;q�'{��"�(7������z�96E '3v*G�T��V7��@�=XY#�^�D�A>2r�b�j&&O���v�6�������S�Ɵ.�s$;jFz���q�3���o�(�߽�CFFX7ۮܕ������8�i�����xj+�#��q�!Z�|��m胵.�fB@1漕�3,A
���3so�H,�a�myR��1�U�4%F�����������(�;h<
]Qo�;�Q��@�B|��J�lxI�mH�S�T����;� �{�-��m)X�cRnEVĸ"v�a�)���z������{��=����d�����t����w&�����Ů�z\9e���+N�
����Х�?�k#���*�u�#��X��{��U<&W& �	�� IU8��&T7Q�����ki�Q�LȺ��;�����k1�ٿ���A�������Ε��3�B�ޭ3SDT�VߺعQ^�!֓���w܇Q4R@+ �]�mu�`]W��[U�{��Kf���o>2#g�Ԯ�kaSc^�Yx�i꿪�78���}��X͞���{bz�����-������k#Պj7K#�)��~�+!'	VU��BKy6�!%����eS�5Y�5��i%���A刟�S������V³4l�%��j�(c8�=L�*7�Z�\�Rk��&��c��GǮD��G>�?��l%g�:�/�"OQ�5� �Ngi~++���1��=�+�2�<%���=&�u���CyE�/Lh��9�FBWe�Z����wI��dq�(y�yJ9�I�WG� �Tp�����\��ʽ�����ߊa�VX	F�X-_na5�ı;wG���`E�7��ZV�	���9s�7i�MMQ�����@�vaԣڪC\���K$�Zވˌ�H�ʖ���[�'���Bݭ{�Ckҙek������G�bΔ<�p��B��p=�YL����m��.�ksw�����Si�?:�yW�;.��8ϧx��@�@𢧃��#�U79e�;8Í��$�H�Y�~�&I�͈�Z����FԱ��%N֞�7	���P*�O��}P��=��h����u��f��9`�qU�&�p{�Q?�q��˲�!��M9;;2�I9\�'e|D�w��:������վ]7i"5�&�m�*��P/��Oc��je�?v�*����Af.�i�UH�_�� �U��KI��1į�%c�P�3ٮ��>&�A�"��������Pv��R9BV��ʻ�/3dx�}� �����s�>c�Qc�Bk��Y�Žq�|s�WiU��9�5޲��뢹GV�!��!�,aI�ks_R��-��vP�ns��g������"�I��=X�n�P8DY��P5c2w
B1�@]L��:�6��-�\EY������j����@W�H�}���8���^���&�U�/(6`�Q�c���#��&���e^!7�3���M��F�N9��y�i\�g�hGl��EZ��vWՌ�dX:���|.z�!�֙2Ը�s�\�XҸb� ���d4��p����)2?Jdoİ\��\7ق�����ȶ,�2�ki7��}�U�v���5��c���є�Zхe ��#��Gl��C%��h4���ӓ�~��/�^|j��/6�D"��F����'^�	��d�4D(����5��%{2��s�|�W��8�/������	ޠ�ֻ��߹5��<h���x��]�, �y��Weq���� ���Z����q�������E��	(ow? �W����sQ|{W&���JO�_G��*4}�N����ɺ�����`��={L8��viH��5�{�.<�\�}�U��&��n1	jՋ�-�Nvܢ�f������`�n�.c��6K��S'�Ƕ�{S����v`�J�'E�˪V��{�d̈����I����M,�#v��b��� wX��>�L�}��92�J����!��
�cJ(�j0����H�^EV�����`��Z=/�Wcʋ�;�z:n��JP8E��m�v ڑ�dG�ǘ�$��96l2�B�F��4�f��ߗ��яM��"��Pԍ��X��|��/��0$Ì�Jz��&�����M9f�J�eh���K�z�c
"����ޛdt�����ݺl��\�x�[:&��xm�������_�����;��#7���tt��9�tt"��z>[��x��W�Y�mnm,bJ�r��Zəha�H�Mjb�D�œ�^�M�3��K���Ypd.�[��p�q�&r�q�z��T�(!
�+f�4#��Q[M/	��eO�A�Y�	�x)��sh(S���F��mI9��7ZD�梃�ز�f�-%j*nu��Ib�Q֜�l"��[�jJd�S�UG�β�紐��6�YۉO�Áe��U��#�݅B�^@�]��TR7��F/�o
5��!�5|>�N�	x�DA͂w�^f�4|C���B\,�w:�(<0��p��!�lc{�@�ɉcJ>�^_�l��V��x���a�.�u7�J�2�	-�Q�:�����X/��Q�r�&��A���-J���7�Y3�È��]Xb,���礰��ȖP\e����5S��\���8�'s��M��6ύW �Ֆ.��J�����v���Ezu ��a�d��{q�P@qd�%�s��{g�/���g㺯Q�Zd��Q �=<,�`,����Y��&6�1Ʈ�*uI�]�g
����1.��l�{�s�����;�DyP3�Q�-��DBi�@<m	� �+�O��p�nx�@�����gk>����C��tG��ex�Ux1���g��O��n���0��$ݭ9NBm��	G����1&X����'�@��kf��tH����bH�ŸU���Z0k����n�<9IcncFz^$%��O�J-+?�JH(����	�_}]���sO�Q:�f6�v�+����U� ?W�nԞ�X��+¹�To��Xk��X&��t�R�u]h��gIv�bD�6����܌�>�Ѯ�L�[T���?&=58B��=!+����<?e*nf|#�ݯi�z��-?�-1�s�L�4�Wdy�T���]��O��DR͜�B��H�+�}W�T����v�&��L۴��ĻF/�W�#4\�%���o%��'>�F���t�HEV��f��4tϝݖr�Atk!�o��y��WC"�`G��~��+M��~}�g��B�Wܾ\�*�f��Ⴤ�^'����{�oY,�ɲ�8�Q��j�V�?(�)���A8SXa
��$�j(�w�x�m�5�vc�ʊ����!n&I��a��&w���
$*o�t��=LE�o=;'=c����-m�R#�nޢqϧ�ao퉓��p���������_QgYl�x��b�^���4]�T�+xx���N�JW��Bs��n�&ĝyDbp[,�3�c�p0+��uC����9������b�J���=<�mj��4��:*[�L���]וג�iz�})�	YQ�nѣ����-!�\a�����.��D`���g��)��kPo��[�2����������G��4KK�ᡅЎ�C�c�L���3�=` �ѤB�g�i&�0e�
�0��A[)��WC����Bm�w��#i�1�^ ��@G��H�!�-"���\�9Rqha���Kli]V���3��7t������	�K�����8���Q��#L40�a�t�Yj�����Bݒ;��)<�Gp�ኮۊ�	x���uUPc4�f�p�Ǵ��h���e�p�z��۟p�|����x�|ta�m��okp1��F:�>u�.GK>�gG#��(����D��������U�^���R�Q#��*8㴮Oz��z}4�Eb���\Z��a0PE�/�+��x�1��4tɸ�L�c�|r�<;�o,3k ��3�P� 3Dp;k���?�����q��k,G/D��3���8;�tAz��Эq�g���hV:��wk���n$zoB��A�C\��gf�J����DI��!���@X�����]���"/�Lf���n���e�ڀ�6�����r��.�i
IH+щ�h���(F6Z�;�T�i,��π��O���̂E:�"��9Ӵf�Q��u�{S4�<�;3��w"��Zy� xG��a+�Nn4j35. c�F�:�-D��*�u��<��q�h�}6�~�!
�?��u�M�4��H,�Y�9k�����$��������O;B�p�)�4Z�&�������po�P0��d��ҽ,���������D!��hM�������Ф��݉�,�����G��J�ˋ��un�?����hXm7�����4C$#�*�-��1���5'�c����"�t�������ߦ��3 ����2�-�!x՛���9�:��/�,^�㳥��Iv�g�1�/}�mMu<�<��UO�:�W�o��0=K$�&x�J/�
YldQ8�dr�tB����p��N��x_��(���JJu�mu���x&�����<P|�����;��/n�9nAʹ��{��MF�j�?,�=�֖���ī��{8�[(�XW?b�Pd�HЏ2tF�[�t[���$��-��zT���(XYwi�Z]ˊo�/+���uR,.����l�asZ)ܭ:�Í���2'��@��܈�g3T �����R�ҚopU
H%\�5ʪ��P+�}L�#����5gi������G�M!V����[�9P�Le��+���}�\�Vpb�d��Y��f��J����������O���V::O��˛@a5��QSd�d�:}�=��f�W.��%$ѯ>�����"��\D�|���;&)(�ڽ��h�bv��:Ë�ᖏ�<#��q[s����ٍ�E�U4�NB!�m�[��%�/�l0��e;���<�Ƀp�/��tp�۳����A9Z��3����~��j���{��-Գ�Q��(*@�T+�,G��N+�Rx���dy�!��d��A6^�DV���f�f�]�k����MVH�)�#�G��ѡ�0f �i"a��_��瘨s�����r���>���r�mg��'�a�q(�,8�S�l���������/�~��Ν[���)�Ϳ��P���w��Q���׼��^(H�+�h�7����La�tI,HLd�I`�~>g`%5[����s���]y6bR�f���.�׮�ȅ�_G�0���O]\�2{�������l��	�����v���š�~t��"�˿��tV�A��є�4IZ���r=���\������{r=RK��M�?��B�d�#�7M�,����}8����Lz��}AbDѹe�Y��&'���~��%v�*�.0z�n�c�F� N��u#F#��#]��u�b=�=v����1�2}�>ϙ��IF���`�Ԕ}7a,u���8��Ca_FDgP�[Y�k��
���y�묗�"�њ���wak�FY0:�+Z����e��-y�Y9�@�����������(�vW�&��R�����-�.��+'�����c���U'�44���3��jm�o|N�$�t��h��s��=��VM��N�^R���udp0Ś�.�2��J�363CC��tG�~����?�Y�m����v�_F�I�?[�G�H(�*�{9b-I�~M��[�v���$:��`��r����w<ڛ�t&a[�SL%3�"�NQ�sh��gȭޠu�A4�ٍ��4�U�&�l�F�,:�3��yb�{=����j��Q��Db�� O�	���g(L�`o��jK�����.6b��QGb�]��
a�kf��~&��&��e(�F,�,�б�~G�px$x��!mcukN4�k�!`��fP��� 6��Љ���7��ܫ��iƢJ����{���C���>lB����B�M߰�V`�O�Ћx�h1�\�b@�0�]}���2rO�	8Ak�<t'q���F�-};ʂ9sk��]s'�å�M�A���)���L�^� }CQ6b�3�Y��w\��&���=@/����R�2.F��L��M�~���+ �Ouc���j�]��/g3K����Z��U��[�qU��@�X�wO�ڋ�d:��8�p��W�wA���iP��\n��Te���q{���d��߈#
��]��:엎�T	eT-�=0
��!��׫�q��E��m@B�I����l����{��WM����\M�bc̛��3:f2�=���SW���&z����=:3aA�j�J�Sl	r���0�hi�һ���AҢ�J��b�~�̂���>����")��Q����(����dK�������o3���6����_@�Ȏ~r'Fު�ˋ�Ǒ��V�L��k$5Fz:����:��g����uHY.G��$�4���"��)*�r*���[��Uk�&��*��+X��ӻ�_�^�x����8\���,�@�`��@�q���f��us���˙&�Y��}�!��}���dA��"[�z-�\�#v�n��&R�F����=rn�G��}r
��#D���qm��yd���^e 0�E�#a8��_�� >=p���i��r��
fk]�z�2x{e�Zo�K�+z�g�QR��'������ud?�U��S�x��8�e�J�@��z.���iݪ�+���h�o�5+���i���|���6�Pf��L��ZU�Ago;�E���9u��p8��Qb(���	t�`����g�g�д:�^�4���lE��(
YC�1�,z^�@��8��Iz9�\bp�#�|�p�֟ʗ �|�J�щ�@�)J!Wڔ��7�G���V�[r��7}_`��M���������Q���F
��$�H�e]��6k��S&�k: `jCqE��3"��]J��_JQ�C#R�'�7�k�(�^����ʏ���SoS.Sf��%^���#fǞ������N���4����s4��л�����-m]�U@}[�5�k� �f�`ԳA-:!��P��-FO����2U���M|I�{��S`̞Zt���t8r��v���r]6F�R�Y���cSTW.�Kߠ}]Rn���㿑���$���ߎG0�l�/䃩Ӡ3��/�F#��G
^���2t0�6W\C��|
d>��x(t��D�L�P[�o��M�� ���Q4;��D,y��lZ%g��+�f=2�/I����d6�h�%��9�j�j�0:��C�b<ϫ(|�h�E[�)�SzbL���U.����h��s�հ,�����ɍ�e��͆��K+:���\��Ȱ�3R�T�n[��DCnj��]3b���6w;�L<Z�/�Qآ����`?`*��9皳�nc��	��ͧ��+01>���ک��X)�lkr�E{���0u%ᵈ��G?5�k�]�m�:b+��y{���34��0��l��[jZ����ؙ�A�%�h�GC�{Tn�x/�"ǧ�m����?��!Ⓛ��ɼ��;۠��H��H�9�������7;t����H`>`���8u-��=�#h���5jŘP�^���~ݏ��&B^���/G�[�ȫP�A���;�h=D����o��XQOS���,��nK����C�si	�s�Xo{�6�~�(��rD����V/Wi�>|b�L|�N�8�Y�I�םWG��4��&����~;�~�s��8I�D���O�3�1w6�r���ȾYX���Yv���b}K���3��m`�l��O��f��iI���i[y��`{��{�b����Mf���/n���i��"��d��R��^\����!��<�[�\�Ӳ�V� ����(��r�4�\���ֳޟ�*�zW�QIu�v��3fe�,�'#�G��q�P�jtv&f�4�;<�U��ڰ��zX1��W����"^��C�m[C�U�����[Y����j�=_Z�y�a���b3g�u�� ,lj��6��Y4�!!Ux�6Ot�I��c��`� 9e�4��+h�����h��Q�q5�<��%L[�?%*/�s�~�������m<��Z�����q ]�)(�s#�kXS������'���/��k�����	� ~�SLL���n�ͥ�A�&�;陻�j�/>��І��h�,z�`u+��컱�]���$��)؛�3C C2(.�I������X��KC�����D�?@�����ɳr+�OF��إ��ĉ�;a.l�H�.� ���	�W�(��+�9᫵�$!S�
��)����ޢP����ʮ�N�Ej)ٖgCs�&Ÿ=)�{[u�/C�t��/���}UqY/~����o�9��mQ��b��h���W6zy���>�^}�9ƍ�G��O���05yn>ҭsGd�d�_U=�)ރW�����b%�e{eb89� ���y����~�wo�+�]#�I�:|Y]�~�m�������~�\��~�cT����[��#?��ͨ��2y�HN�>b56Cx	��d#�,��z��8ױ���C\'��|53=8
���U�3� �ɞLԇ>�θM�qh��-a�V����dY{B]>JFCK �'��I[7��m�,P+���n���ѳ=E��u�]��v@ȉ�E͟�r�o|Ϛ�)7�����6�n	AĽ�Jh i����-�9���ٞH,�T�n���̐�VT�hWq�뿥s^x|�h<��g�a�ѫ��.B��+)�y��.%�O/��nv��xg>?gw��C�������lD�}_%V=
����N W�F3���V9�8Л������=��̗�E��������K��u�5�s�t��=G�Ǧ���z��Y-B@�7= i�ԥ>�ѐ�w��#_���I�Χ�f�8��J�K}h��O�L��m�)�\P$8�%yp�>��M�
���V�X�֜E�'���d3����<������)7�˟��Wk����0�J�2D��ݣ0-��0�Y��y}T����2�\K��pL\�A�䱸V�,!��d'��-ɻ�%���-�������ꌷB>���K��q8�旎�t,�Px��n�S��L��6�Z��zU��"�������?O������,42Q/��Ѡ&E`��~ڊ��/Ֆ�v%���5|\'�\~��睫X����dú��|W�ܔl0�~����̭��)P�{�?�E�����뙑��2�(׭w���2;�t�?���Ũ]*�|��H 	vt�͹��p��z��0��1�\�0��������%�a�P�G|��Ni�a��cg@�Z؝-��U��/��ɯ��	A"w�-M~�˯@��F�4�G>|��I$<\+l򹤐��E��	�Ïl��5�J��T>͆����uaI,H�.-�1! �O�~��J�O�)��J�	˪����x�B�7�s�w;)���z½X?��F�2״$B�=���]�坌PN`׈O����ۦ7O��8�b���8�D�bN*��R����BlUZ���*� |�}�D!2��ԘIz����}A�%�^2ɴ_M�g��c����ݶbL*�jmM5�Tc�`����a��lۨKU`P��W�S��v�A��) 50��-�^����)��1�8f�49^*��pP��k3�tk���6>G��B���#%��I,�EQ�cd�J���oYŋ�6�&@47��?��a0������+�(�u��P6)v��5L]B����-�9�MRh�!d;��H��~�!Փ~S^�n+JN�̀�%���(�C"����x�,��u�\�w6x�Ɔ��=��@^��g_P��o9k�߃��)qQ���N����݅K
bW�h_��$���6G0N���)�UJi:ԎN͡ ��V^J�����*[���jtuה���!�������B�~mD�<�B<5j����Å�/WQ�oa�ᐷS��c�ȴ�����w����%����H��gRkpB��W? |�7k�9�p��,l��[z�V�O���id�D�D�'��Z���H�}B��礠�Sza9��Y�Eh��O� �­���%
��7N��
mۊ0`ow�^�u}��lT{�ꗅ`��q��w��Q��ˊj~G���َ�4UEF��pS��Հ}w@��J�`��'�'~w�E}��J�p^�Cͯ#C)��I8�=���n��5�{�x��ތ�5�B��$�v9��S^�5��1Ѡ�H���	�F�����|Tf��<=�g�xmf����qw��
�����8RV�G�0Ѱ�n�>y:��YƔɼ써%e��Lf� ��0g�'H�Ao}n�[�\�O1��(���:��%W����![�"?��m>.�!���C���8��b�Ձ��M����sX��AE��8f[y�Ә�/��XA�_�1�T 2x����[�#����̃Rt�M�of#Y�=�TELa�\��Gs�;��ʭp?��|��+�[�������B����}����N�����FC��NL=��Y��^��N��Aqu���q.-1�A�e�$�N
��I*�0��:�/}=�;���^��	���v�ƲN��H�Ŭ���[Oz�(�à�4�'���A8�(�~X]��숩��������8|��b�e
�����f��yW�d����4���W�_?͛+�˾c��{���gk���Ԍ��	�+�z͵�N��Fr�rh�iS��,l裮�ۛ�4�u�F������D�������2�C$����5����n[z"t%��k%:D��9ؤ0Ú���4�]�POP�$�n��Z\s�B�PcNe�n���.����|,Q0�4^T����Ha�NW-c���P<0�b�5��	*�l.���!�R.��7��j��]���C���:���krQU+2�A��*��]�r��?�Q��A�!à�H0�(	�\v�^ �b��E������a�&<��੏�8w�N�/s@���w�p: �뷼4�\S�k(c��`O���Q[��y�1���'��{ԝ��Y��P#��5��SYA8V�
�����#�Tx��3�!Ӛ�N�A~�̚`:5�Z���;� �z��pD}���%m �|�X����\��^2@�Ϧ�|�yi�� ی��qI�2П�����J�\��OF��<Ζ�=��/e�e/���7V����b��K�b�_B"'e�p�6�g��ɹN} t�4����=�<d%�((�dj�� @����� ��U���\�~��Er�}!vV�"ЅN�Un�G�^�5�f���e߾[:s5�,��}@ua9�S�A����� &8r��I5]k!�(TSH<T]��хe��i�S��A�Rˏ������M-�qd��4?��	vy�k6���o�B�_a?[(o�8���̚�QT@��^S��
��F�J<}��<�vm^V��4O�y�9�!�΢wx��Gpw@F�P�hQWJ�96)W�L��"�2��E�6��%_���9-R�Q=\b��{۔3)l-ln���?�a���_����&���|@̒X���P���|ʝ�m/z�D��mΛAB�$g�袺\�� ~��vB�!�i�����"�`�d����	�& :R'	-��w-1Z��%6'�iž1ψj]�ЦZ-���a��62m93+TE������Sl�N͍��'�2����zПL]�-�?��|�,��K�o����٤&�e��E��.6���0͐o��c�{�pCB��@�B%��TA2C`B cB����a�]����)�a�DgՅ�C�yR#t�n*/�Р��L���s����Ze/��I��³��LJ�?�+�ė����N���6�+Dm��1�}��C�y�ж�|F��V�͑|-
.@x���6������'�)�Hz�#%�#�l�ݻ�^����ʽ�{�C�#�c���7:0T^U�6�̥��(�4Kڅ�J2j�F5��hk{W���y��{��O�Y��~�0�����㺋�oYD0�ݲ'ƪ`��N?�LUH ��f���^Mr�cN��_�-G����-�����k���l�u� �_��@(dwd�@�`�d�]��%t�Q a��2�9�Qe("�*�|�k�B�B�XFk���g������J��҂+�X�e�
���Aq���RD`��������q�9K�r����=��6'&�&�4u��[0�����y��o�N�F�V���cX�'l���ܠ�c߸�a7����w2V;Q�I�X&+�������db�x�<7�,.an�`N��!ʑp��qw�c�i�u�]�Ô�k;�R�	���_r�}�_�������Y0�wM�5�ip8�Ng��F�`�-GY�N�gi�f��Q�2�3���{����b��J$E�|x"$������	���� ��;�&�:"�[�����Q�G�&�v��O|�ﶆ�v�(ـ���ۨE�zC�]��������7d���y3�Jiy�N��n�zԊw��dcwB����uH��~�A ;B:m���ܭa�ev����,W{�vU��o ���ve��z.����0N3 �W�?�#~�ѝ�S����X�� ^-"P/�wŤ^�
��ؽ ʚ��n74�O���[R�M�x�yUY�y���y�B+���dmf��I�,0)�N�,���A�@�MK��$<+����Fhy���<�x}��-��oqj~�>DɆ�6�C�y������}�:n�G���t���p�ּպ00gQ��Kܞhߠ�LrP������D���`��T����@��F=7iv#A���͌�38zoT�䶇A=V��N�{��3noG�MAc<J��b�DcW�G��k�AaJ�'�_O���|��^���>l��v�\�,��ӑ{��귽iԚ��r��/**@K�8+�@%���}t�L_�7�Nm�\�z"f��C� �D2���M�rfi��K%��,uE�ޏX(C�2�`7Ú&%��WNВ&)y-���|a�)�`7����3я�ݽ�<�q2�0Es[#jpG�(Q��C�KB�~tz��\���	L �S��V�LM7~��s��6eΌ�E`�Q@	*wViBo���>�M|�R��ܒ,��}�ϪTPDq �y<�	o�hm�獿+~�'���+p���Z��s����jo ���̋yrĤ�z/�U,�Y�%�gF�LW�\�E�+���i��O
[ͤ��w�-W�P��*��ջ�;��2�0��a��-�/��P��C�h~�n�i8�[YR����P��OPhH\X�G�i}�onm܈�"7��)�m����9���v.�I ���������Y�y|d���A�Uf�����c���o?�t^:0u�Z
�C�����s�i&ȃ��NӵA���E����B8?Gp��K4O1�K8$O'��_uw������`^���ǌ#aոQ��)R=��U7��
��uvl疒�@�GG/�S���O�+j����;�ս�Y��;W���f��	TpY�𣱷�����XW��� ߡ��@{7�ߩ�!�c%�|�ږ�5+HڙU�(���U9�<�V��I��KhN+����2>�u��	w�����k���S�-�e�t~�3�M:\��o���.=��\Х�`'n���v ���
��:�W⪐����;Ϙ�eg��iA�0��̄��^_)��Y��k;S3��=���`ZJ�(�$��1�!\.��ǧEkm�P!�;9;,�'�^e�L��%��,�SQ�[E����]���TP�I��]�%"��^Կ���v ���YY�FQ\����Љ��oWZ/٢,�E#p�����)�$5.*ǔ��S�=��Q��X ��L2?� ���m�v��� �p�>�e0�ͷr�4�#�3�q��~z���e�X��cV�L�a�tv�l�LE�,�_8Aʀ0t��2����
e�ݘ὚c7Oh��S<R����ga[���с9qס�J�\d�=���m�#���G@;�'Cu�4�A��31�ӱ=�H�^�,��F���tR��l됿DU(涛R���t�x=+۹��Ta�B� ��8����	�̍�i݉�����j�1��Efj��9P��̢�po�q�t�HL& �?���v���T$���Q/�.�q���6P�_���`�S�[霖,��1n!��N5�j�xk2T����HA6Kɲ�o�
��� �^�g�9J<u�42�V�=��/lK\�\�8}��Q�$x
��_��(7G*��j�%BƽS�ҭnK�7,1��2_�ZҐD��Y����۾0����?�U�8W����0	w��Ej� ����-	�5��7��#��nʿ�'1P�����Д�j�<���$/~Me���k�Q^g��J�O�����u��:U����ҳ �=-�&*��Pd w��Gd�C��)����Xs��2H"'l<ɚ�U��lɈP�q5'�#�8O��}� ��/}G�
XkqV�b�g�β8�Ml���L�CR�n��%_Μ''�v8�>cG��5�IXbi�M:�$�+m��A,TbP���#a�2f6�ݟ={3���.p��3؏�&�{Bղ�K:�2l���AS��J�Iy���y��p��b���]���J=X�Np�;������i<Wե�\k�T�D�C����"jҍ0�ι>J��G�mV��8�i��h��8j��Z�W�HҴ�8oq��j�!3+�n봎uBr��0�ij:O���J�2�?f:��SE�߼�z"ߋ��8�@/0���@ c�v{	��0 0>*0j�����0���L�G���(��?Y��T<�ϴO:��ekm�@�)�4�ź�%�z�B�b�Kݝx�}�V�H+H=4�(�T|���<\[Y�қ�+�Q^�9���n�*[�vS��J�R�z���o5bgsk��JB�񇌬#�i՘�T�nQޝd�W �V�鑗�cR����В�L=�
��ek�d~��>XY�l�6gɽH�Ms5��o���+7��L�ܲ^K̯GJI&l�S��~"�B���*���c�do��eJxv�8r�2� ��Iz&gD�,	㖿؝Є��;,W��J9���H���.�:CF/��
�
�>
�����;���Zd��C^�Bi#�a��Tڪ�JK6p;T��	���P��
GBZʓuf��>
���Km�/�}�@#M��k�2<1Ѐ{=9X�Ԕ���P��\�/7�W	#n�<xԎ�p�q`B*cv�Ŕ]'(oْ�MAp��V@������y��"e��T���$�'��Ѓi��Vȓ��ū+'DNT�ж�6����{"��5jt��cC�X��-JUc���q��\�����2w:D��������Q��[�%,LB���ܖԀ�ndBj�6��çzPm �����C�/�Dˏ}�ZXґyoN̐�0ѿ^O��J�������Z���c�����l�C��m��Q���LԨA�"�ϊz	k��F��L�䏿Kd�W�����CY1n�f#�F�����e��3[�`�A,Y}���=9iRs���		�:��$*��5���ġ�����>�@?�$�%̯�5X�&����C�t:�������` >����#�S��9�y���8X�8����sF�P��9�}@GI��<�ׄ��F �X�˗ 旳�ï2C�O����Kf���^xs9�sο���yԘQ\3|��Q#�2��<K�tu��K�:�` w��\���,���JSٷ���#0jX��C���c?�G�T��g1���V�w-2�.�Dq�f�y1;b#02o��>$n�iJep��X���=�;� ���CO�'F76c��m�����h������&���Bn%�̦MDugP�ǔ&��}?�������ߏ#�~DkΌ�%ź�s(G	⃠D٤��g�-`��cp7B%��|�*�1Hd��Qo��
a]���la�eq�=�}\���N�����}�o&��̤s)6K�Q �jk��T��X���Y"�}��8$Zv�̇.	0����F�N����(�w�q��Oe�N�Y1!"���2M��TK�������c�@YJWø�W���AD99U�O���������2�͓�]x����8>�ai��!��P"b���O{8�BF�xjS�g}ǶU�P�V��  �zvT�n�Cwz@���>�y��~����u�xW���˄��/�;��,L�ˢ��'�����P�WP�̲=����/�ɑw���z:����a-;n;Re��393��6��Sw��
�i�Ho����)�sJn�d�a��d-d�x�`�xz����a�"���j7\�$�w~�����U<����	��{�XϢ�dR	M_ʢ��EX�ʼ1ը�itG��z��l��r��R�q�"O�M��Zf�}�
!t��\�6����2��/%4�4�>Aǣ�� ��3��~�D��N��?$ˁzN�R�|����ɥ��,P��/�9� ;��?��v�#�΍��'a�!A�7��s�}�����Pˋ;֖ ������Gp �1<@�i锬��ts��x蘯9��V�Ƈq��/�٠��eB�����Y�H�/��w�W��Rx0B<���]�φ�6�O�^\�6D0\\5.N:�5χ��7l2a4ʻ6k ��(�Na�2ATD��U�C�p.}u�E�P�c���^�:�4���#3���k��,+�q@.u�B�*g�\��;�y6}�<c"t|�ʩ��kl�
&U�:x5����:"����,�L^�>`��O�O{,:9����\�Ӭ�K�f	O/G�~>�L�pw2G��7\�o�^�<,'"�k��tR��Z儿��7��=%N*�^�������H�������c�8-T�t�R��":��َgC�x&� ��f�2c��N����xj�/�ǘ7���︽�R���s�E
w��B9k��iU셽��ѯ�-	OEq,���T�뛑%��#�YG��Z����HcQ�Q.>y��IY{&/� ��= �eƎ� �n�O'��\Y�P3�quH2�]Ƥ� �.F�#"���H�0T��u�=��^��P<���XMv��[Θjs����:���KiL~���v�W|��X���)��l�zԊT��G�gA�Y�b>U�7���
�n��UO�I����MXx
$��=�"�9f%�7�2����S�}�v'�+ 3��#�p����X��C_���s�G��u��I$\�h9��"�C�⊿�����ǆ�=&����W��}�cWȼټ��)2�i����;�:.E�!Kd*m2��m0䛾�Z��>�0	+2}ۖr��m�L
i�B�����������*-�l��3e���o�0��|k�@������+eBY\(���l�� ٧����AA�7�v�}Y���S���Ϟ�(�D�-�9o2\T���ۗ�|{�D�L�>�F�O�uC]m���t�9㼥���~^��k�;�K�;�.0?���9#�[���c�"�,)�Z��=�(�v��\v-ˊG�����Xwe�-�_��.�xEqM�=ϔ�r\���4��^ř:C~��f!;��ո7�!��D�B0��"�� ���.<�y�{�3�ѐ�gF�1$�(/����z��3ނ�amM �m������S��9�Se�����@����>���f�q}|d=�շ�6g͖��}�RU/����b~7��vT��uc���s�~�	��}$Q��4u�EU��Z���V<HE�ld�����_#qi9�S��ԯ[�>�w����|����?�pwpgY5�3̘�n\)�zb���(fP��3a)j�I��~�rV����6f�0���䛹g���K�<�=r���;ۘ#i�Z���]b
Ke������d2"��0�Z3��NZ��uM׮���i�������'�C�_ERg�77@�J����R���3�J�G�8�t��1<�S,G ���߱�sT'�7�|��-H�`{���}����c@��p3�щ!�Q��7ԔG!�p�u8���UjT���F�y0Xa���oZ��E�#���H���_h�}q㉓e���=z1y������Ҳ>�V���r�`�y��11�ʨ# nA^K@\D�����}8C�ʺlJa�dΎ�.�k��	��:�������7ߘ��,s7�Xy�O�2	��"�6�&+��Ȑ��\�Y�:߷Y�ג�8�<��gI��v>^%���B뻹6_��BdQ����"z{�t����Tt3�G��<��W������-x���|��6�xxtL;J:f�-n��Zn��a�B��qT�����&c� ~�,T^"�73� ����?:1���~S �5��J}B����Z'~3��O�s����3��]]�EH�G�vc�˂�!�Xc	S�8�?�kR+���"���*4��j���s�k��#��in�Yo��l��o�.����R_@��%�5|Y�_����ޕ��0��H0�9�V�)�8�<.�G���u5�ߪj]������y��%��8��bz����T�����;s+$R�"�օ��Ss��f�Zl�?���P����QOS��Ǩ�Z��l�d;ȩȉ�5��2���B{RsD��Wt)9�>��vrq�)ܵ��GI3ӓY6f�V,�W�fV9k��E�xϲ�T����V{���c!�Q�9! r5�p�j�r�{)��pT"�E��>�󐽼L7��"D�e�zc���);w�9;`Ђ���~/�V^�����v�J	���\�w-BՅݭ̺%����y)�P��+��� ��S+�Ϝ��D�|�p�D>)M�5B��q����H�4���{���5l��Ս���61X��b�Y���',;�A
�! �S��Yp ����q,
�M��� XV:Q�2�Mz��Z��-�Oh4,���$��	����D�Ssg/�6��Z?x�g�0�˞�	ݔ��{�`�yS�΂`_�7A�f{0K�*�j��&z�F��q����$�<��8�gg�C����q�:�Ǉ�y�$�N	7y�xJNz;�����\F�����Kd��W�\��������A�d�p^Q �'�3���RO���&Ջ˹N��(/�̠.��g�m���p���]d:�^u0���3�3e�xb:�#~-�K�OB�C<������J��r1�j��V��i��5���xi�ٛ�X:�$�vK�����۶<�=��z_S'�&0}<���v�, W3���/!�3��2�>�V${ Ȕ����y�M<xc����y钗�7mtg4QFdVB���B	^2�EY���{|,Sz'!o����|m�͗��p���1���x�^O��	J���g41eU2qI���f�z�B��ho��|��l�{��򘣦�BfFYQ�q�r�<]�ˀ���=.`/Q�e<�1�&fޙs����A�Vح�����h��vJ�vD�z��b1�j� ��r�9Sv�����H�C�w�=����B�o�06��KASԢ�x��!>���\���JP��Զ�[ɣ�_�7K��k��-oc�}�X �`���Th�o����-�֦�!'��XZd��p�,�S��T �� %o'��-�!��a�v?��fLG1���j��Tِ�	��"�.d�bɗM�gI(-D*�o%7��n���p��p?�Z��g�*(�k��"��n����t�A1>~_g��J+)bS��6��QS�����4J.X�ܯA��j%��i�ņ�kNN6�ɥ�G���׶"�����g;�u���]`$(�W�A'{J1�3P'�{)dW>��ҞnjנeY��1-�X6&`3����{p|=�T��wz��	

L ���S�?�py��K����:�B� ;Ɋ&{,�9פּ�c�KQO����=C�~ٓ����0('R�~�Z���I���x����gz]�.y!�B͋i���8o�.���^|(F͔nݙY�fgt�P��`�"C9&�P/!�ז��"�aJcy_���a!���0^�\p����rP��G:L����+��wf؁��v:���Yf��7؏��n���bx��f�����)�� �%�b����,U2\|9TI��u,*I��jt�2��^dُ��Ӧ���ȴ�*O\����o�M.�J��~2c;�h���� ǃ~�G<A�F�h��b���G�Y�69f+Mθ�Q8���*���ǊP�O�S9?(�G\��,�'�՟����¯�G�y2\E�KߨN��	Ā�,}TXق�)�y%��ے��^�@*�����jVA�ߟ�2���a^qJ��Q�W�P��D�f�,�(bߖ���t�.E�Xw��Ĥ�
��k��.��EA�j��{g�t;8�?�4B3��N3A���%>����3n�~�m����(z�������}l��x�pS�����!�\X)@D.�[(�A�O�\)M�ϲs���G�V���bK�̤+�b��e��>+��İ�����=)�xVxnc�����'ۍ��Uz��/��_EF��r�Ũ�q�uQ~�Cre���R�6V���rL`��ܷ����w��#�fe�.�g�!B&ȾQx���ȇa���u��>�t���0PuK��s�de^���}�[w�I4��<M������*N�{^�f����f�r�g.RL�6��4j���'��v��֊R+��b�ר�
� � �֕?�k�;I*g��3҅#��W*,VvO�gK+}yR�[�,�~�Rw�R{=��d&q@�YS��e��?Gh�K]�����7#���r��$wQ�e\(�M�����J�K}x��
�u�q���;tM̳5/g�`"���F���(��C.O5'�a��u5�3l�:_,��j���0���2K�{� �H��	/j��Jk8�_z�c\���|�~�R,�jys�0�f�lv� �,XCUl3R�0�S��R����×�-��3ޗV�;�����E�p��	����Bx�.#� +����;:M�RG�������i���k�gF���r%e��3�\d� ���)��$k��k��p�l��ů��)g�G���r����U7�]q <E�%�:����?3at�j	�%�զ�ِ{���#"��}*�h�lJ�oCKt
�/k'��
I��EQ���H!k�zԯ��@��b�GMT����@��"�C#�8����x.>�BV7��*ti_l����ug$'n@؜5�0�h��B��̼�,���5��8��+�0^����&X�����UK����螔Q�7*`15���=̆@-E��B&ݯ҆RE�9h����ͣ�����9���!����<��_7�0�	Q�Ws�9��|��� �Ŷ4㳬(�`%�W�Ǧ{neu��D`vR|���:�dQ�I���_P -oK�\Y��pJ� �C�Tb3�@��z ���^�9Gn��~t:̞��D]BUm��2���A�T�B��FGp�PZ�>��	T��c��Dx�3����[�#8Dv~��&��OǴ���@&qqL�U!�Я?���O���&�,7��D�L�J�3�PzJ�z���ֵ�I��bf*�=�$� "������zĜl�d�ր�y��`9��-�������k1А�v��=������A�����{g\=�\�"�!#.�/=�_�[&�,@z���yl)�#��Y}S�`q��C��Y�B0��F�
h��M��0��"([��KL�H�L��,L՞C��{�փy��6�����ټ����V��X|�zc����6�@�� �kt��Q <{�XG&R_�K����!b�����<��l�7�E�Q�U�o�'n����&��A���NjvS=J@���z�8��Az/6�(��b��c�0R�A�e0���nr���J<x�*��'[\�(ت�x�}ȋ2m�R����Hu��r2�d�Ec����d�~����>)��1��I��&hŸ��Z� W�4����!EidT�"rG�jI��������6�C�]zSǨ�/���kX�P|��Xv�r���0Z);b�&���%kղ5"�s����%���W���F����(�\��8LQ�i�,Q�"�KAL\�;�W�P��©��r$��k�QfF��-��Y�����Ӎ���'�+�8.�Kʇ�Ʃ���͡%|�vEm�\���٧�����Gw̱�}�*|��L��a��2]<�P�ygsz�V�`	qO��$OY�gM���iTܝ��-?��<'��"m��ڋ;-Fλ'.�;��Ș��T0��Si�~���ز���TQ�����q��OŌX�$u��]�A���(8mܮ�D�ʕL]�^��xK���z順�f�P4�'~�e��<WK�;;)C��АQ9� �a���R�C�.7ޥ�br�	��{�N��
2P(C(
�6W��)U�������q�֖��M��^�"aC�Q7H2����
�z�鼺^�����i6/Ҷ���"˛���kk��,��B3�Ȓg�T��dC�u���r8�O���՞�l����G��m��LN���u����{��e��V���qki�$'.Cج�� ���x��k����z~�4�ԕ��s��g؄���zC@����*���f������X�, c+��3��u�V�����$�����U�%���Ӌ�f*��fe(����B���g~:\�������w72z�EhxK�X��70 �&�Y��ڃB�A���GT���]i�'�J�2s���~�-UF���bL7�2$��R	��1����k�ߓ9����>�|�J�wvJ�SC�F�ڌ�ل��k�	�E�o�"K������2pz�-�f�1����
(�-`�T�Җ.D`訌e�Kq���GH�v߈ұ�mA/\�4�p���蝅�2�A�;�rh�E����l��\4D�9'U��Y���V����e��"���xTRuO�~�7��_ٗ�[���������5��q{�����c���(oGî�\� �����)(�37�D1�p�Ţ���.&�z檥�ih��2,�����p1�� �/`$C�Yh3���_:(��9���C�"tX�*��JH�C�����"'NS=��G�<�2���`S�J��b�?Μ�|D���i��1��M�Qq������$�P�
�`G�w1���I�����K�����PWs�8�ldY;\�fÙhL�$�$�-�0:�~�6��u�NO�:i�A�Y��BxP�7rfQ�	�q���伶��9-�;Ӛ�"���nT����@ ��l��R���ݐge����9�K#�$A�u�]B��:���2�w��%\�c%�f���E����w =D���7��S&�Lq�y��p*�<nyÅ[��S��KД�� _��f��\_�Ǒ����;@��n�CY�ǘ� �Y|*o�y��k���=�
ދ9���t�
=Z>Y�)U5����J�`χޢ�:���Rû&��l�xt%��43J�\�hY�-�$�<�O����;ି�E	����Ah d��67tnN ~?vz�E������X~�X���Q���
������H�V)$�5�[�/JS�̋�	����	2������(�x��փ�U#j�RD�wn��Z��r�Ω%@��N��D���z��e&��".EQ�~�(���/��]:�}��Ѿ�s����r��/�$����[��4��.���[�H%���ZzK@�&�RǄm/��C��(^ �("�a	b�{
>�,��L
J�%�:���4[d
�\��V4;X��;�C�k ���a���Ltm����?d������b[�F%	'����n���^�����
#�jI� :4[�?p+w�S�G@���5���HC��{�������S�J�48��
'��D������:��h��E��8&�!o�k���h��`L�7�2��#��I��_�*mUcO���"��W���� ��&O�M�&jmT�"�(]�`I��l����s��zݳQ�s%g�Nm��K-1�|}J"7[w���Zx?�Ѹb>�)�&v2�{À3r���|Y�U��(]�˫iϾ�>B����-'�����ǹ�U��ŷ|�I��{��`�}TM�K��ͥo�<��jjH_�8�d9��:�N�C�e8\\������ο�_4��}��!":��N����:%s>V���f��=�mwG�18�P�}}�Ƀ;����/� i7d�� ��8�/����M?��}Zf\2@�a���2�~n�J��d'��h7�������Yĉ�s������z�% VO�"���Ai=��?���# C�J�y|��`#Ң��"�O35�����90�r��Ϝ7��늜 ��_L�n������ȳK�d�Sן����|:��^�cg��d�鲳��mm���5�C�l���-j=ɔdP�A���(_�G�N���X40?A�j��:{]/��o��Ę|��Е��Fb�X�z�5�?BY �i��~��HZ�[0�%��!i*$G�ko1�n`-4�r£���"^6:�I|9f5De� �0'���o5�p�{j�ʈ�X�K�TnrM�:�����ۛ��� Z��v�������8X�to��Z����F�Y�pw%�xMU�Tv�&!}�ۖ�G�Z�)�ɩY�vy��y�Ȣ����5�F�c�|V��,zl~@��%�����o>�:7��츐Oe�e�� �Pܑ�I�v�A�����e6g��	&�ڶWn����rJf������-���W�!���¢���d�%?����w�_��I	N���x����Sp@Xr&�p���2&"r�WN+i�t��pN\I��S��"�b��p�d� p�U�3{��~?��t��ՠ�ќ3���^��G�A>8����E0]�|YT(�Y�5^˿�MT�,^�r�
��/��zʱ�Ǐ�zz��cz�]���,/���Wi�&j���o$ܰWy�go��/�J���Ѭw~>ݐ�^�������N��7[�ʦ�l	�p:�,p�����7��Cs��x�sG�Ԥ��E�Q�"�A#;ZB0�f���94��� �d���j�B��'L�����
.�A�
)��_#cB�����D��_r@�}�m)uDtv;���Z��O�����X^�$���H^.j�{u��^;��Ū�.���y2{�K�Q��hR��U�s�����pϬ��V£�ҮB�NR%*�=�4^��0BAl�eT��[����)�0Cv�;Qާ�%�L~��̃n]7���r)k��P�^��<T����ܙ���PW ]
-���!�����=\�_<� 7P8��*���ezQkF:�m��`��А*E�b[�?˫u�Hr�ҐЋ_U|^�L%���g<�5P��8��<k8��>#�x���̍��I���B�T�i��*��^	GH鎺�fC��-�7N�蚍Z��* �aQ%YrF>� �a@5�nlE��-\P���� �&@�J,����7��L�sK�}�\�>�-d���ϑg꟒�c)�6��V�jܷ:�|hNQJ�JP	�-�|�S�v�^��� VV챨�K�9�����ʝՍaO^�ŷ��r�!Z�+��"-t�.l0���q��o.|����~#1�GW�ޤ�,�;�����L��;�qi��{g���	�nS�;��Q�ˆ-�4M��h)Շқ���S*��B��㡋\n6���y;ov�������3n�����Z���.�ķ��J�8�Ii'��4o;:۵9/^/�-b�3\�Q�|'������]X�������A�U����8a�N����єAHb�q>!=����0�)�b3tqDg�*�m3ٱ�b7���U�(ĵ�Zߧ'�+������$�����t��B6Ll<��T��+�+%'�3��##�_B��v��o֯ɯy�UMē=b	N2	�PJ�y���D#�����N���B!���}t�	��4���!t��x�C�#���)g{Vb���o ��Z7ڌ.�.c��qc�����&դ�~Mݧ��S�6�p���D��o����E:�6N���W�
ƚ�V��64!7F�/p�(�j�	|q*�Z$Ŭ���s�i�F�H ��������ϋ酄��;�Y��N�$r�����i�~�obƩ4�IއEI!����@
��Ŝ�z�i��r1S����8��-jVċ�89��RX��x��Xq(��އZ���*�
8{P�, 5nɫ��3���_��1$��h��O[��d|�Of~M��U��>H�u����I��9�:G�wSbn�d����,��t�_�G*����gW��{]7Zt*)���Hc�f���SO6��+Xy�-��i>�����t'�G(Ց{����"kN�r,��BU�3��i�.��t�Wٱ��X����a���`��O	�I�U?!���@]�=H6��oRL����J��B�zr������!h���`):��<��
��!�\$���A���N4-���>wB����f��<t�d?d�-�DD��H�c!H��#K��ޖ62���_pnup�r(��쁂�@7"u�?	ڭ���a0N�B?s=+R��r�7����;�7s����B�\%xi�s��b��C���#Q�:xb#�:�|�� ������%�F�_����8���������LX�c��z�ĸXv�+�r7���	5��z�"�=8���:�RJ�B��Ξ�����3i|J�m�<ǸD<�^q�$fT/u�TX���5�yH�Q�Y�R��*L�.J�(Y�a�W�'�)9��pv�}��3Z�����ko�������4�&�D��dqB���3Q@�r��-���;,S��Gb6l�	H_�Pdh�83�&��
f�&��B���_\�K+�'��S.�n��M?7K+�Q<B�*#�O�_D����%��{�:�A���~ײ �+frx�\y�V2�@��2虥~`����N�=/#�=�1���j���b#�a(����4�JA�f�?�����v�����
�bH�_<��Z���If�%4��,��[�T�5���ݭ�e���#޾��Ԣ�C���1�5��*Z�)3�93b\hL�i?1U]%5�����-Pgҋ��\��xb�c�)$s�O`S�R,ᡥzE�F�d��:�j�tRjO�t�C�����f9c�\��h��f���$U6'E�0]p)E�a�=ݤ6\CU�O�l�%wϱ���g2�:�\��P��O_��	�ܮ��6M����+?��`��	C)çtm��n
9��g��5�kס��/>W������R�Q�c;���'1�����O�ژ���rn�퉫�%@C"�
���>�*:�R�q^Cr��C��{���wi Ru��SX^�[^5e��Q[��Ey:�ܸ��
E~�,2p&J���Ur8��փ*�M��,ayS�D�r�LY�T��=�4��7_#�����-c��3~a6uǸIu�����$"�x�����e�L����G��A���������]b{;��ե��B�K0QI�FF�6�f�����ty��Es�cYZ��!Lt�.a�3)Gl��G�d�4w�}%�Ͳ֘!�Ri���i�T�� ��O����
.�K�m	 JI]JKK�@@�4���AH�dͿ�����ORw#��M�S����Kɕ�8�%����ˬ.SK�[�Hм(S�F�(o����S��qG�D���v��5�) �����	>*繺���� �&��HnW�՛%N�}Q�J��5��R�HxD�V��ӝٝ�8K%�=g�:���k��@h�uZ���b����xk��J���gj� �R�Zj�Vϵ���z[*�b.a�;�"�`��+-�P7���J!Ҧ�H����xGa�Q�sN�k�MK�л���V�zmز�<1U(0\�Vpydb�wT�p<uh:��f��ս݉8���k"j� [
������ʟ6L�9X����`�_Ș���(��=ͨ[�;}+�~�)�����إf���p�%IٮR�'��j��e��i'>�;:��� ��o�)�ϟƉ���r�F���6'����yE��N�A~i=�>�	��FB���l�������4z����K�K.��sk��(�\�r!�`�E;I�����8���+���L����7 �`��\�̽�)�ڢiğ����ى�J=ي����0��Wqv"��1ߞDK>S���I��d����õ�M�`���Q/Ԛ�;dЫ�wf������x�)/_���N��yq�����s���3A�G����.W�ZZ����fL��m+%[|rG�ҩܑA�bJLc�Mepޟ�s�غi��l��є��e��r-�\w ��Y�V�%"m���0ZsG��C3?����VIK�$��­Qe#Ru���N��+�$AG�!Bx�"N��;�+�06? ��>@�DGb�
����9�^oӊ�1<�-V�������e)x��e5��b��#8��4]��hf��gͯ9�EkIrH�~s�_
��Cd���M ޲BX��W��&��^xr��ɬ�@b��֨�2���]��_�����@/:�mϽl���^1�â�����܅
�Iy��o,"f�f�}� j�v/�+j=�@�����]�D����I�P?Q�{�����O_�
����� �v���y��I��o���W�֧��F�(G���䉗�d.׬��+��>��].�T�d���j��N���= EMb^	����k!=."@���	�k�ZƒJ|�&�ʩڋ%�dК
yk���BE�8|�bI�A�m��>�32_%C{f5;��� !m3[�lB7�<-Q�ܮ�[}2��(i����G����"��}�2��hh�Rܐq�&��_�]���[�������Cj�u����ؗ]�]I��ʲV(�։�v��%O#p�2e/u{�؝$��Z��X�H�É��K0��G��}��a���c�=Zlg��\��H.��6�� ���8g�}�ԍI�<e�6^A��\J
e��������U*��>�a�o7��拰�k��ֳ���-?��y{�c���߶ڱş/�xS�ד���./J�~��N=:t��Y'��l����9�b��UEE2^��W�j�'��{5�ۿ���*��;��� ��x�j)c$����s�񀈔����W:Ji�AO6/��|b�Q�>�⨙
�h-�G�� �1��6�� �n׵]N������a��2J<�#+Һ��,L���A�q�lJS�5���-|f\1���O]f�����C��n@�C�Q0v�P���}XL�_���}�~y��34X�wC��W5;�D��LC��p
�g�P�?�9F�q+��^pW+���C�k�qM �rUoJ�����R�����nZ`��3v����u��;u��e�c�@����Tܿ�͉�8���F�Ow8�$5������A��\<��v�~�w����^F��(6��h����8m����d�FYѠ��� �%�n>�l�&ܿ�^g��`f�Ŷ4L�t��BDH��3T����	ɴ�xtt�UЌMס�-WA(�9�� /dJ��A�IQ~F�aq�嘶�7 i�1n��\�~PG	<E��O�2?�b	S���bw��I�k�=�@��o���+j�u�p����	��֎����}m>���^��׵6�|h�A�S ���+����_�S\��̗�}(��68�\3؂&0`x�W
>c]iB?C^�-�*��\v��N9�:�6�f��}��o�0e@]��i���gd|k�ΙzM(������O���t�vt�g/$�b��%���L���Z< ��{_�ks����B�g�Ƶl�7i:YcϷ�CͣXT�hm/�i%���׺�9�7q��12�@���ɹ(�;VJ�pҭ���'�b�z�BϷ��IME��T�ӂ��K���.]�����F��>le#1���S��4�Y�R%�oM9�:�$nhy��b$�5�7�ڄ��ǝ/�#�%�a�]��0���'oD��i�t���(��LL>���y�1>YY���^d�	K�;��y3l#͜�*M��<��KhM=V���J�
r�(OB|��\'���5�)��p'����_�l�;-Y	���s��n���\��(�g�X�b�c<�.齑ܧ�����C��M��� �Z[�@��2��cHC� �Y'Yl�B�
��BiG�z"�d>�~�&9\^1~�Td��� kV����Ϧ���! e��?�=��JW��^�\�:Y�����t/�ל)I �nL3*�:����᭽���P�%9U�� o�.c�����J'�5�/ς!ھ�O*�?��?��?��&��5�n(+�v����l���gBy
�����[�8�up��i�������#��l�O�;�2��j�>�P�^�!�d���z�=u��؎j1B�L�PUgl�������~U��~�([�P�Se�/˙f�YI��ʴ]l���������4̳�jʤd�ό�#"�A^�y{�����B�8^��B�ٝ��΢//W�����Z�-w�9�9yE�u�� ��g�2�c|�}�]4ʮ���Ч��}ɭy{`��wG�>�����e�|,H����<����@�h"�g��ꄹ���K��	z�!�Sw��-��x�������qm�ȓ��XX��r=���,��sl��ne!��2�K��
�"�����ʃ=���+u�$�Wx9���>�do�M|�{���w�:�݉6�����+�d�P�.s�?t���J�%rKHL�y���%�r%�-$�i%މ���/n��-c������& �"Dhk�qרM� .K8��&�Ml�H�����ᑚ]Z��@�}�����(��q-�uo�IQ�,,"�M�}�S'�}�pl/!I�n��@�Q��17M�d�����Y9(��ko������ty�;��?�$�}��Ln�~�(��oz3ժ�%�Z+B�e�2gt��~�
� ^Z����	ǅ�h�\4U#��I�3A�=$#��(�����JzjǬbn����BH |����J(�sRm}�4�S��sA/�p����R�_T\��?N�JԡN^*a �o��f�Y%���p��F�b�o4Q��T�v�ȍ
��Q���m��d��7�]_ʫ ����AS2��.������G;�8���lK�tR~� 
>�(߶�8L��4���?��O�F%�� LC�(��}��p֛肃^
C4���}z�F������єAA��Yע$�N�X8Ȧ��ӗf ���hP�ϩ)M��ݺ��fn��5�{#t�D����^��j�`�.y�u߬9�����N"�Y������b]ר~F���_C\�pS�n�K��ί�.`�c��}u�b�0�U�ϯ�G���v����%����_O�EkGQ W�o���ϰ�A I�a.���3�� ^�Ϸ�?�3Wf����:�Z�S<b���$'2�xo��?I1�}���d��/��Z��Dc�)�k���s�$�Li�*�D���-o��+3�^�u|٤����rgI[�/�J�Ì�^�R��Rp���Z��qy�x�fySZ߉�H�Gp�.�ݤ���)�[��Z47f'��������c���>Q��u��(U8�-��+�y�,���.�iY ��"m�x��CF|� �ԘK�X:�`dxB���5�CW������a�1�� �;X��<�$V(Nc0�/�{e��W�x?��حāZgt�-�.��Dae�����)]l �,�gj+7s����o8�<�U�P�j���[�������4�ɤ��k^6Ic������O3�\A�0BJ�wN�B���gf�URަ�Ѻ����P������~L���]��F�u-�����gW弤��3�T�Yg�F��;���q  �4�{OfXλ�W������ih��/�K�������N-#\HG���(�h�����`=�P�[���ǻ����0���l�问��/�P#1ݘ7��^�	6���t�i��~�t���4��Ь�<.��f`��&�2�S/@�{�:�_ϒJ<2 4s�{���I2�O�Yִ��y#nͭ��b"��<u�S'�Ĳ�sG��#��Q��=��E�`�I�LV���b=|G��*#!ۼT)��2�����L�>��K��t��a��(MBv@f�h�^_�H����:{	�
`V�:�;�.�e��6�v����z}jg&�E���?��f-����!�ש@F?K�5:9J�f>@�r���F�3����e� � ����'s�iE������4v�,�;�(>�]d�{H����;���L���~�%	��@n.\�m�ig���{S���E��㎼�	B��ѵU�h^��9i54>�[w��=��IW��|��=�����>
~-��s�ip�mpױ�=MbP��/�yA��Y���]�g	��'	��S�:�v&n�q6�^�}��a���ZD�?�@z���l����"D4sY�pqqH[���/�N�h҅�m$Dr�1���B��\mT)���t�)E2[�����_m��W3I�Z7�5}5�P�/�·�5M�D�����fU���=�To�ǁ�z��@��U�_6_����.6�9��ga V-9�f-�3�X��W��o>���\� ���(�=���z�<�����T��$�G
�	kS6y7(5�?5B�}9L�v����_9,��臭��^�1 0�/��BGfs�l� ��wWǘ"���?��t�3W؃���O��y��	��ު�v���ZG/��	OJ�Y<�B]F=��R�����u��E��ȅ%�>;�xf�a��c�T��pj�0���uKگ���˯j����=̗�(���Hu5�7S@�ntk:��.�0U�l�e��T�����9X�2V�w�
G�����QɄNy��-3NӠ��M/��.o��_2�ٖ:s���^��^�*��6m��~�E�
�ǫQք�3b	� ��"��2�jA`[J��"�"�)Y��Tz��r�x�� �b�m�6-`Ә��D�=�-���Cl��|z\���8��SJ�!?��k�KCl�9�������O#Xv��g��^�9[�E����$�1h;ښ�zu+z�Xoʲb
���f���=�� �)Ey�z��k#��%������b��[�!���{f��
C1E�k��SN�>B�J�ON��ps��X]rK.�x�.P��s���m�J�>P8!z)�U���`�g�r��D�v	W	�A����6_���&��~�%wH�W�
E^���4@&g)���8����/I�B�_�^�k)^��'�A��:��"q�[5�C[�㎘�Xce.�7����9�2�4.�E�����u"�vS��ϧA%����0�)f{]c%�R�������*@J	F:�[��2Z�s(���k!��wS��Ҝ�����+
�-��΁��9¦��8��\�$�_v
Tٌn�ħ͂����輶��+�`���Zs-���D���ϭoF|i��^J��l��#�j��+�$��D�ğ��M���l�a�0WX�
�瀅"�u�%�]{�w$��J�P���i���9��w< ���!�q�ʳ�~��S{��0��y�HξU�E%O�"�m�6j�h0�F	8�1f����!i@fV$Ro�8��k��r ns�����gu���>��#�8�~�^Ѳ���nBE�V:n��4�d�+ɈH�(f�����]U��M�w##ϡ�n�5YOV�QdȵJ?����_�zK�d_���c�X¸Y��������vX��}�n1G����C?�3M�Z��� m�T�=>�EY�����͈.��!דؒh%Y��l;��mad����/:�0�(��Nۤ���g��daRt�Y+!z�e�j��!3���$�LG�g4�M��w�n�ϻ�:5��FR�|S<���E�0��7���)��i��FM��¬�ت��oNf(�\�Ѻ#���e��!����"/�p�)�gꡢ��K����}Yѓ>{�>�� \Hr�̶�Hpp�Rn[�<�󴐲�;�yX���w+��.�$�"�T�N�|���'&˻N���)6�%�f�5���푊�P0c ®����D��XV/9��>�UJ6��5������
2�&��̘�X����6���+y^怜8�������E2gk��珻n/�0mQS.'ܫS�&j*w�	6b_�f���v�p�D�3�e��o#�8�
��ޓ��륬��r�v^&ޝ&��"��c�<���F��![AN�h�*��PX���\QZ��R���4 ��{Ty��_w}8
���O�5��+��D?
d��y���ɔ�5I ��_s�ɴy�'P��ih�D�O��r�����m#8YE�{�	�7��Zg�H9�'$S��h�.`W�Ӏ.��������يXQU�$߷����%�L�RS!��th�����b6@B������U���0�q.���{/(�L�'Y'{٣=wG���3���"�a�O�@]��oQ5<0�t�?EN�M� ���D�P�5�R�*�O�i����
�,@'��A���^8	H:ez��,=}�p�ﮭE�m#,�6�"Bj��)��/ey�G�O��A�#Jw8��#%X���7��R;����� հ9�ʧ��bOzr\����F��m�Nt3PW1���u��m�G. u1�c1YX�~`b����-�����=l��߀W��;��Uq�<E.����-`�N_�\K5�m�Q�]�[Ώ��9q)\h�\v2I�WEy�6����t��L��w,qJ��*�e���z����)Oaba8�e2�\R�6�c�GR��ޫw��wKc�+*� QgÖH��n)ON� �����Y�_W��
o���������_�#>��"��@1�M�!�6�~W��.��}�	#���ʚ�� ����AO��$b���ܶ1���~oV�a��*��uMh��'9;(��F���eƨ!7�*�a��o/r����=���+��k/(�޷e���A*��#��!�⣇�e?K��߯����*ʹ8��Dnb�&�Ңz���L�4_�p�(�G`\�T�o=���I.�D*�aվ_Ԓ��U�����{���k�~�~��!���������[?����W�Ȃ|O��r�7�I5GH�7m�-q�N1�Ct
�z�o�~�iD�  �}H��Ɉ�`>���"˨Fy�
3����C�x��
b�!� �xr�L|6~�k��������ׂ^I��!�p��w)؞,P5���8,w�������.,4 ���H������IL�-z�[0�`[v��0�2vjo��Ce�5�c��+#'�p�'�Ok����9�+�� �^���9Bs��ݑ�E?��2��P���P�ð�R���&p�2N�sPS�����?�!�)к��Vq{Iՠ=&����)��t�?	pg���ip���%��<�ih�.^�n�����k��s�4tVp�0QrO�L9{��>�x��aSi����X�W(?np���\��xe�f`���u����7��x��F*W��w'���������Y��y/jD=Y�2|�[�[����^�O�>`"7 է�(��t�i��-��Xa�8)6;�&�L@1Xu���0�n�=i�1�}���]�k�u9���F�6���	@��u����pq;9������ay�~�p��i�k�W����픧Rf���������t�uX �C�6{B3��U ݮfKdw��T����+�����5e#���vXvo�̫�)ȍxA��~N�MM�M�r�t����%�M+>��HT)-��5*6Ć�o���#H�-՗��93sI�H������R������@�4���̨��+�����>;�n�H%J���R詫�QF������p�K��}�%m�']j�C�/t�TJ�"Rlȡ�c�������3j��,^k�|9�w;(i�$15�:��7*�pÅ��X)� ?�ٍ`\���}��z�Y�&��y��S�� ץ+ 	8��y�Ӆ˼�F�a��1w�},ۮ(5�듅#��ʞYb���	vh�'����w�`EW�'���#�;g�;7�@|�"�XM�x�� Ebp�t�^�*W@"�]�7�ĜL�BP����7a2>^�	s�3�B�B��S��Yj�rl�:95>S~B���G[K�U=$���sE�њ��	n�l��Zn%��Z�Z6���+�ײ
9��а�}8��|��osK���G��,	�����S�)=�����n|���x�k����]V� �$�5�5>Qc�87�T��F�:ii)�!��|�o!�䖐� V�7q��� c��|�6�T���Q��4ޤL�E��)���rXs���X*�� '{��������뾩'ּ�Z!C��4">4v{Û���=��}��y��-7����;%,Jg�ͬ4'J�3���3*�ogn�z�^V4�履X��-�#����P�O���g��n�ɧΥr�̨kN�E݄����qD�c�Yz���bk��g�d������w�;<%-����0jU 
4�]ѿ�ئ��C������w��Juԟ-L��b�r���m ��'���;xP0[����ҕf�<֢���8����Pi�ّ�S;�y��ܕ��&�*��;.���{�LVM�'EIq)���{�����L�X�; �;Hι~H��\O��7|��f��.�Q�p�����`W��g �e���=7^��s�V��NxQ�/�L/�c^U��w{ϬM������(n)���S�V����U�ߎ cXXW��/4�p�G���@���e_�=I!T� ��erm@��55�H�Ξ����pߣp�*�yw(�g��>������]¯KSb3���WM��'�X�姄���]�I_ |&a�	�g�ͼ��`�y E���I���2�a�zAN���B���>�YK�#�T�T�`�>:��5E;�LU.��C�>&�����r�3 �&�����e�q�5@�PU��V��v��'PI,�eAG���	�w��xK�G�6	�h<J}��z|��}��4*���{H�����R�'�2�����G��aֻ.�g�	�*F)�}��S�}�*ۇb�KA�:"���y����q��

٪[�G� ��M殍,��h�H:��bu] ���!F�~���ʵ!)�aJ�5�l�k(K�p�����ih�M��Ȭ"[�Z�P�'Z����"�T�_�b� :Gyb�(�9���Z�]±?�x4� H��{c^�lٱFT���A�_�F�9F@�9qM\zu����'�M/C�f[���������o1��ʽ�������:�2�pe��MARnG����q�S@)GI�%��q;�Z�s��/��~ǔ[�$������\e{k�W^�Q�Ш�-��L
eP���C�\h��H{��B9��4��:@-�n�;-�6��?��<���A�+U ��Ў�	��C��>=��RkXގJ��nKܻ��gv-$b�pV>k����.|�R�k�iE6L���(x�V��
e5�JD8c����4��~I�e��]��ro�kˁa�8�����T!kwܱ�g��#v9�9p�Q�7/�!��A`Me�<����4������g�'�_�}\ZA�W/����R�v���ä�Z-��l}q�����Є��U+
� G�˴��9��?;t/E��މ��k�F=����q���������a�F�{T�G�I@
����\�pJ��RJl��p.K���L�:��6��e�z�7�X���lK1�ܠ�/��`�I �-=F�C8�PΊ���1�\$�o��'W���k)����/�U^%Y���ڐ�&A��Rn��z�I�R�y	zɚ��G��Tܻ�f.Ɯ&gm���9B:Z�\K맸��@l��a:�d/�Vz���-Uo�@��JJ?��2��k=�-�/�\1�Z+�ݣ��(~<�rA��23���.XK�Q�jl�0l��a0����nv�����&T��}�Y��z��+�	��>E� �����E$����_������
O'1vW�]�H���b(��?�@����Jb���U�q����P\��F�FB�𙵘@ Ȟ�~R�h�k0]��2�^��պ�@�PQƊ2d�1z��N?n��+�-<X�'��>I`{R髊~�攗�����Xp\o�{����H ��B�Ւ�8>�4	��܂�UI��={E���p4�]Hy�f�O[l��}�������"?��T&�Ue�$ӑ
x�^66��Han!���f��i����!W����w� }�QP?ٴ����!N9S��B�*�1�#�\%���C���^{�%5����!�����Ð[�o��IpG��K��Fg�x+ؖ�;Z��J��o�����iBz�rО{�Lǋ��2V㉐#�R��ꢎ�	���A���(U1�d����`Ep�uA3^x)���E�H�d�TP���E�����gfQV��8ل���H�n�>P�x0�Y�{��
 bβ޿���˱�Q�b����S��iG�r�G�ff ����Yr�7Q��K]�$HYJ�t�
���MZ������-}�ą��-�܆	�~ ;B��ݠ@��Mn���w��K;�^p4�(_(�07J��C�Qi��j����L�Q^f���镭�
���r��U �8��uv�ݸ�t�!�*�S�o��ݻ?��(bu"�u3����E+0߁���S�ߋ��8���t)�B���5���&�u���)�G,�V����}x!���{8L@t]�Z�fG���B���D��X��� ve�Pp�:���$Y�-�?΀��c���&���5�c��(�qr��o�uF����GX��R��
��aM*�VIe�hr쬋S'��2�:A� ��Q�RAm,������XB�n� jA�+�K��egy�؄��hA���4�S�$G�3)Ae��3�#P����r?o���qs?��Y(9eAA�.Ĵ�𨃦��f_P"mOM�[[�V�#���3e*e�'�Z��X��.\\��hhm�ϊ���5=Wj�K�j�J�N�4�9�q�˖N������85� �qU�D'8�ʯRN����P�BJ�Fsl��d���m��E����up���*��zfw'����̪����!���Lu�J�6'��v]=L���в5���7��,P�HQ5J�����{]��-癄�Yʾ�MI-��'�9���U.D��j�M<0���8�պ�fy�\x�����ނ{���2��gi�
A͝��xM蔶������D7�6���g���('-��4>2�ioP�r�x�g%�z�b��!-���N��Gr���
���UM�0Ҽ>�6���#09gOY�������L�:j"�M�O>Z%��p f�971�ӌ�y�A"^#(C���)\85fL�Q�S�kX}��f��]�1,�A>'�0���ZL�8dp��B+6�_OcE��v*\ؑ�b2jqv��{�	=���m~^���VZ��u�= ������)��Ju��OC�����Þ�f�TYQ�iOϿ�tD�H��~22`�Ӎ[��.N2~��>2&ǛS?yH���<8�ӻ����X*�6��xU��!��ODЍB�i���B�{G%�>���"���e��q�*]C�jÝ�J����{�F� ��;RMW�DQU�|S&��K��1��O����u�Τ pl��e��!l(�9Mb`sQk��ً@���&�
�����g�|$�{�����UZ�O����u�t;lz�s��(�O�f�	�5 ܗpi�2N����B�|+䪚�w�������e��(����6��;aZ��G�s��l(
Iv��/�(����&�+	iD|�rj�8&_U��_L��໴c΅�:/��;o��sw>&�n����C�`I���-t:^�K�DZ@ZP\�sl�J&&��	a
���ϙ*��`y�T��i���{Z
qcK����f$N�	���W㩢�]gyV�)(���u��7xQ��i��h������e��̺�3�;�%ҥ���Ǝ�-��V\U&�)�����f��L}n-j�����z��j�Ī��B�7:r�ɜr�8�5��3���?�ک����wj �.{��o�_~�_Tb3ǦPA�Y.�Er�cÃ������Wk�P�, �f�=APG��a�]�����J�E�S�b9sq���r�aY���y�\O�*K#:.�'(���^�W�#����q_��z�
��hˤs��s�U5,R`��+���+qH�V����:VMD�H�*~,B�� Ff�C�4S~��f�|=Ga;V��5�ؑ\̃��2l����AP�>�ѓf����� �h�7 ��J8A-�a*&���d_�ѹ�[Μӳ���U��t|v<2��Z�}����\��D*�ˌ{��ϐ��;`h��s�t9Y��Ϧ�Z��<��Bϳn5L-�*ѫ- \w�:q��Qh���O��Qrҧ��E��#bKތ%��ôޜ� 9GU*Skl�\ŋ0i���T���NR�_e���O�"�g{t�w*ͳ�:�����V>�K��9@\�ޯSx��� b�����;[����.�N��V?jK��b[�5Ou�TrPN@�z�@�7�^�����S���
!xO��E�틻��B�}��_���&�Jߞ���ݳ~��
~�b��nr�z�*�������S	oF�ǐ�#�-,�	�r��@��W�J�8}nrA�>�S��;"$3=G��ɉbG���1��P���c����4�OH�����L�d�~X�Z��|Ҭ�I��\��BpH���'�T��:y�P�@��33��������Մ;Ɨ�:��4GL6�V��F'�,Zס��? 215�vZL�<3����+�� aÂ"�Bs�{&�)���)��e�e��.��ߺ�{��E�E ��V���oA@��ΖE8�`���Jf�p؟h�Y������l ���=���������s�a>B^�:՞|�~�K����A=/H����ry��/ ���$�2j���t�\,AjF�����b=,i|Gꍋ��7�&&��T��!�����@K��a���ő��9.�VX��.��h�/C n������I���iY�\D���Q�Y��M��+��B���,��jT�`џ�����@��@jl0c׷�P�@�V)�.P�`cu��z^d'q
L�R\���Z�,�AJ���6�\��Q_@�m�K��W٥R	��h��:���1%�*��}kӡ���ƞ龎ÐK�J�$�}}��S��uE�e#��4�&���"8|Y�Fw1cr|��rU��nهeP����>��8ݭӼ"�5�E�4G��îo��"Gb=qB���(�P����TYgL-���.t�03�=��r�+�qhHY�
�K�@.�ƩQ���)��(5���8�|,���K��n���d:+�#�(�g?Q��m�͝�y/ԡOg'��h�����3�5�w���|�J���Q2u{E���[�޸D��y�u��Y����HGdN$�f k��
_GY������&_ I�0��T��z���Z�j0N�Q�[���}1���Z�!T?cU��s¡_s��t"+��U.hzJ��=��ЕU��/���妈]/>=��hH�NJ?�wQ��gϝ(8�Fv�?��k�M�`�W�>�EZJ�51*��p�
i�|�z��3ݪH���v{���$�㍩O�J-{�Q����\�l��7�K�k�[�I| `4��B��u�S�K�]6��!��O���&.��\����;NW�+�0~���n:J?J��1B���wE� �(��]������J��޳�Ȫ�?Fi�����v4���� o!N��2���%��j�[�ت	�N.] �z��X��K�V�%�ެc7x�7�K_���{�Ze0�k�p�׀ah��Ry)��Q����$�
�8�ўK�A|���@ח(����}�fb��l�z��}�%Sw0zH��G�gV�_��%E�H���s�|(������j��\_��n�4����������q;�O���T�T�5&���Ɨ8�c�v�mP��x~�N�bo����,"�I5I�&�;K��Dl��.1"Y�˫4���	V�K�@�w>C�?��*�X���\�,�]����������r�^�"���F�ֈ����*ye�.Î2=��h�~�ؠ�����E����Is'nDFy�,v��^,��IRԜ�~h�~�ʨ��̈́}ܑ"ao{�uH�����?l[�a�k��VM�x{&y�o�%ߚ���G��R�}���u?�d*�_�ʎ]Y��>m�Dݸv'̬{�n).$�4�$t%��/�F{���zo��$�_�y�^5�؄�lo�''��V,��<I
�h/7H���7��%4�ok�עλa-�J����a�e�":�}Ͽ�#\�!Bж��KW�뙞[2�����OB�F������x�K���S��y1���z�������9�G�L�@g�M���k�m9�§l��y��0�'m�`P�k��8��b[��ހF"UB�i�Ǝ�iG<􄶓QR����\���Pԭ���qI\m��1��g�!��� ��L>,�<����V�2�-���ǰ��,�R7[/�L
��=�+��yK��
�:H��Q!,�-��?�1�taXJ$]�Zo�����%ZF���Z��f�ż�NIm���kש��fk�o"�ez�/��K�/V���ƕ�E'��{h��w�.�����uS�,J�ؐ$�;v_eʟ0�`XX���4T�^aC�H���+�w���Jc�+��GwZ_��^��ε*��u�ljF�gT��t�76i�
c�ɵ$�u����-��v�[��Ţ�Uz�$�
R�|���?��	���ڦ�"�)ĵ�����ǉ�%>}g������ً#dQ�φ���Ϧ��=4p��_8�sΟ�f��ul"3�&���| ��``f�|y����Te���#����e�hō~Ф��>���\�Qng ��e��(O��GW�"ؼ$���LB��*]�5)C}�v�&ۛP�Q�l�F1	K�}?^��g0r� #|���P��2@-�h���s�@(i����Z�U�[���ʗ�QvG�_-�_.�"�茕%����n���ƾ0 �>q�y_�L��6'�eQj�Z������Y�,#ғ�M.�@=���v�O:w)�0@m��"u>aQ�-�<�*��*�;w���e��`��-��`�t��_&v|��/�Wa\-�f����Ӓ%����{��N]#�}`��!�����k��1��+T�Jʫ����w�Z����9X���We�G<�8�wMzI;� �9gn��i,��"Ny4��`H|[2�-,��
J��?��r��~�xc�Q��� B��2����>��/��{vO�Zx��].=�	]��"��''�t��aV��#(|U�m� �&��Mn�����N��w%e�����7���5F�'��UY]O�uheЗr-i�D�k:A'�ƹ������Y�\7B0=��8�>i����W�C�P��x�p�V 8��n��"+a�?Q߈ �FQ��t"#��P6�8o~��:.�C�:k�c��`|_���c�7v�5 )�~ (�VQ���% �����-)b/
Z�"_�>;Jђޣ��\���M4�mq�W�gXn�V՚Y.dw���wq�J�-2�C��2�s\�����ɄG�Kj���� p��km'�a�4\l�иUi"�!����`��b>+`�E��O=�)bJ"7ލ�s��R�R{@�t���$`���,�w�ў	��G��U�(�j���}�����[Ka��V@�6�w�����1FŔ�T'�C$	A}��\�2�\�x/(8Rh{���˳��.����i[î�ɷ��&��$Ƈ_TQP�Li�z��}蛭������E2k���L��6�Immm�0��a�aI��f��I&��Q=g"�M���"����{J�u�4#7LG+	�ȤS��<��}"b��>Cb��u�Z����
�5��K�c���v�b�������EP�d���`4���k�� u�z}d$���a�~3�o�y�i+�}(	�#7B8�7�㽎E�FF)�$u�Rm�gFT��������8�w>(� Zh�ps��z��V��ۡުO�3~m
0[9���6�&	�,c����L�o��>MN��6�Z�t:�oX�r;�BO�QS��zNg�-&M�8�w�����Ա�q�4CZ�������E�ζr�~|/ｋ�@>��@B+����Ea�v(�v-	������	ۄ�37&����CL��:�G* üO*��?:�rA��>{O���x�*��K ��GF����/��p��"��#`,{�������/�7�����[��qP��Եa?Yz����P}L���`Q���&��M(4H�Hh���N����H�G�'�f��X��	���{l@$�R�pa0��Db�{�=�0�s�h��!�f����}��J�4y��.�w��GX�_�C���Ӝ���5̔�-i��iJP@bվp���i�6����mIk�Ŧo}�a����W�a�6
�=�+�����Ak�+�Lz虒��������� Z�s�I��k\'�6�1�*?m�_��Hm�y/Ly��|��~`�����/C婰!f��ռvm	s�����mi�G�K��!��n�_��ԅX;�-��)HH������r�;ϩ��]֊r5�q'!����&>{X�mw��/`q~O���C��7���w��:3}�����~��3����2ٰ"E���mh8q#M4YvJG2��@ӽ{W����Ws�w$��֙�(�$5�m�D�C2�an% �d���ۮFPV5������Q��KY�G�����ǿ2�ih6���	�mg�i>������L�e��R=an���)���dA���Tz)B�#=;����-�� �ifgX&�gȆh��Z��o]������t��).���l���xy?W�����ʈ���/Y�S��)��jOe�F��+�q2���"=)BbJ`&�:��_�#_�����Ѫza3Ue��T�X��9��Kj��j�J��A��8���usX+d�!p�`�ׂ��K��>�g���?���O`=�M���CێO�mL	�m@P[2�.}9	I��d��!����_X�PTd��g�� ���͚�,�gF�}�3�(B�L�,ܾ��(���+�]�)�]�^�JK�Kȇ#��:�N3�%ķɸ��l	W� %�s�l��0�ԩ�<zV�D^�>{��v�󶅅��FO�y����}I��2R⺙C���]����%ڍ��ʪ/���ܓ�ba��V�|��y�8Q]�e�zץq�c��w��'Ƨ�X��!r�b.=2��@B�cߓ��'Ŏ�q��@ىh�Q%e۳zZ}BG�|�K���a��(d��l�9�g�$�
ܭ��}�Ry��8�?��{��7V�����ղ*��Ye�	c�8қO#
��*5 ��Ϝy�Aw��P��5껼�Ȋ��+��Ze6�wb鸌���ϔ>���D�:�� N1i��B�-����-6N�)s�����]r��|S���n�˵�v�q> -h��Wr/d[LPl��xVj�.<ڶa;��{Tè*�+t7p�rp���ݼ$����;wAs�"���b���!�>��8���]��p��y�Փ�$Ɂm�{�!@CB;շ?D�P&�V����0�|9��xFM�Iw֮+�"`Q��"JԳ��-�P)b�D��}�r���"�ߒs�u��/v"	O�G"/੘��ZbԹ=U���\O� �k{0г���ݰ�-,����>�50A��]�;=d�֠i����S�1D�'�}�v�C;=�����6^V�
�2��G\O��e�S:�����_�B^5�Ͱ�@� 98^���� ���o�;덓�Y�9ߪ8&1\��7/r�w?q��D/�𔍺F(倓^�X74�.�mL�����h�)�-�#Ԙ�߫=��=�oU(�����0;�{�U�ؤ�H���[gs>d�{����J�����|r(m��$�9�&H9��H���@3�ڝ�_|�!��;=*���˰vs<�IQ�I��`��7�N;y�_������6�XNh q�*c6��\;D<3k�2�0�$�l�r�U-F���G����&�t4L��k�F)���aZ_/T_��~x�xz������][nǀs�a��O�u�ۉ�2���ZV���ĝ;�O�n��:�Fo.d���ʌh"2���� �#�fƐ>��=�
t̆�JM��>a�I���o�0��A��&I���b?&C�ѳ~A����ky�痃����'�@�� @f�e~�'W�Iث��
bJăz��c���\���aG�Q�^߀���hnY��ď�`�h*�t��c�0tZY
�z���]��ӡ�=F����(&�7��9�ݨx�(zʭ ���ٯ	u��0�0@�䠊Ů�î��NQ_�d�`F߁���C5.�}��MH/�bq���`�Kٷ��k�9�E+�9��mv6ͫxTw�[�y�r���4P�eJX�P�/��W�2�S�;+����	q!BH�_�7�V��qj>��V�ko#�y3��3&Y��*�LveI�À��DF�6'޲�R�e0"Y���|NӍEuaQpWί�T(���U�j];�C�%H��1e��G���R�D����u�;&r6�S`�3��+8:�ϝ41�A;^^ёw��oB*�{��`��G3JRք�n��*BSC�Q��sR�%�2j��Z�eMX���ݜp� �6�$yb��M+�͓�������kͭ)<�`�Uh��<��R��3��$�Ӷ`��a�<<����,K$*�pI
�Y�y=��U��U�wĈ'�#���A.��~�Sے/���6�
j��?7t�Z�N��*��LN��D9����-,��۪��B�A�)�fw�S&����<�sΤ3T��.�rR!�s)�O�u�q��
ޘzdBL[��������%F	Ů�B�w�с��2�����Jp���P͍{
�kU���:g[_����	��\��rܙ�Y'a4ѫ�!���"��@˗���s�|>JȘ�g6?x���!�_�|��u�>
7��y�Mғвd��<=�蟡}�ܫ�@y��A��>s�jTT`�a��lm�RԫӘ�V>L�Ѵ
̃�K���l!Ui�|�#��>9���۲r��}�(�B��"��3�A2�;͘

L��䲂�[��\�������;/*��~h	����A�R4yR�l`f��`�+��J�U�v=���ӥ�+�q�Tꌚ�m�E**yc��n��z]�`;k=��`�mRww :���՘Ư���r5y�0r�Ԍ0�(��)�P*�1�z]���]��N��N�"m5�MWs�/n2�����|z_�Ә�F2��<�z�~|"�oeTX?z����&j	��'�Gj�H�#���Z	3�5���r���}G�"w��L��W=*��7��{�?)L<�qI����UTX�un����h�@dL�_�^�d���5�$i߳�rz=���Z�o�`Q���;���u�=_3@���ǭ��QT/4�+j���_kX�:�F�4���oF���T��MA�/*��׃y�����_:s�H��Çm�)����e�~��o�[x�N���غZ9�D`$H�X#7�D�yu\]5�>)��kuYI���,��Ī#�) ��C��i�l�r�%c�|jճ���1���vN��l�����;飽*YƒNW_���[w"G	�z�xa�cr�`ЉU`oR���Ǟ��\�3���d0$v�{���ΕR����j��҃�Vcp�Ȧn��#t�¶���s3��䓹�=_[�𪊦��yO��z+w^K4�Y���Mm�ql�����.g��%@�q�|$��~��3�:��>�'�`��q�jKQH\����?W���jv�7\��{^[�Uw��ԉ"G@y��!��q�\�aYi(f�fP:�3��l��'X��p��c��ۏ�>�aqۇ��C�7F�4%�����3��yQA�H���	�D箲>�t�vh,\��ALCި��]źu�w��f�}Й��i濮v2�rs�����WKQg7��\���m*Ǩ�z>�U���d���y�z;��!C7��U�v\�Aqm�iE����#��P���c��9k�Y��﫝f�����wNz�.:� �$�;��$�	��T�v�{P��'������{-Ѐͣ�� %j�y��(q�`�&�`�aR]V~I�\l��ʆ��K}3��/��4*TV���ڊ!f�n�~���Ҭ��\�ࠨ�%I!<:�h��{V���v�t�����FW�c��ߏ%ٯ	�tV��uOFe�þ=+��Y��sj�O'��f�����*��t̎�a�� 
���M�ٚ�~!�\��xj@tr@���A��r3��X�S2_�9�ߐ�%Uç�A���7�.��2��4M�N��Sᧉ��73�]Ƒ;1�O��C���g�{�ϩ�K��=J���o����TE{�d�Qv�mN���ٽ�O��SsT���C��&D�� - ��A�D�&�5���k$A�z�p2J��G�~��la�b����Wq|:q7@I7>P�o�b��B��L]����G=/��9�j�9��Y��%m�]^"GM�y��l�3i5�߱��H(�V8�w�^�5��2b)R��]���n:N4�t�-cŵ�����Q�����͑7SX^UJq��h8��A2���)���εc���bk��Q=�l���'<��3�uLRH�#XӰU��� 8�+���N~{�jy{i�kwXp�WF��N�9���緼�N�.3��CA0;�(� ��ѡY4ޅ펚1/i�⟹����JQ������Q�v�t@;����f��k{n��I�L�B�+��yW�o�m������c��?_1�[��N�f�v�`vv��n��G��H�p�}O��Ɉ}���U�:�_[G�nSj�lp��}pS|���{f��ee���� � 59m���.��P$�WY�}�!��_��	>I�A!���Q��¼гl����=	�S�
��7����У�}9.Υ&1��fN��Ok �,�+h_d^��J��;Tr<`Z�H��܆P���"�&������@�ǐ�;P��V4ݶ!����.x����Ls����	��˱~�s�=¯��2ѥ�Ǿ���	��a%�G�)���f���g��Fb�;'DҮ�^�6���sKTN��TO.�%n0 C�m�"N_v�t��,Ia��;�:ץ;]�q�Mgr�_;M[�.��8��ۡ@��u 6�p�5�B�	�H�ru/tRsGx�{Dz�W�P��05���4|��;��k�{��5`� �������)�7TYHtmnL8�q���8�%�N�	%��`"<�� S�D�U�u�~[:��Y�4�����	�|�<IR����H:����� p���d1�~Iߢ��dW$I��UƠ���ۡ�!�֡`��!��+�g��z�Q	�$�hC{~ [��7�j�~�F҇�E��%=���Ķ�Ā&�R��	��`�!;	����s���>�{17�E6���qZV�杚����>N9�udQ���6QJ��KFh�I8b0�����-��j�FDNk�}��7?|�~҄9��2+t�

�[����I�T�RE�'���zmuz����3;)��#��/b�p�mh���/�]�n:�en�>[Bi�O㱘�o0k���&TD��/�Đ�OgPZ������o�4�ņ@H#D��̑èi��^M7SĹ��}!�4���G��5#�i�]�Š;G4��#�!h� �r�)�a1%�0BB�_ե(,�iF�2��p�e�$��`!ͰC;���_�5e*��ܸ��{SK %Ι-��cp�b��Q�u�L��w>���c����Zktw�� /"KV�c"��I��,�U�4���ǟK���y�+�`lA�V��̔j����+�2K0�륗�^���qq4KD�@J�f��˞�F5;�2[������R���8J��v�����n�Wk���Fe
'o!n��K���"a���Kj�x��U��ux;�mK�7�Œ�}x�c,2���?��$�25.U`�R�XqI�d#`�)�wa���H�T0h���y;�o�[	
x5�x�A��hIĖ���Dň�Q���|�'ui}����N2�ԍG��� .������=]�ny����`6�i���x�@������Z{-���׍�[��"�"�N��ËfQ�3E��L�[x�@;��{5�f���~��D��^��zVi��EF8��[f�1���D��ҁ��ڬ�`�Q �!0\`�c�o�D�K��M�k�
��
L��TkBAWM�U��x�E��<.�F��𞿽|�Rj.�G�o_��#�x7:!�&��Б��/�����(�j� C�Aw�#�t!~����_��e#��q��}�9��N�����ۇծ4��d$j�*��X�w�+��zj8�(��������YF���X&}���Z .d��h�
|M�o���(���O�M(�uM�}s����=[0\9UV����SF��p�Р>�٫?��������4$L��*���D[s��܇p��kE�m�:F���?׀ k6�C �6,r�kؾ��?���(Ζ����%��D�x]�JB�:�ߙ�M�K�v8��ƥ��忷u�U�)��ˋ��̙�C��/A�q-JC�_$���QS�/�������ߥC�7ky��V<�|��!�.0]�X�I��I���]єӟu����%�:^6.:�:T���Z�qK�@�nb�?�"\��|28�F��)koE���	�^�s�	�7D\`�.�W��07kW����0��#K=����dʖ&5�c��5D�Y#w@�E$߇�M|�S���9�tO��Ш���M�!��
W�+�%D%�9��z���x�%poק� �{&_�B�W..F�zv:J9�D
�����
���K�"Q�������"���E�U|��k8�����1����W��^_t�{�]�*��L�]_Ħ�4��������1��BF�B���!p�c#*��2{�;�>V���t�:���_�H]+u+���.f8�/�ǟ�&�3P�B~�H�>`,���.��8�6�ݓuOaOv�.�"��r`��^4�!$�nS)]��󇆛n���E�����Z�H$[���׻���d�7vA�ڐ�I���[�c�c`�z$��CW�^Zb�'�_E�Y��%a���+���p�����F��k�j�حl?��eG����ۛO�(H��<����F|`j��@���e u�}l�.�0�A�o���!r�y�}�h���.<G7#��w��z.�������O#̟��F�?��X�AU#���U�$�[6	)z��'� u��^�1x��-h��}yH}`�"W�o�6`�q�iܔ36��7����T����e�!�m���Ťz8���O[H��ʵ|o�&�1��t��/ J#5@l��bk�d����<�n�{����DϾm� Fr�]�8�P�c+"�%,�g�<���̌k�l�@'� S,����t�4��7�`J?bF�N�3�i��_�&�5�ۅ�{m
s0C�M����k{9�^xo �L�X2H>�
NH.�շeAOW��X�x��a��.b��%�	��>̬���ݘ�D����	�@�o�V%��WX���cK~j�(�ǘ�9�>�/�\	M�1�!4�yh����O������\�p���V�	O�u�5�Z�yr�;q?��'��ǁ9
�a�XZ����۟�}����v�7���1 �%��X�P �X�SJ4� 'L�t�ț����`i��q1�1���z�x�=��N�1�R�Qx������P��)
M�i,Ɛ��?�0]����&�U�&���o>s$�66,E�­�1}W��oHD�)��ع�a�e��B��z������1�}�ԝ���mx7��r�2m[�3�V�Nή���N'.ST�;7���8K҇�nD�� ���Sљx9l�Es߯���mW�׊<�h�
�EG�u"d���$9��%�L�9m{�r�6�$�H��W�ЊV���[�\+�p<v�������&�c��
ɞ�4�G����3����%���$)r}�}3�	��ԑ��?�ah;��6����X���^���?@:�U�v��"�5��z�;"���.qܖn���x�#���p��q����M�����?����������bK�L�v�<O�얿������wP��D�ˎ�0��0$������E��U�t0�k�~�l�-ݮ��܂��B��7&��乄�=iY�my��S��]��r|^�����i���)��EW��>mҶ�ſt}�'�>�_Y�;�7ؼЋ�}̓�8�Ít�
�#��s�m��=�p�F����I�y��#��.���WLBz[����	`+���n��h�qE<�B�A0i8B��(�6�0~��Df4A%)�W�-�Z�S��+f�;�T��l��LQ���w捱����������W;j��Ӝ�@�a7j���"F3::9��BFe��(�lDf�']���gl��$ ~4��S����������Pͱ�5!�{>[n�uv�I�S��mz�ogm�����8��&~\�5���X��M���B��2{R� z݇��<���
�FQq*L�^fdWw?��˱Xf=�O
vX��]{�v�>�SLu��&�&���������~ŕ�����T����з��g<UBo�f��D5�[��W���o3E���:�~A֧��;���j �W�Y��MK`��H���T2��[	�<uUU��4um�њ[�w�! ��h�0�	8�UC�Ĝ�NB38�. %���c�N�-c÷�Jh�w~��l�_%Y/^���K�e��I��3�E��}l���y0Ec�������l|@l�q�qP�qݣ�4K.���^�Xv��Wp{��,�S=M�������*V� �/e�2Z�n	(���df�w�"1��KO�g�}�^ͨ�����7���{���J;dt�nѣԋ�g-�%F�
�6R��rX��Fo2%QX�/H�I�2�/�[��v�
�A�zw? Vf��
�v�I���~)W�y'V��:��t���)�K�B��&�\%$\qZ��u��v�	����0��!���67�ۏ9�,�LP/,I�xt�YM.&�!'���`�-B��jy��H��>���m
��;u�	����#]���܏$)�>A��zT������E_b���ۮD6��]��d*����
t�Z�Ի�֒���^ܕ0�vm�fM�Y����ګ�mo�����A�����y�H�cj�0�e�YR����pPo�$"��6�Q��&�x}��J":�������G�;x֫��Y� }�=�DYH�p�ޑc�r���kO�Cp�(���V��I;�M u��x�?� N�/m�1m��f�T�ԲI�Ѓ�#���a�>����r�Q�en�b-d֏n2���R�	��P�k��r����&�Ha�s�6/	��}vj�K�7*֠<���ٝ ���R���ho���X�Xe�����bAQG�1ܝpM6��_;Q�B�Ƭ��%�l2��H�`��Zń\R�/&�C��F��uO9�F��沩M�V��-GG�0���g0��M����	�.�I߷�X���K��ي�gr@���Q��/���K� h�I��8h5�_ʓ5�7Ѕ�`G�͡7� V����Q?���z����Bf׮���i���q1����,=��2�ޫE��օ�/CЌR�����k�a4�� �;lyN��X�rdȬ����Y�r�j n��N(gO�Ӽ!��Pì��Op6+�[��g���~���eU�e$�f �"[-��3v��;�Nb�x�Z$�2n���R�$�2fN��cʖk�zҐ#.��.�Tt��L�4�I�r���o�A'�ˍ�wn� z��ziU���)1��"��4��fܞ����I�3b�j�V��b���6��jS7L���GL��t���P�s�"���=laN7�Z�IF��RT��M=s�M��c��I5aK�'@�W ��#jdi�=O�JS���;�i��,X����,dSp��n��ߴ�z�)��Y��;�48�ɷPI(Ɓ�X1�xAXY�ر&���z�fb��w<`V�J�w���F�YO��ci��rtJx,�^TK5��I@���Yٍ貦�If},���3+�'�m�����)�f���7�\V�ɺ��G�P ��9�L:%}���ȕ�b���>�b��_F3^1(�(	�ܨ[ bua_áv���`�ek܄"	Tny��wiJ��D�z[��n��b���Å�=�`�ӕ�`�[X�Ӆ���� ^�v� z��J+���ЀON�;�?2��RN.-#]$Iy�X6�d���^_v>�G{"Lw�����ݟ{��%�>�C�um*��w5�Z+K5q"����~�7w�.&�c��y�����Y���H8+0v�[nT;S[{�ӊ� SxcB��<���`y<�ĥOٗX��ܢ���ڧ��O.&/��0��@��Gк&FkF򁝡�6�s�BAv:"M�����Ԕ"�����T�/�.$e���=8�i�B�Ħm�r �&�fI�3��ݩ��r�G���﷮�6=��I�B.�U��!�＾۪��\�dZJC{��UI.�P�+�}���^H�2|f$&K�q����}c�Sg&l�F��O������:<�ܩ)@Q^p ����Z�։nW���Sus�S�i�����st����v7U�w߾�&�w����1�Ǯ����JK�<`�s�z�^0�{/�.,�!"�-��K
֋대�^ǯ|:|^]-�IcHI$^X��ۚ/.�[���ڃ��x���ω6���Ǩ$��	U�)����_Rcw�Oٗ� =�T]��Vğ�#���^_�\P8�iB_����o^5֩K��e5D`����]�)����B��Mu�AD�����\W=-��3;���[�'WB.˸�ƴ<�Ps���΢��T����G;2����,�����:E��&*Nt�����}�D#Y�&�(��@'_�[��㢿����%=D��J�h#��@��&!�#���I��V]��O�*�)�������O!Y��yB�����FV��K*�����f���9�ŀ#��+����4��	]��~�E}eQh�ѷL�5�55(�5�-��BY(vʬ����L��?�h�/'|�2N-��H$<������t���zk�=�83F���7�u�c�o�B��oS�C�����U6��� �J��
Z��^��`�d& G)T���э�F�z*Fe��*�✱�/��rO?E�%_�\�K§��5uWԈ����;ЃVm�c-yј�v:�n���,cڨ��&:P�Vr6`��ؘ�G@�w�r�Miv*w�d���d�)(�剹����%�B2dHK�����W�)�lN��]ybIb-��ʕ=��t�LK�n\��ԽdŪ���/g��#������� ��ۇ��p��q��)�9�OS�>n�&�݄ĥʒ/e�B.��dv����vU����o�L��.�*�m-�𾴐g��Uƈ��5fZ�JuI;���T��3u@�l-�Xܪz��/j\������r�s~�(P�>1+/��Y��#?Y�N��dI�
NhULS�
�b���S����)ey���T~��ly��/�]�9�����\���g���Ql)�Y�:��L M��fs�6rs@z�Ym��������B�u]�(#МM}��ap#Q?y4�{���>C�(�X��vkI��V���|�q����䮔LZ��+1TED�K3^<�P����X_��^#���s��c��bK�}�>vHu���j(�=��a���)�7�ũ:t�f���/��[���+������n��x�+�9�y�3 롤UU��cN႘���G��
�笤��!�N2�ά��xԱD�o0�.�֮Bk:>Ь0">�,�/�h���i T�V����j�uy#�\�V�ͣ���ăH|�.�-$e���`� Y%~��}g<5,I~�Q�u�54���7��c)16Jȑ);Ls%���Y�J�:���� ��H-��1��Ur�S��C'0Y�� ������lЩi��q@T�X��z ޿�}��'�Fס�+TJ��&;$�jo��4��~�~;�P'E�zi������"R`�m0RQ��ΐ��Р�;���/X�����L�����T���$#N{#�So�����ߧz���x@EV�S���1$�A��p���x�!&.1�-�IT�q~%�,^=m�t��d�g̦�������h�Sp	�+�0$N����@��&��J�}��Gc���"K�,�q9�:��x�%K�bX$s=!Sxy&֚pȇ2A��^̚��t�4q�Y�
c؎��Q~U���j�������dE	x�����'���DNS���mD���!�−�(!u7�J�0L����W��z��~�V 
&<�"K��:CR�Q�`�@�����̾.�&Z�q_�$�D|<Fp/F<igq`F����bU�Ϗ6_'i9}y`�
����n�/ ���V��5j���H=Ϊ�,���hVw	�uu'�$��:Wz�`��q�Y+�d~���[D���V�RԸ#2���)�J ����Ʊ�Ց�̐�$�� �c�.@��So?�jnQ�Ar顿Q�^��Ŷy���Ge�T�+��aU�M�c���������@��y�S'��4!�,����m��-5�Z�/#���F��S�tT.�x���Q����)�QK�l�;�e�1\�D�!	�`��Df��RyZ�F�@;�����u�3�����"6'hБSF(s=8'��&F|@{E}»frV���[��,� �מ/�frm�aÿ�6���n���M�)=��Omݡ��+���Xflץ}�$�0\`�'�~w�5^[��>	I3���	"�	�,B�8�=0'͐ib���m8���~��A�����c3���ҍx�I�O��љ�J��1b���f�f�����_��d<<���e6��c�E��gF�������T�:M[ɭ�w KQ�>�)ڳ� u
JBQ��۸/����|�[�y):���&m���|;6ǘ����<6z����De��8`C��"_rkB����n�s���G����7�mL�"�>�֬��ֲP	�h��ç:_���K+�{���IH�;hT���ek���+�"�z����5Y8=k��O����B�n����3t��b`����#�
d�;�ˑqN�d���c�.���i��zua�@p��5(�c��oG?������9T����d£P�+��_�0��L������s�[��p���T�Cr�*`d�޹�s�Ć�c%��0����!�5p�˖��Y�*�P��2� ��|���dx���H4,�o�]m�{A(k.)\�D9�ro����Q�����Q����q�}�
o�P�CS�u)��,Ӝ4�$��֧��r���~�'��|�N*����O/^tr+���H��
��`�]���
^n⥞��Y��۝����_vpa��U��6�p��j����k�X���,7T5	�b�i򖴷

��+I�4�򍕕��>�5�K���|˸�ՆnRd�u�������@��X����i<H�c��@��d���[uϤB�nL]��y3d�U�[Q�=�(Z�k�h|�Q�2���褿��V6�hihҀW��}x;}�Kg
��=6�MlK��悤-�	2U���O�����7�[䵱�S�i��)����ʩS��W�1P�L��A=��}y­��(k��GIm�<e[}�ç�J;tR��W:�P-�QE��U�Ve:PG���>��
��OMUy���b��s/	�=���Y�(�ꡣ@A��XNH/��� [d�㒽��8�,*��J���MVm��CS�Aƽj_Q��3�]�_P�6�c��w�3w�f�l�F�ۛ�T"Z_��o\�d�kq?����zY	�~�Ph����>���)�6���!��?��n���H`ʬ�N�H3kw�uҷp�Q�V�7�=��	�f��tLw.� v��C�N��w��� ` E8�nv�8�=zJ�F������B��.aO��ْcoz~z��P�;���.�E[��k�IeY&�����V��7,�g�,6E7 �5�.�T�����6�� /�	�P!8NS�D��¯�k�v��n��5�Ez�ͩY��U&)�}I�e�:�N���>C�(S6��lA��y�e���⳸��)ޡ�D�X#[��'���
���B~�~����̧�������q�q���~�}T�=��:7 ]���Rb�N��/�qZ���t�RN{	���g��ˠ`'ƀ�w�z�R?e��u�^i��1(]�va"'ϡN��2/m_T��0��*[A��@=9��?�4��0i0�fV�0����%=!���6����q�x�x�K���Y1:��c�t�R����A�2�ڞ^��M���{.�5�J�pa�k1jw����ώ��j���$�M�g 5���@�
���6�O���M{<Ĉ�Y�	[E�DILd�p�Mub��
zNdc�x!��B��o�*h| �*&L�*3�]�:y0c�?Gn�r;l$w�ᾖ9�n;��#?�W@K��vo,��=�j���kQ�Ս^�b_�R0��{�-���DU�6�f>�j��qt=���F�9o�����Ĥ2kj�b��JB}��d_���ѣ�|7>�(�G����nv5�ʆď!�;�s�v�������S�d#� �U>0ف�QZe���M�t��MԎ��Z��(�o:U��4�.�~����X�^�q�n,�p��i�l�Fo*�*Ê�r�Ǻ][�Z��Q@tr��D�����g.*�BF�[�G��aO{���&�|t���I�Ǚ���k�t֤�!ʹ	J�Sy����|��u'�_�?�n%_;A4b�J>�OF�qv��ۧWf`x�T|f ���׾~�8�G�vGp�T���$N����PE��(����d���1���[�x}��|�3	�?T����L���P���8��� ʤ�_ut�t��t��A+N5Y�|�:��iT���7K[^�aG���G�����JH���RM}��+�@�x���J��v0�Q:և2��y|0"Qȓd�<����l9���X� V}�|o���$��Fc��!ձV�+8�wxM�kkxޛ��.���ЏH+�m�)�����������_�� �%���9����5JU8��3/��M}���K�y!(��X�B�kZB�t��}7�#���.��IyJOؑ�drp��J�uYD�����[�H���s=r���p�y�UunɁ�LKz�3�ڳ8�hk�������D��ڃ�� M0x\�}bA��C}������GPL(s���&���h���=h���I��ƨ����x0����M����0�����q%(��N�����Q�?9���H���\o)��Y��� ۛDx�Tb2�tY2%�ɜ`(|���V:��Ĭ{钥XE;H(�`:${�_h�(<�Z<@F�ύ��$����h�B����Y���.z{�9X|<gN��YΥRk9YT�fhO'�5��(��=m��t�O65���H`8a�:�*)g������)�e��l�^û�7,Gh��Z����e�4��2l���.��u�#�nR��;ͥ�|k$������΃;B$��`��.�8	n�D��7������&�����C\���s�"�K�����)������P:�)�ƫ�9(�b���.��X�vb�7$'�}�,\ ��qQ�
��>PR%v�a�`�,�4+���ٽ�ej)��5q&#��������M,�i?W�]jQʰ�z/�6�֕`!cֳ�]��V�B����������Z͟������#�z��˗%�b��饆� U=;��7�傳���N�oIF~doK新p���M���U'r��/��]� ���j()��I�qup��^aϠ���������#wNyi�rkq3oN���?���Ҹ{�J�||�%�D[�����W�7-���P�qXq��P�_��]d�P�;�X� �KS�Ej��v���e�2�[����������M)�XE���8	Щ5�}̸�����i��xʋH����T������b|��{�׾x���Qᆗ� ��ѿ�����ڨDe4Z:����Ф��(	�y~h��og�8>&r2� �[F�� ~�q#�����H��s�G����^�3'�xP����X�q���G�z��J�	�͉�O����q�n��բ����$*�E�cN`R�+��p�)X���!؜<?�'ZB��\cZ��j(f )��]���(���鿧<1|b�<0�X''�:܆�@:�7*_-4�q:is�$.(�@�������cֆl��!�0��{�`	��3�ލ@���֖w��t�/��s��v$p	�:Tdzx�t�G6���]�
���F��L��rI�����_�1��=����2��AT��gE<r�nw26�I�k^>�e�T�_��nԌ��i�������&'�59,,(���]	�kX�����&�����=Wn(Ԯ��V2�.�q�@A�˳J�
��{����k�o��\�,���jv�ZE_��q	I	�8Yx7�,����)fV][�k�`�d�-�ފ)�uVY����>9U��aAZD?��nS���#�$NP$8g��[���[�	�Et�z�������ݖ�|���R�}Dal�z�OO[蝆�ܤ�B;�:啔?�bk@�{s���'(�U/�%C��f�N	�����tM���8�77)�EQ�?�<���N�����&he"Y5�-A#�����.�>��m�C�:N�纵���ӏju�!���ت�i�/�tZt�ȉ:/|(=�m}*5Cܾ��>(f��J. o�3��2�W�x���J�8R�������]e5��N��͇k�Z7�BE��B[�)�*��� fT
\'tj`(xׯu�2i$��y���-�S5���?��S�/Z�E�Y�4��CL�j}5.�J���PжV�<]K�������Ȫ�sK���)E0�s��ʲ�������������� <[j�Eq0���#��:u��Xp��+X�Ǆ��
�N3�ثt�~:p!�3"dL��v�ût�T�<���p
#m̀��惐��T�L+`��w�MN��."�����i��F%�1��R�g�w�x�8�
����)Ur|AW�����+z�`89�oszn/���u�M�*���peU�\��Q��^�'7/�����YE��M%e��1bZ����ۂ�
�['��v؝���¼��B<M��0���E+���(_�MTx�٥�5���(���o�4�Ϊ��h9��w��v��	
"�'3��Һ�6���z)nd(��j���OI�����>��?s�Oa��H�]�c�#+o�f�Lۢ����1'�w�����v{W;lao���:q�̋�/u1��ږ���9�`Q��Z�j��K�3 ،���{�iBj�v��1��/1�D��Vpl�ë��
�z��1 ����i�z[����b>-��L9�<��8�P��q����V���}���,�U���+r��9�H���R�sC;��0�|؀�?��Wf�$bвs�6�He��Q�)��� ߌt:}(t]-�/!as�c�$�dY>�e�he6Wׅ�c���GK������k鱴�}�rӬN�8;�wOy1k�5����&$�&0=��Ǡ���6��DLm"<����x+����.��z͎+(�G�Q�l�~4�yq��æ����d@�&|�e~αl|�pJ�r�9T�&L����'�� �#
�H֣F4h�P8��M��А��H���W��.���3�KL1@���AyΙ�6��@kW��w�hbb��so�n�N�W�֎2�p���-�Ck�R�%�i�bX7=�� m0�5����@F��pD#�{���ZA��w�&�UOvљP*��v��Q/&���c���:੤������a��՞�֏x�~b-���O#ĝh�ބgE 
'�F���%g�U���ऩưq쭎��`X?�>�����K<W�z3(��v_zr���l^ŏ����B,���Ð��-�B��#	-�h��R�˥h}s�>+@J&��"�D��x���lN��/��ׯKW��2�n����~�1*���L P��6�r܅J%k_ctȧ"´8�#yX]P�.��������9A�-m��)��Y�/�?�p!>����l�$�>��xM�BHWm{�2%��
F�*Ō��&sOץBv�K��κV4f,���'�Ѝ���@������:ڵ�n.͂�n�Yu��po[��/��cu��u��E	�ٹ���������^]h�`��]�z�ȵ���4{棽^{�#Z@:�hk
���ޱT��kD�}1��]�%
�;?�.޷�/�Q�
I�;�WZ��G0�G��-��iST_��OF�^hݺ����h�h���A�YFU��B��`ܽ�1�?�W��g�c�P����=Nz�7α��'�I�C�n�D�p_K�H �����K-t_\�j��������6 �Z8|s��{�2,s͘$x�ِ�x��=�ŭ�"��jƤ����PG~�p�v�l�5�*�f��񨉥�m�`��y�oNŽ5��e�3�����>�ǥ*�b��	����{�R��m�-�3U7q{?ҿ+�m.`��!��?v��@([`�<��Q���4]W׈ƚ���$I^�y����4Q���i�ю�4���1�v���(]?Ұg�&SN�};�10���%n��z*h�e	T�9����ΐ�c�Pم�,;��g���:<�K�S/
��`�hg�8�g" S��̘��a�ݬ�)��Ƈ��+N����m�.��aZ��I@�d�+zW
,��J�]�6����� �l�i휆���̮�y�Ђ�u�i����Sk 0����w��%�;Q�jP��k��V�U���� gs8&5��#`��xY�44��pʳ�lNŊ�i(�<�Kl�x��)	⊗�Z��aw{m�mkT�ߠ�}��-mn�UW�dG�'���Tv0UK���������}��	�>�l4��H,��/,0�_����k�{�kfL8���$����Ú>�q�}D�$@tX>�chv�+Nߋ�$��%4��H���n��Z�_�k;���
w�$�l���k��+�L��g`hQ��؃�ֲ$����.Z��P����a~Y���c˾=�	�+�t8"w�N�P�����P������C�̡�eS����>Uh܊�~]vW�%a?[-a�|G/�Tp�7=���:����āN3`�g���i7H�:��j�N�9j:HEgW��,��n���*ЊuLk#��1E���I�����6�w�g�� �9V�!�k�dq������`R@#���(�ak�/k�D�]
D��ϝ�����b�st�O���8I����@u�b��l�O��#��1/���oq׮�Z�}�9�[_]�EqG���EK����4�3������S���A��� ;����vcW���_�/; ����@��w5�M
㛽B!s7e��.��?'r�+5���r�/zΘ�9��d��7	j��	��2�� �����ũ��>m�	!0*H�.�w�.	�:�$TW߾ �)�b/������s�b��eO�B ��$ �t�M�y#j��\�*ex]-��4��"�����{t~��p���ۣ�I�	Na(��*ᤸ@��@MQ����� �lk��h����	¸��v<?����i�-��i�IH���N�R�����b���A�'H���U]�pA<ף�b ��e
]m����>���6��5�	�y^/+}r�|��y�{��'�~w�%<�Lޫ��;��f(��k�-f0 �O��O��R7�KK����B�����<�k�`az�#;VЭ�O�v�e�� ë�n �������J
�"�9�6?����qojSm%��/�Kj����PL��z�{�A��=Յ�+<�1�;<Q(~-1;�P�J�|F(�{��RG-ur�8��We�����5���Dq`�{\���0`Cs����%	s%���yj>;�,�iNs0iO������N)�S�p4�;�W�&n�^���'yE$��P���LG׋Rs@R	o�)6��ޑ8��aNgU��\�9���LW+H�a�_;f�6˨��0�yDd��?x!?�3Vhf�	��2^{��CtJگ-U�8?�G��=�b������g��ٰ�a��s�	/�N�d��|�Ӛcs�P9K�G��;x\fYØ�A�o��Y?r����X�<7"4�f�����թ��Ȣzr��yƱ��V��Fk_ݦ�E=:�>�������[|���5��q�SQ%E	���>��G�A"����x������ �ۡ�fIe�8�.����vڢ�� ���X�;T�|:�j$(��ޓ��������5��2D����=���<<���M�sͪJ�`�[�H�+���\���!i���Q/���y�M[R�clL�8f��A����bYb �^���'E�E3�Y�8�#�(��?���?z� mwUkaOU	5�ԝ7�6W�,��u��^9���'���xV��8>'[�7�� ���M���/��Ircck�
��	8bV'T�aQ�g�~Jq��f�_��
5�gJ�ʁH
������T��, x_G߄U&g���#	��}�"/�޵e!B��l�h�b+4��p�5��
G@���z�Kkx�>|����K�ݧ2P�q��q��Il�����%vY��K�D_an�\�3���2�I�h���ς���Axn��i�u=rg�(2O!ZI�#X7�1�nÑz+Lhl렰�K@~�cR���R�p�'���5<`�a�~�1���B����(��xR��:���L�^�Y�d8jL#��J���f�Ұ�I�KFBv+jjhH�7l��[9\���n��5`����2�+���(���?��ê�P��o�ܞEs	�Q|m�WK�奵�Ŵ@��~�7��uI[�L+Œ������(&��ݍ�O��͝����3F�o
��($x����Y�>���Q~�,Ϳ�@��Kr����W<�g;�T�y��Hd��:E"�.�TU�q-*��?�+�
��s�_�@$� e�C�8*�vܭ-��G�}J�/g��`e���t�"{L��;=�I��:P��{��>���M�og���r�s;�+�\�cW��gF>{�,`���8f�}|xk#2�y��!肥���Wƙ���)Rx
���̻�n�b��S�D�m{M����F���E��/���ɒ� @�d}���%��)_jMLE�m3 �����K]+9$}�����kﵣq�y� �N�K8��Q2��h�桒��Ӧ�Nwa�}vV�Z�?��yXӉ�=t9E�B派�z�`c�Ef�1��2@RҼ[t����:��m^}���6����O3��\gݱ:{���ٚ�7�cQ�!���͂�P����H`�R~�rȉ��mO�הO�}z����-�ָR�0rb��A-���+S�(�#�;>�*���n]�ʓ(´}U�����2���v%��F��m=��Ls�vz]J���dl	���l꜏�ĺ�,����y��5�#�#/ԉü$��!�Í5���T%��K.��s�R�-׼�1��NF8��+�659�~���~D��6~�Y��D',��u��nJ�<���(_�+^eT���?{�Fns������B�8��vcŚ&f��c�=j�\N[�w �v�a)�"⼦�ȷZN4o��B����UUM �)��}c�s$d`�&׺�m%��j�������#(#�"
�3X���x����:�$�}��|��_@� ��n#9�I((q���MC�����yKYbEY�ݰ}X*��D/W0�FF"�e��`a��<�XX������5�o���>��lɍ\�ʤ�4�	����Q���|*7`�Ve4nc�Ҁ�b\���"S!��|7�~�CB��ipLzó� ����L63��q��wP��O)�Gy�D�$8�X޿�(GP��D�Nl�w�6�_{D�Q�I^>7��݀
��X�F�W|��/S�3��6f)m�s�a�h3���U�K%��'gA�_i6\���J'7ό�����'�Uf7���#��$M�5G嗐5����:������'����q�Cw͸'�	"'�5Ҳ��U᳆�HL�Yo�Q�(�9��~�pl�=HZ�/���w��E[��m,.L[7A���0P+9���>�m�>d�9�)9�hbZ�a�.?���*5�{.4|�"h��O���!�Q�C�v<=soW)S��H������
#ю�;-{�U�@j~[58�)jh.���r���۞�d/[�obd�jE�p+�������1�/�U��T�x�u�����l�	�!�[�<�����о��%`cdRl;�p���g(@
�OTds�ۑ6��ʎ�u+����"q��4�Dz[��2?}�uL���t�k]N�p��bR�ɒa1R�x2)g�����PY�f�g�ɷbٲDWHb�A=��U��:>�otjb��؃$'26�p7}q�*�����@��X5�j����嫈��x�X^,��A���sO6�̀�ȍV�>�s����jTZ���ZF400z3�q�6��:��%�}9�
t�&��Y+��kö��R���)�,�ìQw=���Q������>��,��-�$Z�3l=�SuGW�&�����#�&%=�,�ei�<������!���y!��s�7�䬡wt�����SLY�ޜ���VQ7zđ�P�J
7|:�'��PD�D��~�B�����92	��aɤ |_�o�a��b��T�U����bRI*�RhuI���{�wV�yl�6ܴ�;t2h���l��R)��D-M+h�N����Yoc����r8�]�u)"�� �ݑ��d�2Tݻ5��[��]��۪�|�M��@@iT�:�hSp	ۍ� ����&�1�y�Z���4*Z�ƕ2e���2z!T�UR����]PY�BH�l0u�h�&�&�3�y��t9���-R�!�V�t+>S.tk�q�xWRp�/sR�E�9�w\��#�Y��]��Դ~�>�	����"Vɾ�<}n]ȹmA��oJ7׏�J�������Q�j]$��Ο)�1�p�~�V}�'�޸G���`@����d}O/W��&��u��|��bz���^��b��%T�Zmj���`�N�^�p�l��"Y��А2֨�9ZH`�Fl׺�?MED,GgO{�&1U�f��� ���x7�ڈ���D�r���d
ZPi`cA9�u�S�ޅ�G���↺F���t�d��xە�:V������!M�Y���E��?�ǴD��w��T'R�	I�ɸX]se\S�wf^�M�#�����Xh�\�V+tQ��i6�/=W'�!�@C>h:��o�J!�<�-ڕ��GwS�cD@�1����@szuݔ��.@
d��s�O
58'~X�~s0�,�ʡV=��r�.��?K�tv%�QA��Hs�Yt�H.���{��u2�M����H�n^_�X�I�&�ˬF9x]%��}R�jX͜�~�Zz��u��nД����ģ��fzQ3h�__�'�-�C�s�&��u|��k���o�A�xA}rW){�F��/��x��u���=G���PϨ�� Ox�XuQ3'r,	�w��qrd�#T�7�(��սT8��z�� �JP���b��㟅�;���U`p��^r����Ӡ��V��}�E��=�bfG�Y�N���r�	E%F��s���Neu�7	�Z¬\�;4�Y���bdJ �|�l�I��AuN6;-��ƶ �����,P��}��c��G>�I�6=R��1\�B{oeU�I�#|<� fVH�ub鮓~sx��纡u�"I����tO��ݷ	��k=#��M��6īT�P帎ߧ�khߎ�*�-8:݋S�E��W8Ӌi�"Km�����p���������L��RU�x��*q-J���. ��ƝDg��6�*/�b�R��Q�WJ��C#��]<����:�h�L�G"��f���k d���yR�<�{�ijl�B�y/��ѭ�~Kq{�Saa�y���΅���Qi�9������*?��]����muӱ�"����g�(�>�r骅N���\�z��&O��_ ��dqM%���2��W&%�ۙ�Y1� C�0I��s���� [B�d���<��>Q�/S��L|9�vs,�K�u��Y2�>}�gNC�Cq�|���;%�Yu�OOE�z��&Í�D6�9?��5z�^�|��!�qb`c,\�����9��XD���i��� =@Z_���"���<g���3���Z%�:�U��R"^��p�VX�%E�`�h����8;1s��DnOhm��Z9x��� lݗ|��1�ύ�J��7"��Jv� ��p���8�%�Í3[/�2}#��(�Pș��;�5C!](�
i��,D�W��R>0x��0D���p��/VuO-5�g-u�p! �BG�pW�|���p6��������F��st�����R+?��!�y���)d=�Omߓ��,:�E���2$���al��"��O0�Hǔqu3���{���d�F���[|F�5Fy���M�v
�`��"���sc��Ib������)�˥0�b�f?�sP4��KH&
3m�E�LI��P@�w�w&��p/q�qL�Ŗ �M*��Q��fi:>��Q����Y	�z�Q&�Î�'p��)�\&���
^&+q����q���aba~D �@)3!g��@���@}��%�lâ�ՅJ3p��?Tzm���m
r�� E�=���jш���dwl�[�M�HK������)��PӔֽ��Yw�;�dݐ��k��0¢�^�4�g�p�Y�xXͥ݊j���3usS���O9r@���Eoݳf�W���1D������L�v�R��Zjo�ĥ؇<�������{���w�bT<�%W��5�q=q��/y����Ďs���f2q7�)ɶ�[j*{� �z�,S4���2N1�")�$X�.R���31X��1�F�s�­�;�(p�dWf�5w(����+?��z�ƌ�XZ�s8G�뤄5�h��֗��
��eqPs�%�\$���%�ZD��eo`��SN=8����V]�H�K�B��94��T�p5�L��������T��Y�o�wz����bcD�.O�����A��>������D��.{Fċo��;H>�k1Ry�%>�a滬V�֎�Jp�0��5�Fv��O�D��Kk�f팈/�	i���x�+�R�����	EA".2g���_TU�/���T������j�����,����0�'f�����r��� 뤧�d�m�w�V8fp�����c6��B�{�A�V��Wƾ,���D&�,Aw;y��������~e�T��s�Xf��C���2����J�yc3�x� T���s�ii��7-��Z�6����]h�Z��_�>��&Eha����E�κ��b�
�̏�H�+��8�ߠnRD�Z-k0�"iۮ�껒+�"��b�v�0?@����b�����ϫ(FS���Q���d�)�/� ���t	�l�r��]Z(n5��7[-c�0�G;f��hʁ�����^�zbEM�<�v���\ ��tK8�#����%�&�2^��T�^g?lV@e�6�$#�����'P?)m!���+�&� Q{=A�˧>O�x�>�h1�s8�rg�aK�#�p��$]Ʉ�Oj��R�����z�����i�Y*S+�Tk�f28�m_{�M/�K8�bX2�����o;~OՇ�H��f�b���J��H�\G�7�S�����T.62��\�z�0�Uʹ��J;Dwu5�*¯�a��C�ZV���qfF�)�4uW൜���d��B~�����0Y��:_�n'�|�x���@(
Ç�>�H����,><��3�gh��+�g�oܑ�B��X{.�c/S 8<z6�d��|,���e���K��w�ԟ���G������{��5�knm��B��땹�T�"v_R�� MY�l�t0B��$;Z���Ʊ�m��hS#5t� ��1��"2��O�	q���N�E�.��fd���x���aFl�u\�E#��8�>�Xl���B��,W�@��rZ�:���߃�Z؆�t�m�|MV�B�U�x�B2�P
�_c���D�RŭJ�_��V$�ZJ+�{i�+���/ￛ�������k�p������s���H�Z/a�I�-����+�Cg�����սػ�Xl��El�A����]�W^��98M1�!
����+)���zX;�����#Qqe��B-��V���͆_&�b���������w$�M�����.W�iC�o�\IԈ��\S�s,(G�e.�����(Ή��`�Kp+�=���ɉ�� źh�obVqp�د�1��{ v�u��&��]G����~���k�Ɛ/�B`���h�a0V��E`�F.qt�pIA��)�0�r��벊�g���涐�ɭ��W�+ � 8RplA�. l�U�o�)^J��	г�����?�F��ک0���T}iAmb4gX�
�����H�O��K3���^�J�m[��Ķ�+��Ԗ=ы;�-�W����,mܥ��9�Qu0�w	g55b�lk����T�;{�xOJ^���P� �֡�rì��%���c?�f$o��,�M�;7�0B������A�!6��
ڒ1�}C��"~o�˺�I��V�C�=��D����{���*��ʦA���{�J6����G*F:E�&`i� ��͔>�F�q��Q`%�ul|k�o!��ʃ�<XـY?���nC]��$�+���K=IawM7v$ļu��0�"�8`�Z�qkA�S���ou����]����Ye��������7Wpo��Jh�>��4�^���mE<O�Fi�Ž a����=��M��wA��7���%�{�E�iw1�c����ʌy�F��>J�w�3�!/Ւ�}�������Q�Y_0�"J��Iver���k���y2��(0�)�}<���'_.g?rWX|ŗ�=7�~0� F�Q�ϊ�^� ��
�j˥��u;�Y�t�8+z�C���SK%Rl3�����mJR�YL�%��+�v�e�uN�im��zIݓ�+� ��W)���)�7ؙ�D؞GY
W*ߩcM�m�걅Iܶ�K���)u�i�:a��sv�笹4�啌اW#ު�&K��[ �fX�C���7~�����ޥ�5������4v�->B(����M�)7�������R�Ѓ0�2���-�&��=��4�}Lx?I�Г��L~l�-�|u���"��}����]�˩���Q�]@!r�������*}��)_3�2�0���7=r�6��t�%;Uaf�&�+VǜO��T���Н�Y��,����c�%
�/M"Z�a�*�m1�e^�:+�)�����M��>}�U�����ǝ8�8��= ;��'�b.�3R�h �{�
�]X�����`�����7�M����gD���Bq�5����es#��k���
�,^¿����v<-�?a����Z̼��hNϺ�#$�Y�&�b�$�̾�F����UI����M�(HYF��Zؖ�/u��F�*'hNy�&C�����%�1�T�cn�3m<�1}����x��f}W;��T��J��b�u�'��� ��~1�lϯ�Ӌd)���@�@?��MI�gϝ�Y�߉�D��,Y�a��C�21H�~@���~Ԇ89����0���/0w�vd�dL��F���G$6���yڤ���+����z5��#���E�#�C/�c�fI��^6�����
��yf�]A�BfWf�7�D��(�]�Զ	<||,$��`���>���0�%x���Tw�Ez��>C:�e0����J�)\�]��Vxm�ʂ��֖|҈��	�����;M?i�\q��A�a	5
%E�V�,�r�|�E#Q�ޭr��� ��n�C}rj�B�w|�7�.�c#4mrrQ����G�?G�2�K�����~$��[L�J�HDZ���bE���5\p�͂�wy�ڰ��ڽ[���Faۂ�l�@BA�bp�L�--��+X��[��/�.RVdj��̛�7��[_
���ؠ��*��5lnnċ�1�s��?2:�^��I w�%b���qF4tҎ�iB����%o�����(��(Z�t1��C�^�q!�)iQ����2|�,��Z�`�љ�uxu�u�q���'�9$�}r��pv;(�H�dPh{�oϘ7l�-�� ���M6��ü��y�p�0��ypS��h0�r�F�*V:�ԐRM<x1�4-��D��́,D�{*�e;���r�;�����v�Th�����2�=�l�La� �kM�#�d���Y"����+K���>��h�+��y���9���a0ES�'�W|D=O��T��[G�!!8���$a�\��͟�г����⋕D�X��R�4��k���=A{=ο�4�ސ}a��&��s���iN�z�k�����">�u��d�Pjkqe�u)?q�?L�)a�๓�Uj%Ŭ�8���ʹ�1!���	I+��d�(�=���ʢ$Ml.Ā�W���Ш��g�Y�l&�PcrA��A���B��@���D͋�AP����F�4Aɧ	(^_f��'j��`��!��2����+:p��mH�%��#�,@��D�K��&�m!r�fc�4�Y�x��I�2�����v�N��l�f#� ��g�Mi���v�}�f%��P<�Nw�Nd�I��z}��f�]9
,���\��p&jq[L�=�"bUFht>_�M���A�.{Y�r�	�M����Z�e����~�������-�b���6��. �PR�� �ŷ�;טSb0l��9z{�	T�4#04)_�ݨ�iML8?uz'S�]F�tJD�x4�
V�7٬'�1���s܆l���~|��jm�a�z���K��b���1��3�<�5� �[�*��iY�%�;�����׶�0aN�N���<�pĪ*�j���"����d:�F����0&:[%`k�g���~V��uI�F��*8�y���ݷ�k[�d�y>��!�l���� B�=ug;�G-%z�F3|�d���7��ҧln~d%�Q�p6D:|c�~�J��Σ���� �l`%o��|`gb�3�̫����s��AZ�V,1��p��������9��`��{����s��y�Š��?�j2B�]ޯ^�hkHv4/*���+��L�2�Z0D�[M e��͊��߄`b�'�W���$�\p�����듖i��[�Ugi <�Ʈ`C+T7̣)1�Z����߁4�&�#�M�?��{�"AgL�D�|�Ҡ$n������Z��kY��6?]u�Ys�=��zh�@Q�7�,�ar�$.��[��T%e�����N��<C��v��i�^u�D4�fv�]�p�Ue1Ϗ��lSsNCS@3+'C��J�䷑�X������j�c�1�t\1�O3	��N�,ʈ�X�k.�%�����,l�u%�ؑ|+_j:��T#m;�=��������و�>��Z	�]42B�k�_�4����C�0���<�������ss<�?@��M�Έ'8�}������砲>-��%�籦ƽ�cf~mQ}n�SٸLbG���r��S�*��'yvR�)�>A�y���;�[x%�U ѱ�eS�"�����c�9�#!�zD�3%�K��Y�
��!Ǉ��î�a�u���,�3?WZ6{]��׹1�����T%8��ۣ\�޵:O�9*��EE�����!u7�)��ӛ)ʹs��Dtm@�1�B�+��'��ŀ�(�*���<�ERף��U0�CCm�Է��:����0����I��>��*c<�_�n�@K�С7lZ�=�`Z��=h�4A�ڞ��eԧ��%OO�q��b�{w�'glp�����&Kl,�Y+N!����ꂝ��k6MJ�ۉS�n�'���?�K2�>c.ԁ��_䒇�Mjί���
��E+��B��N���T��^B_��x}����CȊ�i:�|ǖ����b^D.�_�p���Lg�6�"i[�ޤo	���m�̧�8�p��=Yз��׸^������C��ń>������wO�p`�S�/���*���J�V_2h�U̾���0B����7?��o��v�>JV	ND�3O�f���M"�1-P������+������F�ր']}��Q��]W���Q��U`׶j��7	�
+�!��]"5��]e]���)"� �F����tH�)��e�*�H�
��P���#)�zA��1z��(�n:tRg,{��W��/s���<����k�a���0)X�'J��ǍH��t�>�����{�v9��K1��'!JU��OqfΧ�O`_C!K�/�XM7�3T>kH��QDB#B��L��M�>a��F�dB
�^�# ��+X�=&6w&)kA
�U�[��R ���Kv=}g,�z��#8v�Eخ�B�}D�ɨ�O6����cI�g[�s��k	B�ڈWς�S��L�:�,3Mj�lؐ�0\�������E!�b� ��V��bB��ϪX���<<5\TnJŲ;����X6�m�l�c�55�㹿d�{��BW���TD��� �z
�""�)E�>���BL����6��<!���#����
������(A�� �7#Q�C��7RE:��8\���Mt�qȼ�r�Z���{�5:�*<V�)F6z��$��r���u��+���#ѭ@&Z����� ɭW���ݗ�v�#�_�};{F�f���W֬z�h�[SL3ٷ��?�������,��;EEk�0���怱K��`z����@=0�ͻNm�Hy��]��W�[PL[L�����L@�`@\ �՜L�5��^�O��D��$l�M>�ݺ���#U�rc*�?&�ׂX��1�8�⾹�\:hs�0�K�BJ�`�'{���JJ�����.�N�`��N�c��}�U����Uk�W��יse�^�K�ǹ�n�hy��I%4B��������E���U�?�����A���j����͈$�̷�fB�e�+=U_�;�_�D
����:b�2g|���^�xE�_l��]����`9U��2h5����C�/�HT�)v5(�j�'o��o9c�s���A�?Q@�޴��jM<-����\R��^͈~���W�,}_�%#:)�����>n�R~�r�,p��Ê�mқT�p&��eL�0��u.�K����tf�G�K���6�5o��z�vЈ��4��P�֘S�W$��U���6{]�G���Q܊�P��&,����K�����"������o	���dV���O����E�{;"=��|�(sh��f�F�wZ��|�ް�ZJo\n���mu�*[f�Uu�Â�[۞�	�f�Ag�TW�M'�[͈+�4m�1f*��˜*�1z�M�$.����[���_���I������pq�A6�f���	��!)}qL>d�B!��3�_dm+}0��)ִ��T����Ǉ��p�����q<0�a4j �+l�`�Vp�2���>T���F��,��e@GxƑ=։h�b&��Z� nr�]r�TH_�4��ǖq�9嬹״Q����,���lU��7�t�b�q��Q$]�dd3�F�wN$)���l,��@D�s�hDdA`��R��.a��l	�t�>5�%C��5���`"B;^��|�s�6y�#��:��;`Ɋ��^ �>1&�"������Ԩ&ն�����,fL{��k�L��I�$������΋��0�K2��-+��Cʝ'�^U�q��
����J0뀤�Y�	���~��Ǟs{�r�#[�8��<�Q_ر��g��>kϻAW��ډd4d_y;��pf-Ƭ��J$�kf�p9�r���,����[���S�o�H�T� �W��ͽ��`,����[�,;�y��2�D~3�ž�ǣ�7�UQ��o��[�����TZ��R�|Q��h��<k�$��+]
"72CX_��/_��^���h�;$�"���t8���0�g�He_��c��*�㴓�ܪ�����}���	�1�%'�m��e��,�����+`�BH����wp�O���t�ѰȍSQ��j�{5�������J�=@��»�A�jiT�T�= ��pK��(��+=&�!���{p�uH����Y�<
����p~�["�e���@�����\�,�Z���5��X�K���c�o+xqp�x�
;?�N6{u4�͐�L[>b1�^� ��Fy�Ptn�#���:��u��o�H׉�C�q�Vz�'y>pd���:"\8vl���yE�3���?:�e�:eaY�v�u��{�K[�)4j\Z�T����ˮ�`T�{*�_	w��G|�kމ �M��
�~��{Nd���%1�a��(��ҝ��SA�W�?D� �u���s�F�2sd�X<���7����1�{��Ǡ<p�r����������irA�O�wٽ�j���P�*����\�������mu�P�Z&�gC�i�,�(�j8�aZzc��Ϋ|"�p��Ny$E/��?�M ]�F�R�/�����eqnҖK�s�)y҃6˨���`��`pa��D����1aXN����x���h�:��f��;eI\�E����I�ϩv�u�g�!��{z�C��a��l�mN�¶�%���*���E<oees�y
ӣ���������Ц�4�M�TyŦ]L]n(�ѭW_V�j��vL�ڢ꿍;<�&j�u;L�Z$�X�������/	xErr`��j_��r���f5Y�0 �h�mU�/��V��OJ�w/�>�HB!�|��p���*�!\u�?1���@�Ģ��Mr�M�mϿ� XM��H;���d߶@a�C<�ej��dƥ�L��\���"���iQpD��h�f2f��G�4G��!d�\a�/+[��)4�>���^�Y+JvFψU�a�HDÜ�<9h��@}�X�����B,��JW���^�<��Yq�����*	o�ٿ��<�Z<�_������7hO~�nO?����V
�O\%^x��AI�/~cE�/���on�L�o~q]%}��j��Ru��e)��j7cq�Iemꊊ�2��I{VV?Y����)E��,T�:UvbjE�)[����ӐOb����A���є0d�������|4�Q�"
�\���Z�#��ΝR�^�ڠ��x7+h8�eD��	Br���j�i��V��0si%�3���ز{ЯI�w=����(���hHXr]���H!�b�ެ���Լ�4x�"w�F?]H�Gv�	��Y�y�D�=��8�I���>�K�Iq'{�d\�n
�N��A<��Z-'iQ0J�>C�÷\�B6*m�ڀզ���#���Yק�g���΀��BߕsN?�]ߪO��&��T>�t:��.���	S�W�Y�� ?1�I�yA�gN�����~r�t�M����x_��]���ƧJ���;D��]��o(X�p_ ; |��I�^B���j���K���.��V��@T<'�P=m.]��1ݚx��}��J�d�S*4�^1_-���Y$������t�%`P�I��D�P_Ҝ�R$:M^�I򳵼z	���ŗ+̦]hz���-���%�hJ~r_yZ ��oړ%%TO%�)��z�&'��V��30
����^ⓦ��n�/�d�{5ٳi�6���o�n����$�
��<#k�Hl+����%U�𳽚3g Be~#�]�	��+��s���v����D,[��d3�	�б�^t��0ÆA���8˥���*"
ۯ���`�� I�PЧ��<�E}q���f��Vˤ<tc��,p��ܖYT"U��1J��N�-�B��_Ӛ�>l���+[�T$�ÂlK�cN�
���xd�:����b����|��tY���#lu(�~����+���Y�)�p1���}��R+����:���O����E S���R�$@��X��,V05FEW1�{&���T>>C~�z iͽX�?d�T����(A���t��=]c_�����"	�S�o."z�8�M���k� 	�O���d��0�J] iEG�_�X{�A��S�d��,��6UJx�y�[��P�����u�#�:��:ʬ1�O_�b�?La���e�8��L��hr�a*��щ�Cc��,���M0��,u]GOr��<�a
��r>�J lwZQ�I<��:�q�f�HV���<"���H����qa��ۜ� F��l�?n�Ưb5ƈ�d)6D��;�KRR��G��=�*�0⚴����3���A@����V��!�u=�dY�2���L�vNg.��Ql�'�,R!f ��=�ca�;2��N��g��I�j^:���3hN�2�z�e���*�������{T����J�m@��ӨY&�t�U����,i,G��[K'lM�~n$r�J��U����w|,����2��x����25��y^b����3�|�k��ѹ�V�YI�׍��V(A8W�*h�p�b�&�ٷ2�K�R%GS�͍�Δ���0,8��#%8i4m�=��zxlAܨ��FV�/&���*t�l_f9����< ����<�+jW����oj��e�r�b=��Õ���z�@�Kء�?�|XvM�4���$|a}�I%Y�Y�臞��;�)9�$��ޑ�¦9�,�F�7U8��s�f���gw_�����7�L���źPC!�u��98n��7�VV��<�q���������Zp3���;^9�K'd�Qv���Ka�+�~=o5���b諭����I�������Hb?��P)z��,g���zm��F�ąz��"S^{�`���'��PJ��]�	���7#d�8im��{����a�A�򙱌B�ri~�S�H��pTP��"Mj�os0�Ҧ��7pM��O�c�YS盠2�+ʷ�"!���?�<��utoϝ
�O�$W)WAY�Oy�U��p�i�^�(���P�g�^�l��_L��	������x"p�7���ǻڤ�+�`F���2L͓)+=4i��$��[;wIZ�{fCa�1����h~���Ia�S��������-��N[�ō�R�e�Po��baru"3C,?�
U.����~`���1@T�6?Ø�� ��2�J ��	ff7F����d�N�j7�1p�N�� 44u����W���I�)&GzdZ�J�Z�V�BG�9���qL,����w�1��ڑ �ȶ!���"�H��}��&����y�K��X*f�c;S/� �
dڹ� ��F�gVS�J�i����NZ
1f����	���b��3X0����O�X�R���H�أ��)�M�R�������Y3�3�<<��Y���ڛ��9\O�~�؃|���P#��~y��?&R�:��g������Im�4�>˨J��ͭ���S�k5h��
́��Z��tط��R\��`VΝk�AǴ�0 �-�,t�a���J�֋�В�����B�d�Әh����YD&KR�XsH����[�XE��9:X��8���&�;��X�*O�Z�g�rQ���ʣ�?�aTqK���%'��͢�$��-��YD�'יc�"��ȩV��χZ�]8�#)5M���X���樋8T��0Zq��j�VC��g<}���>�0��Tҙ� n!t�nl�}�nE�ǯ�6_�ܬ�ۋ�����ݱ }*�zi|�X��tnA��Vپ�@����s�PN�d���`|9d��a�9�7���#. �u+ّ
��m1��%�-��r��x�l�C��%���]&1�z��,,�ۿ�{����E����7�P�^4��X�%b��teSt�d�z�=�3(Rz/��r�[��<:�Eg��{�M1Liq.��k@�^t4w'�N�*���N� >7"�����N�_�{�>���.�0�?�o�#�P��Щ�$5���G�R�$�&��b/�� �$������qCb1�B���H�'��e�F�_�������2|�b�-�$Dd�-�ؘ_)�
�1�9��8���t�U���RlP���=yS��`���h�'A��վ��cr�0LpW
�[��^�PD�-������'��Z�~s��D4�U�W�W㭤J<S�S�]��Vc@��I��Տ�g�c��"�R=�x'�`�
QA����� ���In~�9z;���g>ca'x��c��G'�Bֱ�(K�?_M�HP����t4��.v\��
o4�>㫉*��Ѥ��U�c嶢�94�H*čH?��z�����KR ٝ@FM/�g�̕��"�lc���LB�v��u����x��9��s��M��.�-O�=�iw��F�5\ChŦ��]ɟ����'�~�����"ݝoƝ�BP��<��z�P[/�0�������dڭu-G�*.�~�E����@0v�ܵ~#K�;;m=*�c�F��(��9�N�4_*���j�f����������4��*��xr��F�o���%rS���i68��&]�J���-95=jl̡ў]�w�1�0��u��}�}��l���d$CW'#���� �SqOh�E9Yv�=�T��C15(��R�|#��>G��,��
�b}���zb���Q� 6+&�k��T`J]<q���S��+d���òU�Н�o��̼]�K1J�I���â�$�g���8XT[�|2���q��`!&y�/�0��h�0�q��C�xr"�3�ɩ7�]��4�%��f��+>�z
�'nJn�ч� �-o8|V�N2̖���@�0���`�"���K�7?�9 ���e�0� A^� �lR��p��uShbw�Naܰo2�|�	i�̉�͘�j��P���Ĩ�x��-�N�|�־�ym$��>�������H`u�Kc��F���Zg��1��� u.ę0����F�{.�˥�j����} ��{�_���vn%1*m�2�.F^X������o�y/�\v�dc5�t}-H�6���7/�S�����.d��6�a�sSm����q�ܠ�Ѩ'�ʴ�Zs�B����-�RBda�9"�	��4�w��T�g���#B����D��*+��ī�B-�aA�sx��SZSKلI�y��h`л��<M�h��(i[m���͐�R�u�O�iM�k��9򩈙���[\^i��2�+����Z�X�Z.˟��G��XX��Ի��B�p<�s��[�xU��p�x�Ub��%��$�q��;\g�b>�"Cr'n(������jS�����~Rj0$��~㛧J�`�ɔ��$c�ccՐ���pc��	���hF�JJ�����y�R:�L��zv�g�ƨ�l2W���\A����p�ՙ0x����#Gs;�Yʛ2){��ɏK�!���$��_hʾ�XĻ�^�M����5�vC�����̙��3�� /�@W���HB����k#��v�ԏ��������ƤdWI�dL,��#�1��=o-��i�Uua�B~(�4�jlt�K��v�છ��*ɠ��&p�	� ������e@ϑK�Ղ.;/cH��%���Mg΅B$���| �0��$d&�����ٹ�Sx\���"f�vo �M�> �J��x��lyv�=��5�d�Q8�`�G�������i5�+� ���]+�l{q��e71�@�AG���B�cg
,=q��������4�pV�������i"�L֫����`��܏�U������}	���Ҋ5�ҙ}s�ܨ���:,�wbgK��5&c�`�0Ž&����R����HT���1��}���'���oұ�Y�^Z�,7!ս/�9O��Zy��G*1���C��w�3�s�U{��a��9�w�3㚛�<CZ�B��d����w�T�"�+DXGf��? �D\��2F���$��6lⱃ��!�*�P������S����
�\�#wۺ�
ux�qB]�E�S�6c�7��mv�^�4��5+�{�2�]:i͖*�F#�Uu��>��-�$j��)�"���c���vO��ڗ]KAD�
�8�	�Ē�}v���?�Na�Yqd����ݭ�\q�6�s��zTe�|��t��pq��;�&%�|�A�?r�7�lS��܅j��;?�ɗ�`�!N�B��7c��+·�^2)�����"wD8Ǧ�gkbìo�!w�����%���J�e�Z�j�!�{GK�����܅�����dU�k��/�uvκ�Z�iotjx��Z���4l��8���k/b��f�uEImt��f����r���[Zg���v�iG�wO���.4�e:*�k�5_Ъv��;�tNO�Ip-
�G�>���ܴ�Mh�5�Ӿ]6��<���G����3�?#�<���]�Dg���u�A�^�}��DDByrЮ6C�|�A��$L�������BjȪ2���x>��9QKmq���~G$F�L���sz�+�.�QYR/+��m[�E\e	h����5���ٌ^[�����C��G�Rw��Ԡ�<|��M��7�`�=�e�K��N�i~���ݟ����<b6�N �V�X�Dz���^�ă��4�W&�����'$�iroe�s� ���I�l^Z�~���,;�B`�.�D	�l �9�$�&5�0�-�]�'sz��'�]+�B5���R�+^��ߗ�4Q�D�T:I	���}z^v�Y�uHa�)�'ѕA�aV�C�7]�~NQ@�r>y�g�	!#���#W��4W1�[WC4&�\��'��.X3 s�����\q�F:�w��zϒ�\��FS���ح=�ÉL�<x�`r��E]�d�B`�vsU,3ӱ�kx��3�!��{:L�����EEc^{�#��Ԁ��7v%�Ɯx��y��$� ��-o/ț�ɩƿ�T< db
�8��S|���]��}��^=�N�a�F�p�lI_��NG5�/M[�P�4!��'.�`k��e���՝	〱G��ԟ�x�IW�|��l@LHP8?���.5I1d��d�����%4u�HJ��<]جPל�@�: ̦��п<�8��.��֢v���UyP�����.0��G�tk���o��ݲ9�bi��7C���x�����l�ӏ)��k�b�rrXA�4��¸4�\E��J6��䡣*�|MR䦾6Ӫƶ�9Ⰹ�}��碕��@�RP���[U�֬�m��.e��%��e�1��qb�Sw�P��-W�@h���(=g�~ �Zɬ�$�$}?��Na�kK��ʻ��թK\9&h%�/ȟ4 ��u;3"km��`�OT����n\�WuM��	Mh�F.,�PY��m>��P�4��3���9��"��A�!�b��7�8�*���`�T1d�Y���	�
#�'|���M��A0/!�<A���Bfu�i��A`�? �<�'6n_��sg�4���Q)(�������2J8���j�]7�,���Рư���W$����#���Y4��G��h��\S�2�x��K	Q�[�4ֵK\'�^Ǩ�:0	f�3T�X�IX�uǙ���"�1Q��������J�C��\Ɠx�c�� ��׊>�om[�^����Jr�s斺V�3���ԭJ�2H������(��>�m��)AJ�����m5L��̝�٩�h�*_9�0Ä��}��H::<�Vt������y �'�:m���#~NG��F~3��ŗ�6��ݼ�*�9�yH'*4�հ�KuxԻ�f��[.
��GQL�\����BHc���K�J/���Q�v�=2� ����1��I���a��ɆI�LW�t<oN!�� O�'�������O\O]�f��١�ġ�+���].�ji��H�����@���Ճ[t6���e#��v���>�a׺H��ͅ{��b����k��!U��!�ԯv],�\щ����z�f�ֿYb�"e9�W����y���L.<�OZ��fò�����;]Kg1�!Q9����0p�n@+��DR]���{��K��s����*�w��a�Q�E�i �v���<:U��{��em���� 톎i���]�Ra��1�;��*~��75N�_'_8��R�U�ւ��؞��iq�j8�������<�
۠*\��d��#����.�y3H��'��/C���9;���Q�^��;�h;���]%�R��V81�N�xd'�rY�{�+:�%3���7�WT2���'��6��?�R�������]ɋ镢�:��������hپxT����O �c%seoA��:W��u�i�:����T��9<�!��z*F�g����;r�D��.B��;,C7�뺔]�	������-5��sq��Ҍ���E_S���z�n�(�e���f�V�K��SZ�%��4�	۝�-Z~+���Kݞ���p��K��Q]���d�܎�ofI��c�d�黫pU���ץ�Ӭ�ܸqّ�3�D|�Ge7����Hr7��V]��(��������0W��g�00����vj�0}m?>X�5TIQ#��B0�z�<_+��.��Vo�4w�������c
Wd��+<�l*Ʌ�Sy|���A!�F� 'U�ɮ��R֖�4���u�[k�ԕ�æ}����퉁�a��vaۈ=�C��a�%�W j�ѭ78�E����:�\���y�"dL�0p6�H�'�|���hĽ�:������3�펉ZN�֨�W�I��J�����D:!���j����m~�L��c<Gb�ik��@>�8�[�`�6VGc��5�qE���ihZvk(f�$S�k�ǷP��ڽ*BM���!�{�6Q �x����|�v��UwU߿���<0`�7P��ĸ�?�&��f����� �W�a�
H\��S�MCYU8�fC>��'�(���jq<���>�s֯�β�EW���d�����콤;����g���b�ډ�4��M�@��<pT�.����yB2ob~[I�NE���掹~_�ԧc�qDO��>�AD{���<x�Zg�l,3*��m<�x
�R]��|��S�v��oz81�S�I��_�n��d6��e
��Gx)�fń�F��`�ȿY[-5���B,
��0]���a��|�\�
#�p���2�*�^��E���J �Ҕ0���m�61�Ŏ�R ��h׼��q�7�����\�7G@F�Hl��ޤ�J��|��Dą��ń�I��>V��+;��Y�׉�J�G���a&��������PH�%/�INk����"���j�xR5����r6S���(�	�[aѺc���N���חcG��Rq��V���6������ҩ�֫䰁��N
~��eC�2�>G��hM��0�xho�����{9��J���e�|�����]���vN��[�^S�nN�"[JC�OA\;���\4��s l�	4���L�EU���`0: �� >!�ҔF/�����Ed5��ϯ\𾌴�EN���us�PK��elg�3��m4��@�`�^���RznE��Ӑ�1��,��i��g�߯COq5Eʂ~n>\�t�Y�$�>�k"��"�G*ӑ�s�j*��> �Л~r\U4S�(�"�۲���e�:�/B����|b�ADy�S*>�{_�B�FT�0H�� O��w�l��s�����0f>+M���M�%��"v����� ��@�L����#�]�I5p:8���.G:OJk��=��d(��2f�a{��p��X��z���V,p~�P���U\p7�;(��aS��C�ljk.�W&�_��^����k!�e��ɚ��- ����/Ʉ�g�<Kym��oI���lQ�Ɛ�=�#桥X5+���̿�b���kX��P:{4ؓ�t`�����w���-�k���C��ol��^����#��%Ϲ�=����0��^�F^����5���t��o�_����8�V{�;1�N6]u,�{�,�ȯ�t�0��	��"�%2M8IV ��p�u*I1�"}|�AT���0��#&��&|�IB>B�xR�WD���_� -b-,����[�r�\�	�Q�[���!�d��@�0/م8���\}Gh;~��D�6�Z�_�.c�z�q������o�'�Wj�s:�!��9�&v�{���ab�*��k��:a�"��Rw���I��y4���^��l�>���JwCS��+/+�غ#*6��C�32�y�˔*0#���Dj���
��cY�C��V�xhm�L�4�����?�`�P���|d۹�Y"�~�*��d���۠�m�A���������W����K�l��{��[����� ;�����$76��ϪU%v�[d�v;q���������8j��gL,w�^p��p�,�h�R�1)�C-p�
����^:�-�|d�<jn��B�l�`��Y �@���6���lD ����_M���ɋ����n�K�gB�qn��:���aۇ�0�����h`��%��>�1�Ե�|�_˜�dn����21���\g�iibЫ��&�sc�~�~��.Q|�z۷��e��L�Ϸ� ��}�K=p3���!�Rh"ZbIG���'p�߳C+N��6qԪˋG7wX�9��R�~W�|�������U�]U,������Y�p�{sϵr�Ce�<�N��5I?�M�u�^Hʠ�O�5�g�;�7
Ɨ��*���O� J�4(�YEZz<�$�Y�d _�gW����������5S��ٻ�mX�{��Z?�C
��Lb�����sk�޵$o�����-��ו��?s����g�ɗ��}yW�\�3uo��{�f�*�L@�Sڽ��(�-�����mX�TO"(yy��y
�a�3�M�6?D��<k�`�3�o�R��;�@�u
d6�`ߴ�봚yO심'�,T§�+ψ��B������&�$e��Řq��P�a�>�*��@*��eJ������Z�!�߿�_��-H��sBc"���s|(��B�G�Jw��D[p
Y��ȉ�%c)&�/��y"��r�S��K6-�[��X=
{к��Хw���;��C��=���̊�T�|�"3�ED������X�C�����ZyRQ��>��xj�^2���?�\*7@�ℽt��X8���&W�����ꊔ+#NZk<J)c���K<i�I�I��!����L�G]�3o����|`�֡�.'	l��7^����"P��A﷔@TEP����d.,Vz��	�����q���c��j�	��1SP2��+��C��X?�x_��x��ۚ��7��Ƚ�n�@�xq�v^U3A����E��%*�N# 3��	n�&ѝ3T;��j�n�ٺ�S����#����� ��0��Wo����t��g؏9~��<�xQ�,�Y�%m�kj2���34Ñ���D"����zn~�u%�����~�H�#�S�����0�����e#���+�?��i��yU+d���V����!�!G<�� qF�:N/:��B�6�C��Ip��_	m�GD�Hr�
Ѐ�eF�Co����S`�T����ǘ�!��#��Z���E��f�"�r�돕>o�,�,��%�s�V&}����g��K��#��D�k?ŧ�d��ʀ#��*2��fr�ȟ=��t�>�s�U�Y-��Z�ύ&ju�I���-%��r� Cֈ�f�"J� �����zk�)��������@i�=���~B��FM�K�S�^��]�X�D<��rm����C���!�s�0C
��f�jZi����^��!�!����a�?�����$Ri��H��J�t����~��$^�& �҄�-�6 ��3E���q>�� ��U0��
�أI��Z�;WO��No��u)L"��zN'�Ȱ��ˈWˍ�K�{�S�wS����&D��bM��n�_�G�Ȉ�c�;������ݽ�^D�C�n�q����,�u
���˶6�q@j\}���+�H�@I��>�������|�66@nz�m#���DT���6��^��C�n�/��7�����E�AM���<���DwPs�+e�Alp:Q�g�N�!����Ӱ\ǻT���>��M����38=��G�P��P��¾�x���U���A?���� ��T�?W�{-5�GK�Y�hD��w[n�ɝ�E����k��w��+(�����^�:��ZN���
����h$c��]\����l�C�ݝ��is���niv�xBK�8+/�λaD���Dpu��W�!qb!�b�M�cJ�o�y���^[1�k¯E{��wM]A3�x:K�ΒA�"�z��J����N%�N8ƨt�[���UČ��K�i9�]J�;���t����#VMK���ܹ⮡O��
�D(b�~���I[�#��-ɇ������f-Ҥ����(�o�T0����I:��q�㆔�G	�%9P5#���XWZ��Q��qA�iP�=��6�4#SJ�I��c�g�P���"$��Y��&��?�⾓\�~D_��K�F�C��U�Tm�����������O�1��I�TQ�7Zg>��}]��o �)k����I��Q��!z����*�?,�?�h�X��$�y�#� �)�*aѴYrj���1�m���nӽx�?۷��ሩ�	l�E�	p���l@��ůV�h�"�]qM�
�(�>��:���[��J.�i\sPŉF ;�C��O ~�N��5������`wY���X��=$n���ADk��� �!��H�Ix?P�o�Gi���
�̦�h%�t('r]�l2���K4=AkL�$wy�iG�6��bY�����Y~�-9�_X1��
N�A�#!��B|x����{��۹Y��E�
_��`��\�Mݚa5��- �gо-�O�1Lh!�\���\�/2o�G�inin�����%|]��M��,�u��r`മ�6�7�_�G���f&�R]~�J�|�Å|����I��$@P�6�_�7����]*%Dl�L������ �ʏb�:xqzn�n���u���ŦD�gKQ2a
4��=�j����ȍ�},��Nt����s�|Yԟ�M�Yk]���	��� &46>TjJ�@Q�pVBg���e����J�!����3:��SKM�p���t�(B�{���
]
ؕK���%��.�M���CU�g2q�^��n�f��'��������ڨ4�t?[��[���d��hf<�!�\��T�]]����ז� !�!n)�o���םM����; ��H#̄��:^���W����#�Z�ت&/@��?A��MALN=���/A��=I!� �܄u:*��ѐh�sG�A\����[�B\�25�(�q-Z��l�p���c���'��{����#�MK��~�
[�`c��	*i�A�.5��{P�<>��5���6�Rd^�tn��r��>���I�K~̎��h���\$7�dv�6�uc0Dm�!�|�s;դ��;�3�E���ư��o;8JD���	�^�YCJ�<�FfMj�5\ ���]G[Hgҗ����M;[�6���R������&��ExR�+�X��>fTTB���������G�9��j�8s�k��YV��7H��ck3�t�}U��	��RwZ����>�"f
�h�!��/%��KC> ��,Ʋ,xB�Z|K��jCC�D��=�;����+;�W�A��w����]��$EF~Q �s��d: k�ȚE 6j]o�+xv�xjiP\T�+M�.K�ՒN�j�1%�<�+fc0I�W�B6xtP����m��.�zB�|'�4l�Φ��j�˓q�8�?D
��h���T���ӵ�S�}st$�Z����b���� �|J�,=����QG[эf���>�>!����~x(���xm��.�X�� �ʔ�����n�I��و�!T���d�s��;�~*��9B��շ�7u�.�rNs�G����4Fz\u<g��$���J�^Ub�㖴��q`����Ht�S#"7�����~��ɉT5���g��<��p��{����(ф��X9:���n��$` "X2�t$�}w�o��bb&3]�$�k%�K���kV ˻в�4�FF4v�蜰��9�g�kAr���ޖ�-�ډ�*C��^p�Q|�2�1k5��q�`{tF_d�u�x��wde/�?�>d��Q�1mV�O�{�,��=�������nT�h�\-,��G�+ˌ��Z�a�'Ί(�>��p7<�0B0Pj1��h��{�mDp&�!狸ͼ3JS�9��R�/�X������5t�ٶ<&�T(q

Q��7¸���P�.���G�[R_�viyC�|B�}J���4�'=#��k�W��51_!��CcY��ʖ��0a�	�:x�ۍg����#´�lGpXw)}����z���)�I� d(����W��:9G�c��S0m覝�$3��c��&G�B!�ב8�2Z����0�g��K�>�ͩ>�i;z�� ��ۗ��IW!���^�Ȑ�i;�.9���1$p��F�+�:������޼�B�w޲b7y�ڗ-
�C);h�v�(����W^	�|u�?b�p�SL��#]((t�s���ld�v�8)N�#ɖ�}����a�*�P?c���;KdGl��!��2�K�W�7ѿ9肷*w9���2��cy!��mNY��նf<H�� ��Y|t�%w�t��VC��i�s)M�]x\�y��ȋ��mb�0���FY��"^������0w�/�a���mX�m*r��[��[���a�����#������e�	��F�O�h�aR/+3����ނ����� �X0��1�t.�;m����{!n
�����Ѳ͢8�!�p/}�T��
P�(��ޣ��u��!s2�[�(���7_Ҕ6T�Cm����Y�HT���ZD/??fP�>��.��C$ju�pI㦣��9B�Xg�����5 H!q����d7yQ���/��5�J03�Y���W��-�Bt��-[�1�<�=/����LV���9_����;��.�wW7��&�8Ńގ��A��^P������Zk��(��\�Wb��e�G�˂\n0�2���L/�AbM+V��������zܶ�c3{j��v���k`���O�`1h��Q�(`���Ag�_��i�fږL�sv(�`��9��m�{a
��(?��6�Qlhw"1\gΠy�g�d��LX�Q�Ɲ�����ⶔ#�&�R��wt�>���Ze�����Ѯ���O��у����ݼ���S6v��(Y�#��<�Z��M�Gb0� \��+k������X��"1:([ҁ���׋��t �qzՔ��g'��'+���G��&��v>C���x�e5?���µ�.K%>���tI&�=�������e���j�W	�L=��2������A����G����ĥm���n<?�	70 �7�:D粓U$�y��<��<�hO$�~e��z����:��1re������g_���W{TBK�ٗ����s�II�,y6�f�lPRW�ǒ:�����c�RP���t�����D;�����f�.�=�HA�!8,Uw��8�����G1���b�;��9;�3�J�]�rn��lK��d���Kr�gTk�i��D؋��VJ���d��Y��HLU��ݍ��E`Ck��]��cf�+�l�{����k�C��%uB|X�Nl]�WO�J\�,�Q�aE� _U��I� ��gR���՝�it(	5�pLN��L,}�?ɸkgչܡ�:.pf�6c�ӳu�~��]P\�7�8����	�H�H�ZK=�b�͇�m�0Y��|7pD[+Q	ΆQ�֥���5ќc�XU4�1Qa��k��e3�.���l���n6�=���e�$���Qر�B~=��
#�C���~�mU�(X��:��$�z�� �>'1s�zм[���O�wa�l���нC8H*\SH+%}~��ϣ�B���q�2�R�`_�Z-�9׷�)��d'������N�3hab�J?7�k���e�����&4Dۈ���S[�v��h��$y�#�l>#���!A1XQ� I\�kS����NǼ@�R�-���ř�h��&	�,�{'����j(�Ѣ4����&�Z��9Is7�����1�&V�L�x���f�ߏN�8�E��e�:�DpI�*iE�)MC'�8[�`��}�~7�L��_.�#�X1�xB!�-n�R;.W���N&;|5��BB,��}��0�X�F�!C�"O����'W�s&pۮ;� N�e;D��r�(����\�������K�<)l�ЌVA�Л���>-��+H7Cy52�;5�k�wW>�A������GA��ţ�AR��e��9Ot��Q�̐W�s������-W��,� �Ԉ�P%&nĥG�ܨX9b�-���	���P�j��!���Bɀ�L���2�L�<�[L�8[�d!;���s4WD���}L�4lZ�ޗ�>Vm�җ�U��~3Z
|Zq��̾�H��xht�Ps��?��D�p�I[�eacʪI���r���5���r+JE�	8.K>���>@��A�]6=G�<��e̅����������d+m�$�(x�H���Dv��b�<���l��#p$	��9<4+vė��6:�rL�Q@�{Ru�B	�qs$anV�}b7;$�Z��Б�:3t�\?��J�oZZ��z8��5A���IH�(�cؘOmG��Tb�W��g�I�$����O�zW{��Ty(0���=�9:�eAy�I�&�e8���9ɟ4'_�_C}���9`�b(>&��%����Z%�|�x��>��n�6��y�Hd����h�RN�-VЍo�[�6�W�}��uk���&�c������%��=N/'�3����\�������Jm1<]K�L��]�E��3�4��G��OYx��f�6��2y����&����Q\���/�5aI���B�;��(=�ٛ�P����`��	��.�Pb�5�D{PL��,�\Y��l�
2رtO��L*e�#��GV�,Iw@�^i�'e�l�:����^�F�E�cʹ=��%e:�V{�B�foqS"���ɭ�"+�Y��bֶ��b����]N�4S�.�ܽ��B�?ù<�c9�8�H��*Ga��K�� � �Ŵ�o��Z�7��O�nv�SC�S�t0D�F�
�~�z)g\|6��[�C������~.`2.�Zr�Sc̼;���i�@+��̯h�>&f���ܒL?=��_�t�a�ņ/�A� ۊ���GB��A׋��ua���`N��Tf}h����t��֜ r��a�J��>�K����qR���~ܾˉ~dM��ܼ�}^��|�"��:F�aR۱��I��^҃���������ȻKh}�Z}���\dt�R9"en^1��ǂv��	���39�V����=*��h�/�ӓбv����7�.�k��窇ێ����g"���p��2	�+R~��9e%�7t��o`T�?k��-(��MH�݆��7�PWC�����u����z�59��\�^��W5t�.�,� �c��.�j��=hY'ź-k�5�#���8��6H;I�T}J`$�\<���wJV�D!�G�\ڷ�1(���ԍ<��ⰳ��dIL9nH|����6�6��g��?F��I�V�H�n����ܓ�_g �T,�oC�½���p�B�ص!�?I�O�]}���	:�.��16�/P�P�^�Qe�7Q��I����;�[B���\��N��tѪ|X5�;C������ro砑�վ�Sr���[�sr ��1l��4*�߁1�`�nׂ�W�A(n�D�G�Q��0k}l꾐P)^��g��{��3b�]��s/3���dEI�lؓ��^���"|���N���Ik^7]�fߪw1A��	�"2ݗRJ�'Gf,@u�+GX��h���^"i8�F"�AFi�Dp���t�|�E51'MIL��weWR�\�����i�@�0d�5	����)	�5N�"V�DC�5' ����K~K���˦tP��\]�Eݢ��(��	��!���Z�]�twI���}�
t�L��e�v�
-����9���IG�Q8W�.~S���Z��&ϸH�7�������eX�wpj�f����@�<��ð֙��B��ۉ̅K�������#����}�Ç ��[:�/.Q���E3iT��:$�,'�*3��)���)�2J��"�FyG%�ĬAl|�l��6C!��\��ǯD��RǌD���.-}��.y�NN��(#К@�6L_6ʬ���&�aB�M���� ��3'w���#��:t�ʌ�e�l9��>]�Yc������i���?$R�~�m��ց�@���
9�za���~�)�`�E[��ay�'�m?9jS@�ґ�/a�9S9;n�ς�S��|]���.Rd�e��e"4G#�Λ��9�nR��ZS��*K�6�M�ӿ��t��Yt	z5�W���Gf��s�"A"Wҋ%�&�VQ�r��mo��g�+;��Ћ�xD@"*HF���2%Xd�Uh��N�t����+4�E?x ��2�/KD�W.?������e�+idy�;?Ӌ�Е�B����Y������w��$4�O�>�E	�D�ޭC�"J���c�2����a��W�J����7훳���{&b\�ד:K�V+^++�����p�*��S�=������.��BXl�U����qL���ԠF|^\���'9���Tf#{Im�����Ր`���8�ԽF�-��!;6
5�)]����r��8Pw��?��˻��_��~��'L���f�mX��e��T���&�W��7@;���B9���Zld��X ��f������	��&RV��?_	�Z��,p ���Q�DY�$mڮ���{P�x)�Z*��>�ɦ	�r��x��S��Ъ���ԙ_�9hGhdӻ�!����	��sy"͝03�53�ڳn���@w�@7 ��?&q��Mr�*nՒn�SG:r�M����#�)V�AG�v\���� �ԧ�0���i�υ�I�(�5�RU�	�����'��m�uhqNuN�/�gZ�;���W��p��6ȓ��W��#�!Y )	}��8�":�^-�ej�2t�~�,���̘�P���R��HR���
H�?K��d��P�+�N9--^vh,FTD��<�s�g�)˲�4/܁�A�oЉ�	m�Pg]9���B��%7Ό��O��(1��vɜ�ht��Pf��8��Sj�X*<�^\��|]�S��{��q���wQ!���F�;�+�,O��m�x��lk�e�
=�WB�p����b��>#�V]OGHl���'����P�i�)��:�i����_�u�BsK�|�5cH���D���?��#/1�-c򯧏����'
>�����SPNX��((��k�KW-�G��B�����3�:��V:���^&�\�B�X�"d�xw��8��5>�`����˱������֨��j,��lhχ�hz_?Jɨ�{�;���VS9��V�Z�*��x:�x(+�͵^܃�" {On���Xa��m>�˝����͛Yb`Lq#�J��E��a��T&�t�Z�nc��\�i�����fU�r��y䌄,�[����\DiK}Bci���ҷ���o�r1��h��g���;fBH�ڹ���'VA���������g��<���sU���ݗ���1��!�2s�7�즆�|*e�r0�5�8J�K�{&l�s��D� 6f��8x�X#��V��Q���6�̃{�@�-"M`�16��k��(��_!�rL�}Gs�BF��\�V��@jX	�>!ME��o�|s�ʍnL�����X��
?�	��њ���Cy�l&��)�qm+F�g!9��������>��~¾���X7\�Ѝ���\]H��W2�\��D�}�6���>����ُ��jc6�t^ 3p�p�\f���dX���&3���C)�-/��En���41�+�v�.�6Xߥ�Z�/�nE)+��a�՝a[� �~/j3F���nn���+)G�E�C1@���R"��rӑ8��(�Ց�*I���ȟN+	��ٙ
wA;,���B@����)�Y�1Z��:ﴵ�f	�4�BoE���̈��������^'0xn-���M��5���ܟ�+�u�����o���{4���$�{�]���@�mK����O旣YJTO�]�'��0�:'��	�9��t.K���[0jX¢H*R��Qd�S��.u扭`��+hj�M<�UL᎓�֨�EbmٶHq�Nܩ�N�h�(eW��S�Ur�R�����+�M5�Ů�o��� ��鮮x�)ٓ��s�S��������@9J�㴧<�����4\�&�<��k\�!*��DD$��l�4�ʿ'o���
���oO�ٗ�ZQ��.A��K�gӧ_JX,�,��P���phmlv}c��_��5L!֥��7�2�`����:j�W�3dI6ؽ��ߵm�͖:pr�p�+���n��u(R���p����R(��?���sa�}�F��\���N�E����=x1�}ٔ�a���U�t���02bo�;���MW����0�yسI��gxP���B�)-XKy��X��%G�.=�촐t��\��	b�6w�I���i�=��wm��'�����>_ln � 7[/��in~���_)���:��!�ОVT5ݷ�@�������ڰ[�'^��D�k��f����@l�ZI�����є)��q�٤�T	�m����d�k���C��m_J1��-������F�$���2����9��Rc�8����y � R(my��p�j���~Ӱ���@�@�i5��'R�����g�����:��y9\?�~�qKl�[%}�:�gZ:��&��������v��A�fJe'�M�8^�.)�j��n��qc�U�XǼ@��G�3t��]�ġۑ?�;�X��@�qj:A���D�����H��i�5�!�$�>��6-��7%�z~@���^������kef���2B���h�\�4hp��wT%!Ġ���q!ob���07�1p%�r �n�z�n�l�������=6f�\{�##a�Έ{Kx}�X�f�2��k�T��F���`�~r,��$/ڇS*bX�<)6�˂����[���K5-�M�7t���>hg܍<�*@��Z�����r`�ئ�c�H��~^r ̶� 0q��l���'�4���0ѲlYM�p�Q��:�B_Z )W"�S;��a�%����_C>Å�{�L���U�Fih�����
�2�a˄�pF�o>���MR��ע!���8
�ڸ�٨M�H�����5�9k1,h�H{� rMY����b�u$:���1ȍ�24�El�L^+�< 8�#K�S`�%�a@G�XI?@���1����L���6��e`"�"?6�h�U������0��Q�Έ�q����]���;����h`g�mA�� ^6�a�� UR�g3��F���g�$Aê9��dw2�{��� �����w�e!��:i�!H"zm��A������nk��L�o��G7�N�T����)��.�Ā�%̀�h��%�A�p��ݺ&t�<�s"� �����x�x���\ya�p�+Y�2u)`Ϫ�!^=��Q����g��c䇕O�.�Hk�Q�㷆�$����4�y��|�pǙ�i;͉���Hz!�μn�SS��E�k�t7��6��)v�˥�����d��c9�G�K'�m3U)޲�� ��Z�,�s!J�/|K�َ��3-4<m�<��~��/`�MP�y�2 ߌ��f�͂�{�@�(�+kS8�L��[�ū���Ӡ�4�_�o$RD$���x(r/���=��+����*����Ϡm�١��%B��;�����f� w��L��G��v�"&[F���Y�iv���儋ĕǮ�J�n��6�1?Y6���CF
FY��^����"`F�\�{�?To羗ge�|ݱߴO�`�o�H��յ��af{R��p0W���ZER]ua?g!o���/�_@)�4^�y5X��Q&�V�"M�N�o5%=��������'&=�1}����$�a䆓\������9F��6Lf�����X�@H��������Bu6 �A	]ԧX��aa�tM��Nn�4��S�C�����jw������ط�EqA�
�0�_�?�<�Y����oF��b�穎p��O�b���A��_��� �<��f0*Fm~�{!L��W�N8t�+��s�!}��g����EK���%,M
S��O6�V��̋���=���a�>oB����&��>�cRΊݿ4ؕ��o����<��q!N�3�s�^j����l���WM�Qޠվ�_��������h��
`i��_��Q/�������HU_���N�p=qZ��$����w�	�`�3�5���mI?ȇŨ3��; xHܓ���0{[D.)����`�Z
��m�����0��U�@Ԧ�P_��uz��JL����8<!�⤥��E�*��2�1��N�Kh�e+A�&>C���ʥ� ��i�$��LVH�����b�ὄ\TG;�����٪4���G��Dا2�,�'��� �� �B\2�i6�#:Sv�b�^�|� J���[�,��bO+�W^0+�՜v�ˮ��3�@��12"�@�����C��D�*n]�/Cw?�x����!����H�������c����g�'�>��5g����p�1�;����a��73Q`Yh	+�%0�x����m��>0FV	����{'�[<}Ms@~��X$q�����ZN.�ke]g��'����k���/�{��n���Ⰸl|�Ər��֭�S
�>D����b��!x��x�`��'a�=C�5D�9mTEx��d��h���s/4��7��� ��C�����{��W\����;j��:ZZS�	��Z��g��m;�m����x6������m��S�qO��qlz,z�)AP�P�9���4DZ���4[a�jf啐ءa�6�"~#�"�3y�^:f���u^}(X��u?���Ř��9u�'g��N�}Xn�+��C�=C���	����<iq��'�dF^C�t��S�r��g�>��<�ԭ
��Io��Ϧ���]1��ѿd@/�ҟN��B��[w�_��v�Б�{X���Y�[~��u�����uqi����ÿ��`&�B����m����P�l�$��U6W��.����e�זG�%�oE��Idn�/r�9KM�[fE�ܩ[I��G�|�B�P�N9刏���G��� w���(�������ϽŠ����>�t�3�S��u���}��D9M���B��׾6��D�I(y����7.U�t"0�v��2�`>��$bQ��^�� ���ޚ�V�[����c��Re=��<����w%��c�%X��>�����{k*�T���	��e��H��<��A��De V����*�3��lD$�yK���l�~	�UΡ�8a�#�)o��}����٨ͦ	5G�ރT>U���Y�O�?}wS�J�	��W���N/�"�]�p�"�oҰ��`��A����ǝth�CUP�����K@�DA͑z�1���U b�
���ȁ�>P�~=�cG�@���Y��t�G�L����G6�{�n\��-�x�ʁ�ϔ�P ��/z:�`�P��H�I��˫�$�dB��K�MXv��h����X��o�Sԟ;�żc�^�Q��b�Q<��OH��f�`��U�qŞ��}����	6�7x����xn�A�!f��*8�����D]&�������N�ĨF���*o�ƧF83r�Ѧ��ϫ,���+�t�Q��_~#�h��gI�����}��q�!R^R%�>��|l�.��iB���e"*�c��n�`G��mC�2JF�!ܑL���L�o�wҷ�ĵ3��9��ԯ�yg�Ң53���1�.윏��3j�r;XbDe�|�O��Z������_�n��Z%�{�-R��`VC��n��oM��Y=�<�6΅�P��Uݽ���T���ǎ$�д�M��E���'q����q��Ri=�G6�(( ��7���*u��Wʒ��,��'�j���NÖ��g�u7�����W翩TbB_�Q!}��̤��-	�ؽI��'^�̋�W��d����2�&`�L��rSW@VP?��V�P7��}�$�һ|�dF�^1���q�n�^��&��V�
B�z�!�U���+]9��vb������
⊥��{�ml�Z�f��9�t�mR75���WV@͓dg+�l1ɱF�EsK ����p�Av����7�]�j�P�AK�c;��[R��Ƭë�^{{�y�����\6��\��՚��׭4:��O�"'o������I�4H�\�<&w�Py$"�$���C���no���{&��jjb��M`�MZ��Tv�Q��SrJ�C����OY)^0MB[C�t~!*p�ȉ���αr�������g����<E��-�$����\��#8���(��$f�l�t��7IF�a�d��S��T&�Q���^������
_�^
�GA��X�SӶ�*8��*'3� 7$�U�9w�2a\��D� �]Z�Ls3�?$p%�@�{	��bR��<>�=���	��s�D���	L�C�7u�Qڿ֌�3�6�i�!�Uظ��N2{z�̫]ͭ���7j-��d/!8W"b��,�fR|O9�K����Y:W������v�tP��,�Jcs:,����UV����Յ�&��x`0���Ζ�d"M�� ����#�6��ϥ����A�j���&AÀ�q����j��{���&<��p�S.�#3�ɊX�ߙ��[���ZoY4�>$)ɀ�g�L��d
y*�O��ŗ�&J. 먭�oE
�r'�n�A�I ���l��1��3	��`��!_�#\"�����O4x�;t%d�Zv���H�T�aC��8E �����h �f����"�t�o{3�֞���QD(R����j���] ��n)]����B�@��ڗ��Z���Z�O?���L@��b�d	e3,��<�h`��Ɇ;N�>�S�禧|	��DB��OR��s��qSm>�ңQ���!�4<<2��K%�g�5  ����&��8x`�2�4�rz��'	�����i:�4}�=�����n��@��Ebᗴ8W�\=�W�l��\BH~�¾ڇ�:���)-!�K��;+�u�F
b1k�t}ep	\���@ɴ)Ygz^C+��:��b˃`�$$���",�W�|�iD�#�-H����4�^v��6?c<�΅�;x^�i�ѝ�o����k��Iq�WH!�)W�OK��4,Ǣ�>di�w�>1q��zk�Q_O�ߧ�N^��5�W��ʳ��s$?�����I��?��b=kk��ŏ�c֓�Im��83�T`�oK@�������ϭ�� ���� ���u������3	jb4����n��,� �c�띋�<-���c��z+t%+��IE����u;����^[�Q�����S^��ǽL�47}|u������� ����`5�TZi�
�E���J���C׆w'�/���?������K�æ�\!�Uq�oD��/"oNK����1�Q���.�.;�pVH�Σ�������p�)-KApr���.;a� F�ζ�p&d��㔕0�:C!&~�0��Lj�r�
��o�5���8l��$�����+��C�ߎD���mO�4P=��&)�D&���w�Rgáݡv���TM����F��󭱒<dU3�����-�|L�wFx�@��_�Dd���M����߅Ą�׏(8�K��eh9���绣wQ!�ҽ��f��3$M`.{����6'����?�&v%��fp"��q�{��e�&��8�+���W�9*rX\��ذ����M6��:VjiF��u�KY��@G���x*{���(��o��_V����C��w���.����ۈg��f�.������_m=��θHW�	,
�Q@2�A�9,�X������B�Jg�{6�-��F�3��M�!�q�IZh�K`&�胺vԖAs^�{c@+�����1J�����Y�T@�43��ߢA�L�cͫB;ٰ=�<u.�M�'��O� ��v�哮h�Y$��N\2U�Ԁ�g�~i�����S}J���UF2�Ï&j��㋨�/Y*d��C�l%��pi/[{�F/fm	�~�hta�J:�v��cwPL��]#n�����:`���rc���~���]����0����O���Ƕ:#��7mݢ�0��=26nU�5pO��zR���6]� n�^ƌ�/"O���+�����'M�9c2W0�AY���i�������hqccn�[^G�S�9խ�+�K�H�)��,���>�T��X�Q<���Gn[�;᱄c����
d^8w�7ŭ[�ͷ���ű��GD9JGc��W�8�W%�|'
�8;���Cj�Eɖ߹ʲ�&M�!|� �G�1�h��̸:2zAfpQ�_aD�e۔`��`�\�ޚ�:z��p�$��]�w�}8)�s�b����-�[�/}�?�и ���p�k���B��!HI�'�&iM�*�	\�7o�3��,��	��A2N�HG	ɪ��.l׈�vUO�}�� Es҅;�ύJf.h;�vWn�2�A�f]"U+��q/.B���a�+4\�4�92DAdV��NH�^�y��G:�*���J����ŝ��wU�ri���4Q��t��·�y 9߭(��Bl�&%{�C���,�(��WȤ�}�4�MWi!�҃{S6pg�J*;�*`S�;]����'f����p4��-ޘ��,�㉌+Ȁ���ۨ��i��{a�l�͐RY��$�<�6ڜ�j`�e-]�+$�	�䥹�����J��K ��ײ���9��q���|E�5 R�d���O���6�cQ��Rs����j�t~/1|�+���%������2�@���
��:�?,���% G7��[&��j����	�nE�+��I��d��0�*~�cV�#����3��<����k~�~(���� ��P�����'
L�,�Wg����n|� IpkpaZ��L!7Z�IC[�{�]koC ��X��aߌ[�E-�>?Pb
܁�g5du��N��P���Z��#�E������GT��iM�����?�J�~���׍{�~��[����%"��g��rf@@�V��Pi�T�Dk]�T���ء� �C��T��B�~��vY�v`�R��W=�+���[���]|c���>���"�g��������'�ɷ[��]b"Z��b�P�6����%��7�"�?Q$��c�<��%1N	h��pc��p��b�	���c�k�m�9��g�PEic�P����oG���R�Nص,	��w����9O^���~�&L��рZ"l*�{�
�����S�%�7�n�� ��3���c��U��/kOw1!ͪ�uhQET��NC�<���
�\���I��y��t%���szƛ���@hU1���,�+�\=�r,yRz����e�lɟ�PR�	'uU����� �S���xFF�t��=�۰�����~��	��M j\$�65N�Bdv�}�4`[�[��߄� ب�zp��B2N�:��_q=w�<�n��ԟ@��g?C������D�����;
�y����HaA�G��7r���r����[<�zb���y���V�3:]h�9�I�[KF��`w��w{��[_Y�f�(Św�T(�v��K�������V��&�|��zb�!�Cr���*����@:Ԟ���H*�P�8 l)ԥ�H7# K��D�/��֋�^b8ύx�� hi���]���Z�F}��ib�٢R���G
!��:p�n������QU�����#��=N��y*�|��?�������PO�PED���>>�(�w�'��Ds_�\D����ui�hb���G�Rw���r��}#�GvV��R���cl�*�3Y��ur�y��@����Z�����������Y1� �Pk'gH_r���o��γ�ؠ&&�vl�k��]��X��r� e��,P(,�tmя�=6*�6�ڇ�m�-x���}�����$� 7F4��B�$��K-��RDu3)�I�:�|&%@=f#��kQ����y��F�!��֩j�b5�Ұ��+������=T��G*e�*}�y
���.wX���J������>�.[`V-չ�w���#o���0���"B�{D�v�:2o��D�Vq�_�%?v&$�L"/�������5T���zod~r's-��BW c?��~��36���-Qi�䪁��DM����GL�ܹh"�UrmUI�#�}�&�FT\<zzF:u?����37e�h~+x���)>mP�r��ж���Z;�$��3גu�CVBj����p����PH|W�+�0݂�9�����f"��a��j#Hq���?�lk�϶��烪(�ӭe��;wv�}��h�RG%� ���J�tKR���!�݈�L�������������8�|�9���=p�p�|��Bs�/ew����a̕k��r��
�8{����蛨��
+��85����O	ѱ��i0ْ"vk�H0/��7��-B��P�,a�9?��k?���[0y��"Nd?y¦o1�x~)4#)O� M��T�O�`k����
�0O��#m�����[����y^Ϛz�i!�.b��SFѦl�@,��z��l������|c�
O�����J����u��/���<��~E��i���a����,�������0q�9���́|U����O�r�H+tZ�ig����U�9eS2@{�+�l�xp�.ǿN)���;�^���~���ȯte�c�.06f`��S���j��?�h:�h�;`rM�y�N�{)<�܏�4<���R
vaP�CF�+�o�0�R�<�u�k��!���Sxv�X��	�h�޼��I}N� uY~?хX�>��녖��<RO���?�5��������	O��t?m2�xZPV�B�F��T0v�L���T�odЧ�:�J���=�Olշj;|�kn0l=�8.�PP�Sݰ�(}�R�B�͡'�#�r�0�Em�4�\2�/H?��'�<�$(>�,R-ϊ;�5 ��6�"�FM�,�ju��ȯM9�����?zz�&�~8�����aY.D�qd�F�|�vO��Y��X���4`U�!�[8�� oD�u���x�[���[�W��b�P9�<B<���60�C�Sh���gu��sX���Oȸo����ݰ.ι:18g���O1���(6U�$�6~����b�T!����!���4}�	�hTc� a)���qA� ��t�H�OW���гG]o�_>������x����-�R*���i'�|ɜ^�a���Ȃ�:�1&fɷ�\�x/�p���۷0~�ܙ�=@��X+��4c��1�׆����"/��(�$m��b�X����m/!�C�`0sŲoYo��3�z��?Xx�Q�&$�q�WV���d���i���2�`�4~��b�O�N�L����\rl����~�{ډZD/.����z܀ڒs�/�9�R���;��C��
"�kZ��)!�.Q[ {D�:��N�$���mG��ϫ|.�i~�GݝN`i�ɛ���9���r�����ቾF�;����NH�Y����NsZ���������B4rj�Z{�su�@�;-9������^r5�N	o��������4�tζ�E)my���~��4�>EXv'����8Yl�I[!&+3^���n��SP��5���hA��Z�w"S{XK�L�g���y	��.�5���?_4d�>���Z�P�Ps�&>��2��׽I-�\��'!��y�����$t�8t�D�UY�`
 8����C ��+��؋�ۛ��!sQ,�M����/�r�>�.��k��v��A�x��
0���,`�L��gD��EOH�o�{���=����AW<���tP�5d����T���L���0��*��6�Z@�`��n�ݭ;�� �>����Fn����2?�
9�v��� � ���m��F� o�BB��	��m@�Q�����JΙu({U��ɩ� ��>�M4������#s�fԶ�ҫ����#�b��͘�o�u��\�$_�h��Gq����>�X+!�3X[�Zk��ʂ[��2e~+�EQ.�3. {�L�ON���j;դKyw
�@�v�`�v����B����(�?��K�iN�Z�|���KƏ+/I�\�c´�=�R��[*��^;�m�q0-	��d6{���x�ZM�mY)E���l֬v� �gn�c�1�K���75���௱ˉ#mr�a���|68F)�&lpAx����&�7�B���ɩ����.��]�a,���~���qTX̍	k�3��:�I/�2=��x?r�R<��	���f������KD	���,َ\r�J�����#�s�lz��)�dl�R���x�O�7�*��7�]���/�*}AW��pO�)%�a�U���p�6�kB�r��hך@�	�q;W c2�/��
��Q�M�4@�.��)#���&F������BqR��{U��������x��-���S�ai�g���p�%^�S�<�9?n��^9��-�_���Q9v���̀|���C=��sG������P��jhA����������T����=<�)y�;k�dUҾݮ��,}�fm;��7���O��NT~?��^Fȑ���^t�T��Hj�������xBm�i���lk��dW���cY�c��D��o[�C��������3y���So>�-���ʈ[��q)�.�1Fbݐ/�6� ߢ$XSY�z�5�4�]�b�׍k�?B�B���PH�����a�Hk���d>����A	zz>�G|~X'�5�K�����\$M������E�E�~��O��'��;i5��\�uf5Ge�_H~���[��P9l��;uVM4��*#Pd�u##,w����v�C;2���j�(j==i�>b#�TlY�#Z �-��x)��`C#����&��S�W�D�y��*�@U2�v��jYஒ�+�V߅I�EC�n,�fҪ9�2���t����gv4�qG���,o����\���٧��������l!بE�^/q6K��*;?�&(m�z���Y�6CN��j�.g��j���1Ն���I��r�C�������$�l�Ҋ[�n�k�������GgYN
%�m�D����f��zs��v*���1~V���|NR5�9�ֳY8?�������7lva��L��P��-W�֠���ԯ��� ��
o��������N���NY�q��0��O��j<IӚ)�e}�n�	��1*M��)���,�^�o�+����Q��m/B�-���"7��O�l�4�l�%�.�:$V�n��OJ��	���T���ǳ�le	���P4&þ�1�Ik{m�>����������㭕I��A\�Y��謮��#��LrA$�r�D�v��G�>^�����X.c,B��#ү����w$����M�M!xIr�����C��H��T�"g]�N�%(1 ���������N�����O�&/>��
u�4��Y5<���p��.���{��צ�	6�]�Hj�8b��,�5�Q��Ѩ�h���¿�Pa���;�6�A�_���-�i�`7z>Z#�C.���8�w1g��^��48%�F�V2	m0k��<��[A�O&y���,�{�D�8���'�_{'�_��@�>׉�p���Kn�2�izw���$Ń1+|�Ŵ�,���Ab�3LϧQoY*/��Pw�F�,���٘�"�^@�'p�,�G>�p�A���u�%��ARpV�h���-V��)�M�e[�Ge�x&��*{��������Rs�q�x��3� ���@[�!,����2��~�%�M�ƝS��X��E�a��τ'S��A>K���=M� �����.ΐ��[L���hn-��?����ݹ��fU���D��) 3)�e��_gU��p�oL�0r`ٞ�o�i�_HGסdlb�p�鵣���hѬm�Hs��k󹚠��������������}PI�<�<=P�\λB����k���h�r����mIE��
O�oA߿�s��Eߝ���w��(2��obu-����F��mQ(��K<7l�I��\�m�>߽[E�c�_t��B�!\�����rm�X!�I�3�7���E�U>\���u���F��_����tm�Q<$�7�\W��Փ�%��R����Kr��v��|
��&���%��1��t�YBM1[�i��;��X����V�� ۦ��:5�Ss�u�H�l�E�P��ꔟz >��n���o�7�C�U�s����/1��V����h^]��z	���+$+����5��C	M�8ΣKE����� 0݀PU��:�$s�>��Ʌ`��gԢ� ��b�v�n�C�2��~X�nk��s�Ab�z�4�W���Gv&^� �����٠׎<��V��U8�(/���9��V۷P/��Ty�\��E��H�������:�2���uU��C���jzQ2���;�*�J�$�Ȝ�Z�Zv=d �bb%o���l�^�]���_4��Y���@�E��!�R�`z�$�-4�G�F/N��2@�T�=��C�S�<=�2[��i�j�Ej/I�	c	�b��v���\S��؟ر+� v�묗F�8����T۰��fZ{��l�{�e�|�T�&k ��
���۵��׏I��5�lT۫ M.����Ь��~`߿�����>ڡ���P\�Tg]��Z�TŔ�Z�D��K�<�����&B.c ah�SU�~g0�����e>���wO�قcJ�٬<���T��@p:�)�w��ف}�8�k�=�?�G;��/��-;��[�>^��Fr�u�euڤ��F������#Hl7��w�K�Mv�(����*Ѫ𤄹�L#�)��Зl�
����Kw�[HG���u��Q��nkigl`sg��ɲ�׉G�x��co23���d��T5��>�ca��/���l��v�/+^�@�Ӝ�ӿDuZ�ޢ�v%+7��G�P� �o'�77+���ȘvL	^n�alM���b�>���ׄ�7�-�P��٬A۝��������L"�1i>(��D�C�;t�k�_�,m��y�0�|1�������Ǆ���Ϸ	K
�J�@'��i�!��
ZU�$�*��8�'��v	=���4jI}QVl|��۠���O��v������hf�KX��z��H�v���X��Zc���������.�������*G�o0���c�Z�Lkرr��1�F��4�|mA�&�y�g|'ɩݏӺ�ՙ��0>��ɉ9���M�x���-��	�1}�(�����#
gIw #�P���۠�K�0��7�~��V^�.|��iLE�3�	!I��Gυ�؞���-$�(�t\�K�(pXg<f�1�]p��9絴��A.pc"�v����W �%Q�SF�6��h"�xjg�Ζ(!Q�<�#�	h�A�.m���2�"@�n��$<�jf�ba��qA�2~�Tb7RL�Q;��9�	�}�x��:-Y�r��G6���7�+�\�$� �C��gY�φ��.6��Oz6�R��2���b�W���ڬ�HX��Su4`^ϭ�l�d�Ft2}���Uəe�* �2�v���a��ndȚ������=�Z2��M�	s[���G�/�g�$F�މ��Г[�u���΢�j.n�Ґb�YȬ[�R������x��X��P����i,� Ch�Kn���=4%�P�v��5I*�Ơpe�I�Z'b�{%����%�:�I�C�(��_�ݥ�;�8Q8����z ��=ϣ�{��؝I�
���ө]
���2��x-�3`�[ynv�^�c�[=�X�*��1eL�,�_�NC\�ǩ'շdS�m�@�Li,R�O�	kڌ�P�]�U�JY=m��A�o�0�&�������"��f���RqN���8I���"0�
�A�[�?��m�cX9q�ջd��W�j���|Ţ��0�����mWv����q���E��wۂM�R�K.��`#if`h�U����$X�����j�s�"b��N� �7YйZ��P�^/����r]`��
=���nIn��j��X{�%;4"��	���~(�aDhO � ]�%i	��Ӻ�C��WFH+�n��*�Ԋ��d	�n��ޫ*}a�*��/ȫ�M��ܱx\��R`՗{.�=N�0��(
�D������6�������-!���m��
����H�³ր�DL69�ع>1[6��0=n+���0�L�zP6��@L�Q�*��.�R�B���=�
9P3U����<�S&�f��n
A2O��pyB�@X�V]s�O�T��A\�픏^�5g8�hi��)5�SC����j��l��#3�E� �5��25k�FB~F~=4A(�^x][a�L�{�;���Uk�����k��gS��`C@q#����ƌ��R��}-�1d#�&�D�CEDm�Dً9>�,�¶��o���{0|��h�������W�����Ĕj|�*ۀ��#(�h��ډs�"����X�S��v3z��	s�4@a��+�`����wa�U�IH2.{���5�-N5�³%1��Y���F�ԛ��U3�xT*�l�C>Q/�9$ǉ�8�MV��3\����7�i?�Y�5~[A#��y�cѝ��5��n:�:�)��̈l9�(��/�@͗�{N���#��x�n���H�m�r���83�prT3l)��u�����0����z���̞��^Ht��ǯs�Cѓ�,\�L�U��+�$�$j!��)Ͱ\.д"=���������5��ŀ������G�2?"��ݡ� ����� ������wR�- c��kO���+j��8�|�i��5;��;#ѫ?�$��`l��$w�r�'���9$G+��<.������T�`I`� ��gl.Zک.����ɳ�wE˺K�Y5���+	h���ǈ8`�v*�L̂��tWX��a/;����]0�tY_�øY����	�a����j#�RA.|�����!Xd{�RFC����ֱ,���-YBUZ_����c�����h�?�����S#�mDi���Jn
ڥ��/�|�t*u01
U�Ӱd9L��j^�c q���w�e8z Ո_�_A�������F2��
8-�����q�_W��<��h�������_����/o��L�&2��Z�ګ"�~n�S����m�ڮ����(Ŋ�70�,�Tj/E��k<��#��cB�x�o�И/$�[O_��U 1f���X���q������g&���R�Q�w��y��q�Ij�{m �l��ڠ3N�a���-9���@�� �p�kw�Σ�̪�7��g9�
7�)����c|��<�'$��M�z�x���n�D�$p�5�f���C�C�#�I�B��"�B���9�־�0��y�|���j��,����ʩ-��eRKH��Gէ��&�d35�B���KB�}u���g��[�v`�����V[2B��\)p��_@����\`�)L��Fo�����n�	��<���:�����ҰZiSǅ(�U>�O�ɰ�EO�"��%��V*�o����m�t*�X�#�S7�,aRC��l���E5���_������]����j퇋}3yX:�7� ���7mcYj7�Gx�e:j�V2V{��(N�
�j���B�6hV�Eg`��JvC[�O2H� �y$~�1¸�:��9��~��v���魥�F�_i�d��5�kK.,�=z������ʠD�����n��y��NC�(�4�r���]=A���_%�#c��<û1z��xw��Pi��S6�U4\Kz��L4}���ȫ��}���W��a6:�@|���]]9|d�����^<�U���Xx��j��}/�p[���v�qB������ܴ`��[����!�jKr������z�����A������Pڀ�t	���q?��	<|B�ǙA��ͬ�l��pa
�mo|�I$X���N;������sg<̘]���Ib {f�yY�9e��(�9{�sE�6cշ9��ؓa�� ���v�0��)�e�7��'�E���G�����iT�L�l��[��\'<+�[���U@��(�Rs�6PD���g0�GT,U��m����5�O ���em`�@ćȓ.~���.P�ޞS�C�Xo\�ȳk�p��s� �>`"����j�<}C�N=Z������ڇ�O��"yp�2�%�w���u�օ�B��,&C*�3$��D4��O�w:�9m�z�q|�E�����`'b>��`��5pM,���NG���M��L>gH|�8p�X̸,B��NU�gʶr<^ғ%:�2�������#l��r����� �ed-t���đlIK��s( ���	�
2��h�s��6[�a��a�	�
��8�S�v9�.# B �!�n��<e��}�*�I>{�6���ԓݖN�� ����E%�5�K�����0�`J15L��[�㵎0���&�p_��i�5���:��IU/]4~���V4�{RM 9+�4g5SY%�4�M���T#4{����%��!��V�AK��	��Y�R;Cy�s�T�yn�'��k<��&�%ڲ9sV�t,���nղ�4ᗽ WfS�ǝ�/�5W�,�T�q��J	�Z�W*HY�u%>��% '�I�[��.�⬅%���?��P���-U�~d��5JL�
��z(O���˰�!��i�%qGm�.8eqp���g;�Ѣg
ե��s���(����eߩ2��}!�1�6@�A� �ăk���ȩ �I%�տ��˛�5|6��~�ڬA����aCްy!��sP=(v�-AFgy��V�'`
��!����&��1��U�,�g`Ht�(���ɏ&� �g���V�`���b��[�oַ̡)��0�b�B	�����jL%p�����m���5�>�u=�º�cA������Z�p��:W?����F���}��)j���ʮ�cK2�_����l"1N������9>ܺ)�,�G���X�S:�m�6>�P��~��Hd�D)�j^��&�$O�͎�9�`���Gw��5x��]Z6�4.[��t��Ӌ��}�6g��]�w�b��>ZJ��ɔX6�umR�fG)�hf4���*$�.^�ĕ~���0,��-8�5�|ɯʏ���z�I�tY�$Y}���q/�R��)���R��v�d�[:���5���F�Y�/T�6A�����;�!�.�W��j�]q�w`����V��#�\,�O�s��������1�.�f>����\oW��H�i�R}�m��f̝ȌYn�"�m>he��v���ѩ/��l��6�,A[�YHNx�A��=)f�S^*�Ԕ�xY ���4����E\&�J��e8)��9�`�y-Q�j�$؉�	��kc��aaF��~a�݃���V@sk0�ޭ5�Z@���-�L���3P'��	S���s�9����f��2+��1��.�)ds�8��O��	G�rA�7瀏?��R�)�,~�oB���45�8�V��m����w�ᾠ�� �P�@� G�_o��h?��J���g-�V�ĭƘkUS^�&3B9Տ�����K�Ńgc�n�����n��ܜ�1T_���j��e�#�]>GS���>%���'a6��Sg9ݩ/-�BS��<���XD� �H*�'�
.�Xʆ�W�O�]�-v�^W�~eu������~��� ����o�A��Ͳ@T�amX�� �sQ4&���A�Y}�s�������F)-q!Pi���$�3�*��9n�W�%��:;��b^�n����Z�%�)���\_��y�����w��w��_��5����;q�\��Q!6׾�,�N�8�X���wl��[�L���Y��JEM�^#���~1%i�+T��K��f��!�[4�1��i����%��J�R�ْ�;U�M��;����F���枿�6n����	��[���8]$as��ظVwӽT!֣�8�z�_��
��d�������a\�m(o�������?8g�q&t���/�dPQ�k��vs���ڜ�z�S's�Cg��!_�g'ɦ��C����3���b�w�)�MoX�귝Z愞}��x���?(�=m���0�&'ҫ/&[LYH���W�@/��|��Ƶ��cx&��.���WR,���K�*���1���FO�z�t�9,:�6�E���Ky�oW��p^������T�7����Ы���'��@�'|q��)���'ץ�w�-���B�B�6�F�s�f�4��a�,�+2��T.�iZ��V� ��{u�hUI�[d��q1BWي�|��1e;��.�S������к�+��u��>�P7�#����8x�ã�"%� ʖG57��G�N��� `6����_. ��ǹ��A�G�ǳ���/��i�ͯ]^+��Ꮣ�a��}|xgK낔P�T ��J�v�M�;6�P���%�x����T�����x�.x��k%BB����X�6Ra�4��V���O(ݞ�E��d ���=0Ѵ��o�O���~���[6D_t��I�O:�W�`�Ti%�����sn��x�ㆀ�J/���~w[V�@RR�ç�pKT�1>|K䷶��I�u6�x��[�;�R.�g?2l n�E��]U<��%���b��ׂ-����х��O%j�C�?����� ����^��<�z���0�硰"u��������^�y�� �f�F�p���p�e�Y.I�@q�q@Ћz39_ 8ߕ�x�[����
?�����C/
r��kWI-d���U��AP#l䴰��՝�D��T3޲��C<k�@���!�Ŋ��Gz�����da��v��VR�#t lt��xȼb��<�\�2zLՃ�}��c	��Go^8���4��B<�'"�w���#���!�2�I����q��j�����):K�O��L_�}�����D)�e)B���?�E�6N!����g��`�:��lچ?18��W��b
(��8��&���x�Rtg�(ȭ��8B���9Т�4z�~jA�<��p�,^B˹ �i���3&����]��{y*A�l��c�'����h�O��?�D����Eg�SQ~�h��
���>��w�n,�7���c�fy
ֶ��+��� ������,!N����UPg0c������>.XH�;���N�[SU����D�O'9�(����Z��.C�ap�W�Iy���j�H���r�B�9��,u�'�jz#�X�hN���2"��VX��O(�Y�C��g��{B}V�e��&�ӕ�䪝ld�-��F��`�E.0��j?	�J�d3���7J4j�-Y	G��Yd���� �r�1]�������c�?�'��tB]�ՏKQNO]%��{�Vq�B��S�������3T}��aM��t��
_��j̲�m�%��9��t���=�de�(��y�]�0uc��|��@������\|�_��8�FeN.N��6��-p��t������	&�������q=,^"�! d������lM|���c�F��YA:��$������/�ZV��4��ڎC�!�lJ"Јصv�W��%�����C(``|�\CO�v��_�=����6y"'�i�7$yw����1�.���Sɻ�Z!r>� \��S�A1��e��hɅ��L*k+�A	�i��
��Zda�	-m�p��j-�S�����D��*l>�'ܚ`#J@�f�������<0B�(/sIzs��n�:��%��_�۸`�$~<�*�jY�@�`�X�QE�䣇�Jܹnl3��	�f�T%�-���8�J(7��H\�a��54�ۙ%��{s��r�������ˋMi������L�a��}��:�~��k���9�S�@����x~�^�+�D��/R�^5�+�Q㼖R�4h��8�u�\�ˀFGV���z��u��������aA�7M�
nΚ�l�e�mtz7O@S@���H�%*�f���O�h��d6���/"�e�hY�On�<;��"l�p7��*��G�����u#���6$���������$\;<%�e�{�H�YǈU!h0�5�뎟4;y����N�P[]>�_��' Bҷ���	Z�����2K_���$�5p&�V�5W1Y�߰8������郚�px���K����r&�X�8��mg1���K4t±,�e��J7MYۄ@�Xu�S��/��J@ Sʪ�-��I(D��pߧ��u����Z�/@���h��~@�
��ϜE����	�f��~�~���7���)=�,هd��_=!J�J����r�s����e��c�R�A��	��XV5k܍w`�����E��m1�"����(�T�ȼ���M�тHW�����İ��
HJ�ܙ$,[�U0=/J����*N��o�r�����B�{�A'��x�;�IO�}Â>�[�ż=}��MN0u���Q�j�j����� �k�v ���Bb��KUdM��1b�/4T�:m�@�@h���>uU�z4$���#C����T)�$�eͭ,&D���eJߨ#'}�<��~��1/bf�e4P�7\O��`�Y,`.��a���"�qjw�d�M�!�b�<� ܍���/�U�
�:,Ė���w��lZDVclq����L�տ�J�;B�$�Mq���ƫ-�dkcX�:�	�="x��}3�;O-ͥ&-'H�
5�D�G֒����O�2��8F%>Et����h���^@%_�(��	!�,�k��z�V���i���ܦ���2��.%B��[�zɣ+��h�&"��p�  �df����MN��5/�M(�դFlf+�1�1gg�P��R1�L�-��,�8�|H�B��TM�a����O�H�rc�R[J���>nl���,a	�L��I��-3��
Tѓ݉p-���}�� 3�a��F�(W	����u�m�.F��`#�����3��_��6{9!��~f[�	�X��wx1@`s�f�|q�a��FQm�8�'�N{S�a�"!�;��X�F���iv� R�7����c��)���p�a��(���%\�]1:�l	��;����c����Ly�Z���Dڮ��)�<ӆ�q����)� ���,
���~\~�v1��@Q?��@D5��Ni ����X�,�h���
��� �Hn�4��rT5��.*p������t�d�-O�G����H去B�2��:���.W�2/�֍�|��_����p9�a}�!kT(q���䬰��|����$���o������.5��vNb���?���͉7(��+���f:���S��G�Flq���g�i� ��N���u�X
9�ᚌ�3{M�1E�)�~V6��f�C��Ɂ'��
w��.�Q	�l�F+2�hw\%��b�įQQ��B� @&�ui�_��[zb��C�v0�B3��D�At�:��m�GL�sƺ9�	=*�����ٿ9#6�t���W�ٲIǡn��������7�@���w;��Ev[`ǌ�d�PB3����MRɠP��C�,Z��>t�1F��6�%���"��.D"��FZ�}�
�+mU0��n$7��J����_8��TW�S�nw65����{�0pϛ`�J�qau�Ќ"M�9��Cۼ�i�,YMM�27�
�pM�0���W�I
BgU�!��Ǿ��H�J v���<��Wg�߀k� ���g�ۂ�.��2~;Gʱ��E�Kp%��(s���A���D,�{�e�Q�H?H�S���1q���~>�沯�֤�/��:��Z_k*:n�{���a2wEL\y�Gp��wջXK�S���������-�|V�����8p��B��Em�z�@�Q���!��_���� ��/X���w��ђ[�*Є8��
��EjI$�I5���/:�O�kL��[�>�;,%�Vڞ�I��N��ۿ�TV����
��m�@g0�]�{��=�|Ic8 �S�<�\c=�7�PW�;ۼ�&���k7�����sٗ�S��)J��>C�'�W�
� ��f?��<��!��{�3=���,����Լ�t�_��`�Ȼ�8nB�#���L�nۡJ�Xhq��R�tM�����nd5�F[YH�ѕ�u�ID<g�~?��c�0�؝�|;�������[,��W�G�ǰ(�g��%������8�����=���]���wS�.��Z����HMy���ND\)�T�0l�Tڊ��J�`�j�mȷn��K==���>�Q��d�l`��{W�D*Uޯ�9Mu�M�>A$��!&�N$��r b�����9S$!?�Y�y?+�R.+��c��Pn��<�������'������|��{c�T������׸��tl���K�q��~�x'�a���UߕT��|Ђ��YO�~ԇ�U���.,����CB�·��2H!�xF�N�rFR#�jz�N���!�	�B��^���
W���|�\��J�8q���'%�Y �b
��?����ige���V��س�Q�'��움#��U�htx[�/������=��SQY�L��0�X'V����X�'�_Ē�io\��",n�	L:
R����zA(����.�';�b���ԃ�$BK����@5"���0�B���sӘL8,��Ud[U?��?C�S3hmD�0N���R>`0B<�:����X��)�H��3h4��cuK�^��� ^.��f��p�T�su�Y�E��RSim�t8;���nOn.�/�y�$z����&�A2��Bm���y��cw��$QJ��a�#�_�gi�a��c"�Q���Gx�K�/1���H�%p������ӧ�zUo�Ă=�R�F�G8�Rk��$m�ǳ�P �:Y��o�r.
 /G��6�L�6v�C�:�We�2�m�==k����?{&�y,�3�����oiE��ۯ�R7 GY�_����~FJ��8f)�<$"�b��&Cbn��Ag� f���$~/�w�B��s�������B�}��V��iѯn1��M��,��2�N�@푆���=!,T��p1:6�bH��7A��N�����i�yk�'�5��*���U�õ,K ��P�N�X���n�U�+�~*[�\�����b��ńEӯ3,!��j`�D�\ d;þ��~��Dx+�z}���I���mE	z��w�-Y0hbz4�c]��NB��!�2����# y/��z�nrAv>�U�ր��ʓ�*�z����Q�hX��1��C]����^���'ɷ����Q}58��1�� ^�����p?��j���P�= ����f�t���{֋��2m�e>�$\�k��ՙǄ��Nk�&���_w��w���?۱5r٥�m-�y��� P���BH^�(��)d�@�<�DO�k�0[����w�]���4�~x�������߇�j�W;O��S��g6Vp�b ᔏ�,*���BI��-|�j��p{d�"���� =ƽ�eI�
i��d|�t&1�K(	Pn*��	���~�]J�_��������CEu~�ź���b�����Lbykub��3w�(4`��lz��E��$�0,�+<�_���#[��Z��Y��T����������K��M�­(��A�UƱ���Ч�5��6AT�%�͊�ug���r˺��{mB���{?mV���˘�u��In=5	e��@��A�ɮ �Y��lҷY(�����!�=<M�, ?��q���h�9eHY�2Wސv�'��"6eԚ!-$
�D��1M"v�:��L����~��2iJ��P��s�{Â8 ��Y����8 �.5-mY��J;��x���|�*T�pg�V���ڇA3�]�y= �{!�%�u�٦��j1�7~�/5_�`�R�[5���gY�֟˼*>W��$���a9�<B�!�p���KY	������gwP�����0eaa߳�0R#9�i��|��UWߤ��tA�4J�U��G����p�`EL��T��p+���ݽ0�0���̐N-�A�� �Q�<ț8�762wp�4���F��όfr�s ���tD;7ۡ��L}֋��í��x�]E.�"�����_"f�J4�j����P���_U	%���i\�t����s�r��DT�[��\�;�?�'���S�����b�G�~� �����'8k$�`n6����F|�b�A��cʮAЎm{�C�I���VIc3.֥R�qٔ����ʝ?�1[
���`�x����Uo�,����?Q?$�o�9�@AZޑ&h
�x0>Ƹؗ�7��=&�k@7P�h/�搡�(��.�������Z�(/�+�:��^=�3|sl��Z��g��ޣ���O�)�|��P���足�
r�15�&� H�*so|'�V1z�@	�-1�	N�Q~����*�Z����uEƫڧ�%U~ٯ�p��#�pG#��$��|�E��6�*�ݗR�F��!B&&�H��H��G!������H������`������x!�̞\(�aq�6��G�NCJg
�C�5Y&>�#4u�4�o����ct���Mv��M+^�C}@���^��e,�l���ޤQ.��G$^��,�=��秊Q3���Z�J�J���񐴙�N�'F槾���ba,r���a/r����Iz�o
M�B^����i��s�Z��%#g0�m
��VO��8`�{�D�`X�KjgW��`r����#����6lS:�N��bM@һ�X$��̪�p��z�D��&�<���F�R�
���ǚ�~�5�5������P�7�
�~�- �>Mg�<��9����������ܚ�VG>j0�g�0�/\�M��?6{}{���j���xt�.���$0R?���X7��hZ��H��d_��.��9�V��B��cY^�4=�h�T	�����^p��v�^�M�0�ov�q5۟�7�x9ڡ�;��G�?�q�`��-��K�^D�K��HX���}$W���o@#��b�C3R�8�?΋����ܖ�l�(`%��WO���hhx���k�4�z�j8;��(&E
���#������:C�c��Í�����%��u]:�YF��
t�3�ё�<y�%1\;3k�Æ�M�I���a����6	��=�)�T��~���������Ί����𠢖�ڍE�UR}����J�g�-kb� sL���x�j�`A{�7��1�D��U�GL�� ����O|�3[qA�dzc'1��G����t�.��$�甍#7&���E��{a���O���󥋓O��7�_b9��Z�����R�&�O�K�n݆!�����H%��n"yˣ^�񵠞�@^�
�P���f��m>b�Ww*�?�Nq#���p̟~�+x��\n�n�O6� ���$H�Q��s���!3%�m6�C�1����iȤ�<}��:(��(c��n��ޔj�bI+o��B�>�fF|D�v��ڔ���m#JC'7�˱9�͆l%85gTR�YB��gy�O6��� ��3��Ӄ,�3��e��1X�e��n2�h墧̴�&�m�n?S�O5W��j�
�D	���DW|T�}@�k>�]FI3����~ә}tN�����1O�?���5G�<�Ǳ��QH�����M��;��Z�(m������_�
�__�����J���ŏ}�_��An6�YϘ�d�	���wm�����o$�yc�0��p��ސv%Dk����NU����~!�ǷK� $g,0Z�<m?#$_�M��o���: �6���.51Qm|0��!e��r;�H�6hۏJ'',�Cc0U�wL�j���򅘠X<�;�U�\���o���΅����[�ڬL��vٕ��陭!��K���΄����a��p��ݶ��A~%XE�{����;ИB+�(����ʖ&:It@	���	���_����Z�N|�_��oi��)QY��hL�q�����ߚ�=狕�_���|�uB)��YV��e&N�~�}dRQp��U����G�>�v�I��jM�h�Gȍe\� ���`S��b����e�>��:"�O3XDx���*ǧ�/$�,�����ݕ�-�"L��P�C�ݿ���q�S����Ɔ�cs_N�H��řюp� ����<���
h��{�J
�t��s��i��aqM��Y�Ҩ����_���  	���B%��\�s�c<i-i��*��nߦ�)d�ɢI�^{,�#Jf>`��<W��D$��b�x%�3346'�R���~6�'�N��F*[AFl7%�*Q�?Z����3�s�d1�_�ሯ{Eܖ�N?Ò�]>p9Hc{�b|K<@c��lj���AMX����vJ�'P��l��tC�����:*OR��&��Erɕ|V�·�1=dHK��!�%��l��Jẟ��f��d,�Iz<��j��	+f�����C([,�5�%��M�[!�q6t��D��?G�������yuS����	i-Ŵ�b@�V�:�7�y�	�y�x�#��*��Qklڸx�z��v_�yF�������i+����o����@�ׂa})1��
����S�����|��j��탺|�Sq_��O�w�^�ȝh���5��#�}�a,�L(ڇg��]��R����t���C����HԾ��Hɍ����ڢ���|KU�-��Cm,��%(|��_��F�?g�T`�î`�d��8/�{P1�}�Q	Qh
�Ն�� ��@2%�4p��:�@j��BT�T��Ԅ%P�g;q���~:Z��g��!g�a�d>k����G��̬���a=�0�����?�M�zԢ�?�{&���l�T�����!>�v�|������3�� ��<s�pAA~,��k
�K�с��ٷej���#��!��-��kB����#��á��.d�h�A8�N��5x���E��|�����g�&��a�D�\-C@{�DTZ#B?.EEN�cVH5�$���PC4����i�Ġ��	�9ι�H�k^�׽K!�x�
�{/뷌�Cvf����R���D::�S�ҡ�����g��MY�O����s����c�h7;"�M�qN�7�-�^re��^,<�\Œ?B~��|V�\YV�=*D{����.]S��V�(�(�2�@���.p�R�N9%�m=��ٺa���F=�vZ����2&LO�����iSC�L��w��B��Bd=���ފu�ao\�>�TP�jw�ij�jD�%���1���+����MYO6��<��P�׵,��b�%�Ӂ�v���8�V�����/l��R��W��G��;�w�����|.��G>m�yĳ*q>��uBQ[�`�9���$�h\�������� �~�ۻ���F�9'�SL�P�[���0��Qn�FA���H������";�:>#I`��J��0@�r���� ���6���zJ׍��!����
9���Z:�YƔ5)�x�S���(����Ϋw���&��4Jn���>ic?8i�������5` x-t�oC���6��n�wX����2��J�R����xr��{�恪Pլ2c�m���Ȭ멌�lέ��G�\>�o��J�+���`�t�h���5��SNNU�d:v�a���w�#E�"�z�M�<3o�ڣďAR�/R��Vk��ӿ҇���1i�v"|N|p٫��B'���������^BGn�Y���B��:��i�R-ʍp"�])PN�9pI�(�RF/�U?�n�E8M@�g�~c}(�1��2�Վ~�2�3p)��5ޔ���
��/Y�� Vr�Y���� Vy�&=ہqc0�t�����չ��~+r����)ag��G������L�͕�L�E����u�_֣���O��Ǯ��ix�_��7C+,��6��z�L��N��Jsq/ٔ5�"�۹��ULg�q,�T4��v��:{?`\����BX�p�(
G��� ���^�d{�X�ߩx�:���}����ݯI6��}�`�X��G`���u�Q����m<��s
:sʈêh"���H>v8��>*�oϋ��(������v�\���YJC���s�k��w��
�$�(}�(���O��*�TÑ�5�v��a|rǸLe���������'ߪ>p�X�5-wofp���;ܣ��̏�T�������HQ���!K��r�T6��݁���*QvW��y�
�N��.�W�4:�VgrC�płgK�T��uTL�wZ������F~�_�H��p?>�9�@<���P�,��;���n��;D�/�'+�d��	��'�$�푟&*��YG�LÛ��E�����:yp����#T<0ȸ�@m�h�q�¥U�F)a/W��������?5����sG�3W�����4s��OV%Rہ�^x�ǽ�aYj�w�=��&\ZJbBN�P���k���a���S�}|,bDrV����x�V�.; �7��F(,�<]X���s�LO�l�6W@$�\���qi�Ԍ��'u�f�ŷ�-����7��c�<g37V$+�$&�皤4�b�j`�+<_r���R:�t�jl$m�O~ � �<_��93<��̥�z\���l��*ǵ�_P�^w��X��x�FD���Ŋ�?An���`�������h�ܴ�϶]塭�K!�-���D�
 ��ai1�ΧIE��k�ۥ�3R!��
�=f� �O�m�ٔ_��P�
�J��7)�^��k+(|#���ȃ:�dj������kA�%�[��ؖ��=���N��\��|e�m�6VW��?lss`�݀c�{4-���v�i짌����MNM�)eK�c�I�8�9Nt�
��W�Y�dK?���~�*�}����ѣ�F�Q��'�.ؙ���>�/�0^�L *;�l}�ҔC h��-�� �Vt�Ҁ
I�T��mA�+*.�z��.H�0k
�x�XL��)��B����gHxtx�aj��|������p�,�t~�
R�oP�'�R��ާd� wr�N�˸�S[5��IJE��=�$�/�ׄeB�M��o�����le�Y��U#�Y_\,l�L�m.x��2-�����Y�8,2��9{��9�T��*���7��}S��I��?�{k?��8a������:�M�����s9��h�l�2;�rMG�Hʉ0���vA364���>Ŝ8v��a���lx���:p�M�L%Z$Z�5N�O�����O$�:�P?�
��U�~�T�6��	K�dzY!-ݘJ��F��)�hL���?YJhng���^���x ��mn9�BXB�so6n���:��Ļh�\��t�2��K$V�5�)�^:�Xb�F�՗� �����'��N�/��T�5��3�!P�h\9\��R,��-�6M;��D��X]���Cj:c'9+TϬ��,tf�@g+dXbh����� ��̄���_�ý@~mV��8�v�h�t��w^�Ժ������<N�?p�_z�c�)�=�Bs���!�s�u��|k��}y�HZ��<����vC��$�?��|IE[a���ȅ��(p��f��#�֜����6-�S~#�4�5��U��|O]ߤ��T�_]j�@�vE8��B�F?R�BN{K^k/l"���Ni�2ёY@���hI�����eF��D蔨�ٌh���t�&���l����(����B���S�;A�J����nn�|�!��� 3&�#�E�dE���Yp�v����{Ч�F#��l����ZDo-P�$���u�,����(&������B�;��V�<��A��"�U�K^�n��'�(;S9��s���n���om���K���I|󆭑~�W�i�立��B�J��z�(�8#����B�����m�b�VH���Mx��e5���^_�*�I��&��W�?I�i�Y��cv��c-���cn��Y��[�{XR_�ŦA+������z�?��Ip6�d�i��n�[?=xWJ.kփ���[h�<ǚS�oC���Fe�҅(��L�c���}M�,6�Z��x#*�VY�R}��yR��VJ���<�x�~4��ҳ��Kվ�͂����������3xkcr���hɁ�?HC��S5�#[�'%�#���k��b�$$|���<<n���ﾕ^��eA��ퟲ)�4KG�ZH����%QfE�MY��(���=@�ʻZN�S$�Ɯf,�W�4&�waUU��#�A.@@��\��O��<&�Sa�����n0*����1�ꁪ�C�ۆ=�����^�_����C=i9aX�O�۠\��$��"╜9�ޯůi�`M$殷���l�L9��h��F��TT@,^��o�ek�[Zr������'���u۹��N�ˀ�s�+A��	�rx��m�K�[,��PM��܉"4�jޙ�e��ۤ�����,ۆcA:|q(n��/r�٦f��(;��џ�%���Q*���E�����d@�})�6ɤ��)ʖ�u!�u��Ms9.~'�)A)		���oDK�>�@� �GO%�D�fP�E����T�34��@�`
�';y���H�\|��E��"Ԝ�54�S�m�ܙ\�(Z���-����?Z��(r;�]0�!呭z���P�ի��`�9,A�vzWK���ԓ�bb���A�Io���nLs8�׃���Ǩcs JqG�q�⦍-�-��;q�x��X�k��y�J���*��Em�1L�ʋU4����V����7mf&чع�>m����Jʲ)��U^����Z�"��H� ���jO���M�kЖ��(��A b�W:t�*n=��,^�)��a��.2��be��a���S��{�sf�:~��3$��\`5G�_�hƎ���#�jφ@�8!�S"��0��_3$RyOΉUd�|k�!���}�O4��a�f��<�ȁ4 FД^�������PH�O.��Z�$��K�X��W�o$��x=#��Gɖ���<8y����ʌ��tl��V��jC����,}M���Cj�#����q� �d�q��@�P���bô�l_����\����
(�>����Б#-Y�޷�ߚ��N�%��ȿ˫ɅM/[Rڱ�А�ڬ��eh�[��[�WֆA�@\v�
����Uj�Ф=$.[jwSՖ?,mYL�W9�䱙���R��x�N�[N>I3߹�O�O5 ��%q`�v@��}��}�ڱ��Kv�.KS�7?	���F@��.*%h�Fq�7��QJ�0� C�� P��Q�52�~����4M!c�n\�����邌M���>+��Vn���:�'��7e��W�ee����,M�W�=�bb�� �%+�S�c_��F,Ҫ2Ȑ��G��C���TQ��#�~G��C���i1��y��B}� ��މ;*|�=�8?"I>�B�� �g�A��ϩ�fh��E� �ubhN3��YN;�3+�\"�=&ԉ��s�[ride���\�@3n�=q��P���%t��a-�%��.�$��Ť�p�K�!����G���e$�L�y��bٗ<��#_ݖ	�����^�F��z��y��UxB����I�~`���Z����Q\�j���5����/5U
�Y�?�£0xP��j�n��B�_E�w�H81��P�]ƞ�����o��:(5����#��_f�cq�]������U4C�m.��X��O�xiA��\l'�?��D��D�v��R�����*��X?a��<�TSp��X]y`aO��"�!_|L�+O�6B�Ԑ�p��N��뗒��������9 ����KyJ1۷��J����W)�GĜ�m��w��FK`�6@����"��ׯ�F`6-��g$@���$��v��[���<{t������8�-�D���e?
��wq�bW�;ޜ'�R�!@�������a�YFM�w�39�q
c��Ԇ��K@�g�_
Q����<
Y��P���eY���<���~��g�B��0�Mgf����G���թh�hK�O�"�?>q&�b��q�@4i��^s��2�e%��m���:L���B�6�y�e��H�E���\l�iE�Ȏ< ��۩��d����0:�r�}���/���m�]"ޟb�L����Ih���	�g�Z�������n������
�!H *�LtH���b���� �m���m2���{�"yQ�+xP�F �#�h6�h��Q���Jk���	[�C�W�' �N[�E8=�Q�me�F��8*�y�g��i�p�j7+��_����w��k+6�Dg�{�*�7m�v�ԄA�f#�fb����`�4?v���w���T}��\��D��-�V�:�)�"7@O��i�`Y��DB���� ��L�S���wJ��3W��r�:�۶���&��ĕd�՜�f�#���|��~�7��xa�b#c&�Շug|$��������	q��� ����/,�K5��w,!�ۇB9��d/a��Aͬ����3����S`�O1#{�aihw��>�z@}�p�zNa>�r�:�b��.JRIF˲�2>�m��l�d8e���Ө����j�F�ς)xH�El"O\�Z�K��|�1�ʹ��_�v�n� ��oOK�ډ��>+x���F���n�A(�	�0��k��(�}!��ub�pDbMTn���b�?�z������{Ҋaq��wt�:ZL���7?ݤ���
*��*�J�	g��~!D����7�/b�IE�l��4U�� �_�K)��06�g�?��g�ν퍉S������E��h�Ȥk,���h�~��<�|����}9ғ0pf-���[̼C����͡Y*ySoN�����\{H~@3Zd�(��TU!Y�	��g�Jk�W� J��2x��#�'�5����}�J$z�����vSý��҈�:y��i������H��{�۫!�:�C?V��3���BY��T|T���T�m�Cz�N@�c.w��M[��,6Ӽ��5`ci�"3�N�� �7��2���z,%�dg�o���7��Xގ����ӻs��^�l��J�烾����׭TKZ����������>��OV{�~�7���81��xd@K`�B����c�cI��'j4�+V���O���§?��`���K�pC� s)��,����?��
��jo�"ĳ%,@y�&(����z@W L"�F?17�'S`��kQ˚��,�MS/�e�Z�7�u�jT�0X(��D�~j�'�������&:��{�D'�x����6�.�6=�_�	&zy�X�͞��액b]�S�����|wY�_���}�R�䏋�a�g��ç�;�B���z
���"{�	$?�}�1x�����jR��o|w}v�����F׸a�Xqt���b�:�rG���Ě�Z֖f~NĠA���{.��ғ�p�bo�
'��x�c��z� m��ܸN�84�<x�V�O��$�D���HU�^-�RC.�_���[(�л�y�i/p�:P D޻]|BU�T��:�h$�����������	U�E����#�Y�� ��.q	5�Kղ�N09�7�e�)G*%ш�Yu��Z5�C5J�iW��8X�ʋ� �y]����ѹ� ��Y����]p/=J# ��7�����E�W�F9G@�D�攗�M����w�J-�J���Fہ<�W��׹��Wu�u�;l������X3�L[�y�C�o�8��7R�	���ˌ�?l�[1��� P��_X�JE� �D`\A����� {U��˭�g�o}�P�����j�Yщ����|b�s�j��C%�O@��:�X:�Sm	3
+�"23 ǩO���P�
Ĕ�]�iB|���."T�0���-�鮏�Z���bv���T�Gw�T:?�4�kb�z<�����W����Ơꔅ���9��2��_*�"&(L)�CG����N�Wm�r�"Z=�8���bP�����x�REV��*&́
��c��~��J��+��)@Jp���C���ؗy�]?7���_�K���)ˆ~
��cK./�@������i��hE��$�Vf�%�&�/���T��C���Z���"�>�ѳ�Vi�eZ+�vBF~�1P�Bʲ�� A*z�_���7��wsl���3�X�R%���!������;i�G��W�����Z�����/����'Oj���#�Jr���}�:M�H�Β"�@���kb�V�\n�{E�8�?�+�;�	�t���[D�e�Y-�6F����*-����G�5���4���z�%)�4��������B3�,���S���o�����
�����Q�T䄦 �ge�����
�l�B�'*���d�����RS^ŉͧ${nD��o9t\��m��ȑG����5}��>c&�O˔��wdD"���b5s�\����ٴU����7�
'�kn]�ֹ6=* ��^��=�����i𥺁��1��
�p�Ca���#�y5&W³ �'�݀�4�/,f���7F��������9�*���Ij?�.�
��.��F��� �&�n|~�_]^Л�N���+�3�2�0�J���>��1�Or���f�/�HI\��ɨ{�M�Pe[�h���&��<����C�VL����������v�6�Nx̅e_u+����}{x��i��K$���:v �@e��F4�֭�,��)����Dh�0�PBA�a=�j6"ٵw�$�m��_�ki�F�΁>&�T�T��	2�������	�V>g���R�t�B����;�dօ� T#�=�$5;�~]}�W[����b�gQe/~����,�8�f�{N{����ڄ3��h����Y}�#� �d�Vŝl��H�q���O���5"�r�<?oR�WRZ� ��&�5R�X�Gכ��L�Oӆ2�0*���q����Xؔg3\j#�Aʯv�R��i���)�/�̔�
+ߋ�����GWB{<i�|� ��x]k֕�\�a^��$�U;����r7:eB�R�O(��0������N�5�rj|r�(@f�]Q<h/�B�hg���}O��g� �*"{�������wPǁ�}���ړ�'L�7����CO_�aQa�E�;ʓ!�6�W�m��=5!P���s9��u�$P�^P�:uvM�O���%��V�i��L�Yt���~����@ŀ��1��@.9����'"t{5��R��jco7���Uiy
9Q��R�5.�G�2a���P�uy�z�8 SC��XƊ�c�C&k�p�zs�S�=a�3�Jjչ�	R�ܤW5��7���ض��<�0�1A�|r5�X`0��H-�;��άu��%c�m��0���\�j�̚hߊW��5k	�iЁo~����~��5�� �as�돝�+��?#�3mS�yhtD���Mx˟B�Zl�N���s)��D>PeYC~~�*5ͻ�P�b�0�[0�ڃ
����Y�?/OB�8� �J�hͧ=�DY�������^B����Z��U��(I7����q RN��Z;>���eP-�~��h�g��JS�X� �@�-ӿ�m�`�~f%/>kv��F�|��%4��e�s����o�7�玞�b�w�Fqn���x��0��ϳ�.<�KW���E
�I4�S���E-�(Q8r��SQ��*GП]Q��1�t0p��C���W�2y棩�Pq�&���mk�*�8=ȨP�Y,�-8H��%3+�gq��4�ٿYf������$d�[_��|@�M���n��3xWUqd�6 �#����=GWͳby�+��E��=u��a���@x��)8b�я��f�����X��Je� ���U�,�Q�K����CŗƎ�h漑��m���h(%��_.��T�o��Xʡ��	W,�Mh/nP�GC5�*��q�����'����Wl��
��ۓrgk7X5�(����Wp��j�:�d;�g��S=��t������n7JX�A����2;��RNol�F�@H����jPx�a�"�ڧ�zU ��)m �G@A�	
�n��}������$*/Yİ<��&R0�p��~�� ����<��A�0��Q�Y�O�*{��46Lӡ x�1���t?Wt�L&O��O����u�-���LZ�ߜ�B9NУ�>����<*�x�h��'9�)9�� ���������5��<�;��k\�T/Z��舢Z��]bI<|��>�v��Gc�m6��ş���>���l�"7��jkb�?�d��~'V�2�* �����QZVE�	��_a��� U)�vB4>���2������Nމ�2���.8���5��­Z^aa>�����iZ�a��u���^�;�f� Y�r$8%�g�X��|�n^����7�:N�F��d�d� N�����AȓPn�C;[t|�xŋb��/�i��4�N�2@�N+4�1�Ц�O☃Syn�6������U$���?C�3�]�D�w~7Mr�Fc�R��L0�V�t��'���l���q��$���Prst^���rwBq�������m��Ɓ�f	�m'Ls�0\�xq%Ӗ�8�����%�8���'�+�" ������yb��j�(εfG/���x_R�N��ۋ���ϟ'�oc�4Ǜ�����r�hP�obz�$1����񢱟��Iz6�a�(AN����y(P�g�1whfR��_Cߪ���y���0��i�f�L5S�]H$In�q�^5��-�a�e1��^[�a�9'{���I����)��zU�#4Z��T�yq	�^c��g�3cŰ��_XDX�!d,��c����3�.׏�#�	7�@a���8��-���iEC��ih�� '�i:����NZL�H��}�_@/�̓bDac}zN����%�<�"�C9}���V$�~�Ǽ���L4��& vfi�$�]~[7o1�Wo���jyGP�~�{��~�!�ɇ�,!����ly2Z��<f/)��
�oOx�V���/rhl'J��:8-�F� }��!��jt˼^ ������v�I+�ghܶ�h�p�����p���e�#�L�������d�D_�~�%�*�I�+LM|S[LSh�C�Q7�#�"�;L��r��Bo��7�d���٪I�o�����`MV6�y_��i^���K���x.���p��0$�|6\��k�s�k��-
�[��|�YZ��]̍W+�X���E͆�)��i5��['2��|ϳH_�"@�`j�3�-!ET���<�v�!�7 �L���]��Aq��R��e�.��M�4���f{��W���]��nb߰PZp���ߌ;G#���yo_�!�y�Q��"��}���)I�"N�{��=����i�>\��v
.�!dܙ[���k������s9�_gߵ�� 	v���>4"�4A��[���C���x��n��^\]����N9��v1H#界<�eM^�;Cw��p"�7䢷-!Rv�=�G�Ew��SF����!9��B�a��^JΥp�fMz��/���e�P�Yx+9jX��0�c F��~���*�[;�+8~B#�i����T�?�	��E?�#9h�C���\����t�Q�����Ls��,�����z�m(3O�}Rl[�<�"�O�*��a��)ǫJw1��ͽ���I��>��P�Td���U��⽢�x����>�{o���g�>�8*�s��,�v����J�m�)�IhA���_��%�n'��½ڐ����.���,�S�,�����s��>-���������
�y+�>���MN	-~�$��!�Xv{^9q
�<\weEWh�����)~��qZ �Q�J�̂Hՠ�2#�m&��9�e����+��r�;����u�	���"a�wAa��ɞ�j�9����O�q%{������Vo>@��4�ׅe�Y���.��=nõ���
�\�3�w��P@�� Ph�)n*�P|5��V�ˈ���:'��]we��&8J0��z��#z6��=h�a�\�c��_�Kz�b��kj5\�ې_���ܳ�7�]�%?72M�'e&�a��|joq�3�<�&�4i�k�F���M��YQxX7�F��x7��3������]�$ Y�v�;��P.X�������f��$��_��|i�`�/�3g��̓F�-���4Y�c�3�n�bۇq����{)(`_�	2	𴓘��P�W$�ba�*��(������)tIG�<;A�)�*^<�u�,�e�ᰗ �fky��J	�R�q�#���	�j�-)d�3L���⑻�*��tՅ�W�u���IH�T����w�V���]����)|gT�*<�١���0��OGe�YQ������A�z���Ʃ��j9A��!EZ��|Ξ|뭜M�A�^F,�D�́�?��דBr��9���׀�v�!��,8�6�{.�[fm��g�2�X*��t�C��y	�a�{��� �x;oU������l���|��Hn^ٴQ�����o��T��+����� {겧S��5�u�<7�tڊY5o��sBR���'W����_���o����X+]�=E��}ο*Rs"1��\��(0Δ�:�ۜ䦽v��oS��P�q�ġ�7�;�H��[�:2�@�Y_t#:��ݥ��i�3��c�?ʽT�e�Ҵ4��:FX7�gF�	��M��)0� ��W!�4Mo�DNRS��/���&�
�+2b���M§���8*������4������Sվ?�-��Ǐt�}��>l�iu�Z�T��%k�a����93L�=�>���-�g�#��g�Aty�]����T�0�W����Ui���`L!������6jg��/w_,P�
�\jd�@אe�肠40x���mW�Dk����sW�"o���KM��}���уX��^��8�F��7�<t�C��v�h����	��`�����`���j�����*x��O��iO3K���)dw�|��=���%-��J��3i,Sd��� C�=(O2^�ׅ�9M�� ���H�S|$l�Yb�Z_V������t{�x'�J��U]��e:.D~?�
(D`�-J}훥�̏u���w|�>eCe֖�E

�Q[z��=.$�G�Pu;�9�U�W����)L�L�C��x�(Q��Sl}����xѳ� �O�0	����r�����
��^����]�3%�ph��W<n��X�d�*��籰����)�ǀp��*<��ߥ�6*Gb������A�CQ�Ew-�������J���:��9���Z��zX���u�ۤIwί��@��2k������(Ga�e*���"ԉ6Y�H��@�N|�Ʃ#?|�t����A*�������g�q�X��(����/�� ��-��J3�7.&��b�o s�[���]2X*h��Ɔ��<��T8�[d����Փs��g�:���L6?Ÿ�?G��б��y�`���uq�1�?H刜����K���}��<�7\9X#/�}��n�EB�/��-< M �:x�zG�
�V��?ZN��m*W���t�8?̋9�k����گD[WTѶU�F��X�5N9�$O�@{J`l�x�G�|�p��\t�e̪x:��}���%����\��'�E{���N8���G�p�<����5'��-5�g���D8ݥ��T��hd��T(���2����.����uJ{�D��9X�7��E�"������3|�=}���%�ڥ��\O��i���<a[�B�Z����P��� l��p!;�f��ʡ�ګ��)�7*��)�3.Ş�A�� F�EN]f�y�⫕�ɱ�(��@5��]X9k��z%栭ۿ�qU��(�Py��i���Fʈ4vY�q|'Zڒ %U��op�\�������3���U��hAb����Z!�0��Ǜ�x�����N�7�U��[ �K�?o���i7�5i�\�˝*%��:b���e�jx��b̧�ʕ�e�D�@7 �N@�z���Ж��!r�a�Bu��e�'5���.Ռ��7�1e�L�:�c.�yfrW�u4��w�i�-W^���U�_���c	���	��g�%�_H$Wюn�}��6s��H4(�.�C*�d4&ٽ΍q�I���32A|�Qi,Y^�G>�+ڃ+ܹ�����+[���8O���o��w�w�*-�R��vb�dA���������x�Q�%&����N6I��[�~?G�r��w�a~n�5a��}�ve&�P�s���vK��mf�w'��h���a�܂?���2���K)�G���kt��EHa�!Sj��H�U��bC��#��f�OIB�3A�m���Y*"�0h��x����j,��b�1�d�˹m<MM��9c�����`��){�8ce��3���V�r��U[�Y��2~�=B�T�k�̈��q�@`U�I�������ᛗD1�|#
;iq25���>�˓��m5�u"�b|A!ƕw��7g�n��B���o���E3I���n����@"��l��G�ʗ0ކ.��1��i�u�lSz������i�梂~9u�;�R�ȸ|׷�A�bE���}�_�,�&�@F�_��t����2�<専���V�P^����d���� �u3s�;+k�^>S�h�+�7�M��ꤊ����l��?4�L�8m�yd+7qU���tG;��`�(Ef(����K6�Q��Dp�ۑ�A�_7rf#Pi�LƕS�dh+��ص��co&LA�eT�;�ƶ�&gB��D�?76�i,�ͣ㯉/g��p-���������,���G����$��+	]���u��\����,����v������ ��)��d��n�`�.PѧY������w0�+���N�Ji�!�p�2H� o�a+�'�|v}>�i�XB�a�+c��u������ǺMP� �א(�KramJ��9/�{��韶�U��F6ZJq@9�)yIu�h�p�6��

Fa���묣ƅDl6T��eT����T�o�JLG���� �����n1�oK�#�_	�Y���S�o�G��޹nH*�?�r7�wQ��M�g�[��mU� 
 ��Ҍ	VQ�/�,�Ε0��U�+��./��E*�P�K�h��ϊ�2`����5B�����~@��be��(�deG�O�qsz��Jrjr�ԝ����ً2,}�j��e�T"���1�'�=?��^L��bL�߻��`
w���vjܴ�D+[c��9�-�&\��A/��`��F����`��;ʹ�(̘��v�K=��v�.���yto]��*��xi8-D��.2�K8yJ=?t9�"�@�`�6-q~��=3�� �]����(va���rib�o���$�|���)�,��l��=��!j�]g`���#sp������Xa�y���d=��
Q�TM��/���i�R��~%X�}>DH�w:c"�و,�%$W��|�NaQɃ��p�A�E)Q�k�F���jh ���I�ڔp\�v�����/��K�z��f��2���A���s)��oA�d�	�ș-�V���X$������W�S�xHAS,��� 㯳壚�3��	զ�V ~3��$����"Xゴ%*�����[����
 �pzۊ�4g����Ɗّ9���ޝ�!-��`����y�J?�l���ʟ������Nۭ|6Msnr�9�⿢_
L��Q`��&ۙ�ڄ�����8e�#EC���CǓhx�O���q��q��ZجW@l|�Vr��c�'�����nf�WX�@���������;)���/�X��%s��a$��(I�J��do�V+�07z�ǒ��{	H�D�C��@��b�* ��7`
N̝����ؒ�����\���{y�����:�%�E� �eRlk���&[(}��6w�F->����w���X'-=��m\��b;�Y��xx[��k8j��Q��YV`k�� �S	��(��鄝G�P:��jM.Q���^x���)�N�דD4=u|���e��y���"�hb4��y�!>w���I�}���nQ�z�[�R�[>���A8�HQD��w�C���q�`�Qv�.p��2dF�����͋�<K�.��
�DS�w�����e�pC�}��i!�˓��tYo-���O�eQKm�@mD|0\�g�˻�h�eWh���� W�ӆ�h�}��u����[Y+�rMH
=�"��
M��ݳ��%�����ޠ��ل�,��S8�����1��x�����~�L�V�A%~,׫֔�$FꤏP,b��<m�R�eU��tG��� ��?���GO	�*��<�|T	��yp��I4�N�~޺���Z7��o��a���8A	�J��^�ʧ��p���ˍ^��F����#
�6�U�jCs��q~E��<,��}ˤ�n�>��9�ݹ"z�����r�f��ًێE��T+֯F
t�z��x/Υ˳�F�E[�1�F�wZ4
��\��%��Cy:-�$!�}�\S擬��6�cSg�P�]��gͲ�jR�?��c"/�F&)���E(⠝��z�뜖��Z���~�:$9VT�q6>��h�ֲքSO�yG1���n/7�g��h�.���4�-�V�����.~I��<m��
<���9��A��eqP�8ܥc�*_eL9a�FW�ғc�T�>-��+ٵ�)I���i�	m������5An�jP6��W)�D�L�+ҥ�7��$�-�:1�,��?ֱ���ʿ���	@O뱜�?��'�*�E���Z���O�f�^��7�Q���Fn�8��vXׄꘟ�}�\�*l�cz�%�49�&׾�w_c֗�;�5�����s����H��dc�b\��{c,	� �G��1��Ei���h�ޡ�1��}Fj�3]��)��<c,�+�kB����*���.v �?�{�՞����yY�.�����f淁�f��bEt�������r"o�Z)�t�~�bw�Ywɤ�dr̸�ZK�9HȸS�C<^����
����^[��A '�_r�I������E�$�C u��@�+���q�p�D�������0��5�SQ+Ů�o��V��V��]��v�U?@)�ȅ����*�&�9��m�:�</�\8�L��"�;���Xy������}Y'[����hq@������E7N��p"�#ua��
{���Uo�+��`���&=����\g�$��)O�p��X�_c�{w�m�1�;q+�w�v��2��ly��$���-�{Ʒ��Lz<��bH3dg:e+�^¿C8�.T�x��f��A�}/�}��q6M��~�-j��ٛ��;�s�J��*hY�9�����䍃|���ӕ^k����R+[1�؅�=�%4�>�����LQÁw��v�����I��=I�dY Q1�y�+~�UU���ʌ�B��Z���?��7�E�?q�"��sʒ�.V+})�P��B�5̦��Jx�ΜK+��E4p*�aqN�O2O�lYS�Tp�ğ �������z��4{�aDٸΪ�Cl�G�@XZ�(��،@H�	���0�v�kj�sy���i��^�S�1g�?
 f!�#2/�L=X!֡��8�1;A�ns2�1jt��6��g���5���Bu�Ay#ÊK���E<pe��L�?��c&�<ӈD�O��$X"���`��B�E��y���~���w䙡u�0t�K����a�A-���b88�<�5٥�h�_����Ɨ���^�/�m'�E�וS�֬e�0	������Ո/���O��&'�%�����m.��ې�+�^8�z�/CO�K��)�~��p��Cx�G��;�����: ~!����Z���^YO��*�٫SKn By�����>Rp���3P�^�����;���AA��V2��������`�_�9P�Fe� &1�i=�R���E��ߙ��Sj��'���aM.4���y5�{��G��z��N�+�3�=�ʲL��(;�����34�I)�:]�hᰈ��P�[����̆�@���d�gM��G�Y�֯ �m�Y<.�|
q�֑��߹���)���Od�`ikN3O�Y���������E�����������)c�E�Ȫ��\v��i5���N��w�aNrk`�!9W��u�z<�A�T�>�u�Zǹ�=	���]�!k��.*��J��+�4r����9�"č�_G��> �#���S�͓��R���ѩ[�
������؛�����MW�J��$>�}Nj��1��`8Ǟ�� k%0����A+�+os�%��rj��X}r\�.+fd4>]\����&�7��%^�]/�GtKq�gB	�p�K�aK��A/����JR2���o8��<��i�b0�����g������Sk!ja�C�1]}W��Y�Eu�
o�1�^&�K{�LmOy���$�}�,��|����>�\wI��|�-9a�n��)�tt8���޽ElG4|�)����g�+�,�nH����;�Ҳ����S�����8�'Ȕ_A��/�dJP�Lz7@j0?s��6���%Y��� ���Kl�t=��N�D�6k?sC��g%��y����*�O�=�BQ�R���_5^P�y9Y�{k<X��awR�H��{�j;�@)�Q㽩���9���d��H�NN��,��Ub9�i�[o)�N^�M�̶w����@���Mg��U�J�W���boP=��
v֧7���^ ���Z?в�MH-Պ���P�Ph�ݿ�`$*�/��|�4t�������,��b��r��9l��ZUm����W��	�s����Sߩ/d^�����A�%��yP?ؔ�Z�{\V�!�Z/�j�X��s\���u����e
��;�a_l�D���Vu��v�N�[\W���,�;]���b�9���p��:�H�V��F��*7��s6u/�o�S���lC�'̺9�A{�Ͻ&��6�����n؜�6���5JN�t,S||
�)_(༂!<WC�ϒ���^��e?]�7���z�a��� t�� _+�j�0ć�v��%�7��B�����|ܳ콋�W�z�9$�Dǎ$xԈ��)���yh��z"� ���^���ߏA�lǵ:�ޞ���JД��@]�pLǋu q"���y �����'>V�#~94X������O����4����^X)���L����E�ktH�df�(�|�܍���R���:�C;OF�8��2)	e�"}�'
	gE�K�~s��146������+��L	�,�����<���R�5O����oS��yc59�޻YܞX�a�s��(�Zp�ݡ"<��P��g
鞶so�za���]L�?S�������N|YT�Y��E[��q�>�_v�
�~��{�<\$��X��*�j�0jI]ͻfa�������蒜�mt@s�9�}�ɗ%B��l$��D��-�Oa�G�ę�`�NO�1T�j�.�[�{�D/�H�)�L����3E�-G__V�ڔyB���)�ȃv6���T��Z����O����|;�zeӦS8YH���/�Mi���8�8���	�*��zt�|��4>}1���FS!�4UHVk��������Ю����D��	W@w�@�e�iEk�L����8>^ �|�������fw���6*�\��.�+NOz��}zU���m�h��&��Po
-�S#N������k�J1+���U��6)uK/�/(�b+zF{�E~�pJ'�07�~�ܑ���[�o��i�Qt&
E<�^�zm�����i+f� Vf�=�����G�ڠ�x?��X]�b�K�Ku�P祫R).��ѿ���=���~�����ɾ����o#cu|wvO^z�h�y vR��Q�FybK]�f�B������$�|=���ke�O��Y�\�]<�S�U(;m�e+�ޒ��0�l�3X7I�����b}�mos�	���H��r���\5�qe��a&��:�5����;G����pI���#�i�#�/mu����BS*��o��zc`�>t���i�I=$�NBzx�� ��}���L岾9���ޒ2�����5��@�ܑNdi��ﴬɓ$!Ԓ�`��)VL��FĖ@��OLd��Ӝݾ��.9������V�,�ʗ�^-��;�tGp�F��y��b�~s����p
�i�����zMW@ٻ��dp�0%���'m�綿�G�A��]`��`�~"sWח_��"�B��֖ 5l���~��g��K�$�s�&�Y�T��*�X�p%��#7���;9�{���I����?��No��G@����
c}�6i�=t���Q���@z:d���]C�Í������B�^��PS3�޹�(�F&.��;[��#�y���oS�v���ۯQ+~O�m:P��4�%���ᶠ�ܖD�H�9o�Tyb[e�� �w�>DO>�����p����@Yt~?x[R@2/�����[%a�6��J�g��E���#���q�c��ʣ��m�9_C�B��.�D�ǎ�Ka��z����o5�%�d�=Tkkv��li�(��!�_=b�P7J>��4z� cZ�L9�A��q���N�`�yMY(k��Y��@��(����7sy�*�R*zZ������̞��us�������w��9g��h<�͊�&���A8�Q1f4�tW�GȎ1Y�ѩ,������S���gdf�%7��`:V/f��
�]b�њr���FA�tF��ԉ�/��l�X@��	��/�̢�eF��͞zs�+uK,UB��i���"	�룼,��m�8��I]��	m ��IWO�l��p�scAW�	@W���@m���'�]tQ�|��V$RK�v�,dɟO����Ĵ��rcg�uGQl۔�)�:/�5G��ʵv��?�3�1a�b�����,9�D@T�w.���6"�DL$u�Q4PU�a �2���S
OC�t�ĉ�6���Q����}��y���DV�П��^��+ߚ�\s�iu�%�>ڿ�	�k��{�b�Zj�m��Z�X�`$��\z��&iw��2��:�;5��[z@Tʣ�p!:��(�ֆ=,�+���~�UM�_�����*x{o��ڽ8R��?<����4&d�桹QU�7�5���7GW̿��7���y۹p	���>�m��չT)§J]�ߔ�H��2���|"���(פze��/����\
�Bͅ_ǚ��PEZ�KeC��fP��cֽmz!�	�H��$��w�
������H�#l~�|5�hU��H��!��W-ؖ7��zO	�m�yYk4�����)�ES˹�2h���!VE����]_���Iam�p2g܉��.�����Б�P�9���1�D��lWG�s�O��ԯ�8���ʒot��s��[@���[��U7^�0��Jn�3- )���c�d���Ɍ��g�L}�����g�ưX��q)y2y�����o�]'k��js��	|�kϘwzL�?��H]c{u�~�#BKguc�>���24���á���0x���¡Lp��s����=)W�(7U=��]٨ZP�*������%L=�s7)׺ 	&��R��/�Ly���.�J��1��mFp_�i�E=,-?udJAe"HE!qư����~g�e@\��8�';Oh���\u�{P�(B^�>6X,�t�]b� r?F����Q��D�b[��Js�?�5��ꆦ�[�ID�k�C���ӌ�������bʰ� ��pVpCG�*��z��4m����(I!����)P(��_��� �+���܉W���O}�'��@^��B},$GM�"��P #�����e�A��_�WO4��3���6%�P�C�\�T�6v��iޤ���I������M����"f|~1]}�퀨�&T;ˋ���;�H�%��K.�D7������"gO9 �K�T<����y��Yt�jӥ�O�/H��	���et��0�c&b5m�O�O��<��d�A 	^$���}���\G�©����-v|�{i�Yʾ�o��w9�R���Z����ʭPn���j��eLT�����_Z�!����!a��q��?T�C$w~fDW���v�p���%~ӡ��w����t��D�1�7ppV�b)�j��bZ-X]�iph�C��V��*é��"p ��,TØ"�'0���.C���3�&���Iʄ�6�(f�6<9����<�	R���
�>$B�(xM�dƕ�F�(�#�!Z� K��~��3�Q���mY��#��~�@��gkSX;�r�ћh<�GL��ۄ��"
<8�{��7��w�1��0�����:&Z��i��~��Ϡ<��݇�#�j�{U�C/��m6����X����zO��_I��<�)xӔg�|�N�Z�$�hc%%��Ѩ׏6Q��gbUw�3�5��7t+��@��U�YgI�У<����2�N�g��)LPwAhdO�{�*�I!Xi�v��F~ ������`��I�y�ӳ쯧N�\8t�uf..��uۅ���KW\�X�V��N�/���1�` �yIO�G���AQ�-2�͇�=EV�Aba����ǺGq���Mj���xU�|P�'mC�����v
4�Qy��Z`��,��Fz�mIN"���YyC�P%r���$��,��+���i���'{۪�N#HnQ)օyG�oa*����~�p��X���М���n�ܫ�쮔��Q9l���ʶr)����U�w�QH�N���Q��������2y�xB@���y0� �J�&�̍em�pm�\ZH9�v��9��թ�(�Q ��1�OHF�(�g-�����ٱ��Փ�J	����k0oq��u�>��h���xl/�q�;��'���� .����������O�/]��!������5�-~YILA�Ze�_�Y�`�~Hxݽ��U�T[����q*_K�Qn��(�o��Eb}��*z��Z���4�U0/�k��H��1c>J�p�En�#�S���(��R�W�������B��pl� (kX�ݞB�)�u�EjH�А�P�|���ae}0QM�݉�C���ƨ&2�
\�H��f>��к���[���E�6�II6��ɍ.��hU5ܻ(wjgu��i9�45��wI���h��=Fi
s�G�jzDv�l~��=/�Wz�!�Z�	n�u����r1���w����6���̟?�!��X�}+�8H�f�U�{=�����Ի���2sJ�.V���vS\���[�o�9�7���Y<�}�5�yŘ�RYͽ/h�¸�@[��l����ȹ|���U.#C}dlv�(ɵ���7��BB���M�B/]E��qT��K�7���Ez� �(G�o�<�Sؼ}��1��Q���:��|������
�!m�
g��j��QT�0�OJ��F%3,����yR*����wR°���6��#����e#�b�>ic��w��N,���	lr�{�C�繉��1������/�Կ?��Z�B���t����
9;=�� ��x)OU�`gҽ�#Yꈻ=v��w4�R
z��N��~��ޙk��	�9?c[�>�EDSb��!���L��?�q���7��K s�r���}��$0�c�,�5i۸=`Мi�#M�h�g���^��Q]Y��#e,�,oO����Z:�21Y��Ha��E�
�"�wfA���rر$��x/�ͼ��p�ޚ]�WȎ�&�2�BV-[�~(E+�ޫoo}e)N��N��
(��&�1J��&���6EY�)��1טK?�J�)c	>���}���P;>X����HŅI�8�L�v豪���K&����ٜ�P: �
q���	���{����_x	*�dI��>5z�V�� 
ԅ�1"��Wh2��h�Ƭn�{�����.|!���nS\��>�j�m�
9$�<&�ރ�XGc b�;�|,������էx~���{�I��X�wT����?`�LW8���*$flற3�`���!�Lkk�q4�X�79bQ����]Q|v�P�K��Z#���t��b�fi��߂90n�<oA����ҫ���Ҙ���:��{�AQ�E������v>Β9ua�ĸ6({:di6�r"��^vɚ���Uy<��Q��#ك<�p2��ꭥ ��EP>Ѓ�Vȁ�^���d�+.�S�,~� E��|���?�^������d.H!5;��������8KHs�i��/�;���Ow{|�B�����[.��F�VE�1�T�������!)D�����T�����cG3{�~,�b�G��ב�����W��qq];���o�;�"����5��g��f�v�
	���A�Yў���ٶG�5:ˠ=�b���v��uo��W~��f���z�k�E�Ѓ��L�[�����μ�=n��>���\BZ�M=;կX��ݙW��������U�A�oU�t��a[�߶�.��~�*��f	�o9f��N%�����rq����]enh�����r�E0���-}�Y K�$�^t�@�Z��]�癆9^c{L6�/�0YAOf��n�V�9#���Oi��>�q|��8���_d��	-Q�_7���؍�#Pk{𒂗��ݩ�Ƀ	񱝝�yv۬��zb�'���;���
49����"��83C��T~������f�;�繇��I���F|Zx���&$z�h��^�`��:���'!~#r}���;}�:ϜQ=�_X�r6���8H�D}�.��fR���\.v+)b�Q���f�ܵB�~�,��t��~^y"ܘI;�a*%6��kl�K�O �o�m�%?����h��O����3hU�`,> 5�: �<�[d�������X֔�ĳ΁ϝd	+��J}�:�<���Qm�	��������a�m�-���^�!O��좜��N�M�zQ�CZ�J�VH;U��E�3�����1z�֢HHsYᵇ��]	@!y����i���4Й~���S��.�v�M�����~��YM-}��@��2�ji��j�u!��M�Cw�i���Q1�[�_i��3_s�=7J�9��I�?D�xA���0N ;�$F��z�������leY��/~[
���ӡ�'L�����β̆�u^:������[Q,#Y*m�j��R���}s������a|1T���/L"��0�9����@�9;z�?�u��C=1&���4c�*����!��9:&|��f_��ns��)��M
�xC�o���䢱ƈ��@�������D��2�y���lE��r�u�R��9����	��[IݱS�P�����E2!D}�c�Lf�E��y��<���W��-r���}��� .i����ŻkD��l�����\e�#����x��c��6��2ô
Y�߾�m�^�S.N�X����W�\��~1a��v~���,-*K�WG^�}����B�qv�w>�B���~i����hr-۟B�ݪ�� �sm�3b�`�JD�����]��Ͱ�I�< u{	���i�sSE��8���:2�Փc�|iy�] *������޳�0�MO@R(�`�x��H8n�'}�m���zSP`e])7h��Y
#�k��K|���G�r+�;���`*���"��*N�4�Ղ��J þP(�$�r'��X<��ᖸ�s1L�w2:"�7�v�dy�^��g"�&����n�K;;L�u6��TK��}u�UM��N JF�37+������9n<���w{o�x�<�����l�%�w!�iᎅe�����.������?:/���J� Y���@=�`��@�J͑�%A��\B���x�)fa�T��0-c�\`E����P1�RSo	��qq����r���4k_��U[G����ǅ����)�����p����S������ɑꤦz��]��MnnN#�_z&U�u���9d)����0�r�q������3��_�����pHZ\����3����2�E+$��xt��G"'��(�\>·��YB��[~�L��6F���t?�@���)l�����cM��Y��f��B��辏Q��/��=<sЮ�$�<�Z�S���@��#J0��[s�8Mwvy*�������s�a'0�P�P֎�k�(��~fY��4w�Y���}��L
4C�wj6L{�O�n��ǎ���b�?��?��D��p��6�k�x���Pu�����@���K��@�Œz�G��Rk�jl����X��^�LȌo6:�<~;�u*(�C�1E`m��G5�W7�H����
���9��9��lie���
l��3BC)�]*mDb�"+�|=Z>K+��zG�f�^��]�YB���2�E����K�Q!���	��0{�,�x�\q6W�Ϝ��e��Z]��>	�-��׋���c�RJ���S C������6�s�+��&OoЫw@��nB;z��!d�<�@�(4tT���|k�ƾ�M���tO�Ѕ.@m�Y�?� �c�|ȭz��%�����P��r�u|�R��T��C�l����d�^j�P�q���ΘF�wk+?�������>��Vd��
�iê ��6-����	�@Zt��
�za�iď�_6������ �hƻ�����V/딋���&��~�;|-�iӉ�;����z3����4��Sq"�U��$IBpl�0����k���ma�9$�[7��>ԑ��
�s�!	��أPc������ܖwc�FMP˽e�E��*w~�!���,5�AD�;�q4�OӐT����"8�gU�P b��51.xb1�*`��	2Ճ��*�
ާ5��c���@9�j9����b�A�-h��[��`De��������/���� ��Y���p24���L��6�0�^r�h�ap�/^�sۘ9Q�b;P�� y.+�-�9�y���i�t%�a{��+>�r��.�G֖��s�d
�-��Pm�&Ȱ1������Z�����\7�I��:3,�y
o�.���Ѵ&0�2
��[�6��a���P�3���l�8E�]Y�j����[�J�Ί���3�󭌮m��R�53��|q���������6b�!j����lg���@��l�{�P��ۃl�6�8C��o��0���_�����ͷ#f�mL�����A}Ǳ/:vl�<l�(d�$J��a����	_��j�-3�����:<_�]h/�X;E��T`�+��<�+ɺ�aj9�<��/�4��6���Y̘Ua���{��&�6y�)(��.�Y���Rq���^�Ucer��g���"�J������fN�~o�����~`��.��DeE��6�N>�?8�Ā���H4H&��� ��M5���"�e&�0e��.�h��z����XP��%FX��<3�����)�5���s��'E��֮�\����v��6U�Y���n�GyAn�M��6<e�w��Zet�:��<T�4�|T͔0@E�Œ�	��4��o.�X�\�����lT4����U�7��vr�2�R7��r�k|��.���cux��xƗ�w��xi���4&��3m�q�t��[���}�l֥�R�����#2M�U�5�+in����D�x�.���@kF J��:W�����|"�����5���dD�u�]�l�����	1fh_��j/��l^���| Z�&4�O0!�����ǡ%��Ü�X�m?��:�E�Iz��;��m7�p�Ds2�"�m���ݸ����Svi�ۆ��=�%8ܨ�X��R�x��m�J�F��F�]�H5����=F��؄W9W�r�/���Z%L7aG��Ǵf"����&ھT����c�����]6O*��ǚYm��!!@��+WEN�?�b� ��FD͎H�X"����p��^�C�O���RK��X;���(D�����B��-�����;�_72��&@�u�J~�t��UG�����0[M�v��M�W�#8kFZ��{ee',[��E�ڐ�
ف�7X �F$rCή����!��G0�v:�O�[���BzgFu����+�c���}���0 �����t<8oL�í�@vE�!��;�6����Ti���{�Q@.X0v�Y�Ld���?�6��
g�L���i_����(�E7��{���4}�R���6��`pn���@5ų���-$�L|����lH�ݛW�T=-�{>{�nO <������� �i�>�R��Jś��w7O��u��&�椑�˞O�XW7Z�#��B�'�5|��c�C9-r�f��S����V�2y��H��ז����[#G&��PNV$�v9����2t�x+~�3��~�C+�%�xA���@��V�F+aM�SO"Yο_�0d�������QD�iڃ�����fN�-�I}�͜�`�`%�aL)���_��w��8]���o�9
����]��`��G)�P�}Y���OJ���~}8������f9�l�����2;�O������H*�>6t�E-v��QĈ|
��}z�H#�=��Պ�Z�L�@��躪���F��e���g�4ĕ��̍����*-D��H�����eO�W�{��{��������yS��ti���s��R�����],��,%JJ��4�7��eu�G���A������A�X��O/��35�h�y$=%�G�'�j��ijΆQ�ie�Ź��(ai߰��3`U�VT-E�P�b�v�p^ޟ�F���/�4�M���Օ���G����|2˭h���7.�F�$�=���c����c(��27���X�	��
���O���<�9A�'
�hP&��J�q�1��tE�����R7��RV�3E�a�xy2�2���
(��J����+XdTa��/==�S0����]׸S�Ȣ��+��3��Bh�}e�ݍ1�K��s�������N.�l&p��E�{�]|iՈ�@���b�F����U��g#�|i�wF�����\[]�8¸��G�=��������{�v��;?��{pBՂ0����<Jm�r���0�Tdw�#V����ڴ�!��؆�
ZN�`�ݍ)[8Uq�J���s��r 9T;���C��Dy��*\��~�i��J��^x]�rǙD<�F�����I��zN�/z�e��ƻV�Ϟ�Y崘˭�hP8��#CaP��Is\UF�i_|�I2��u#As�6K��[r�j���ȆC^�r��`P�<x�W��V`)���R�A�bx!� .��JӇ�A��XJ�wY��	M�����6��`�`�(�5d�XW��(��~��,�߽���l�Q�58-%��P00J�g+jȉw�D.NcC!��~����-�j�-�����t"�s8��J�i�,��n�Kͦ)�L\%�Q��-g\@���u�ݢ�4�'[4F!��@5�6qbӺ���n��UD{p����]�}���v�C��I}(����Ej���|�����%"�Q0)���<����';�ᓲn�y&��b�>�0�܋��ob7�`�Q��[�rr�R3��,�ő��u`�ҏ�{,�ѸZ�,0"v�4c��Z]����PiN���C�Ћ��s�Z��ed�m۴��"�2i�Ý�4�VZ;���7QJ�Uo�����;-�/���y����h8�d[$�����f�lLS0�5�����n8�� 4x������ыă�w�vW���.�a\U��Ka_�>�LK�aXW�#�L9
�,��,,YY��	j���삫�h�m��oϜ�+>��	zhH�cEJ%7Z=B��D��;c�-�H-���>���mf�:1~>R�wD:׈y���Zp?��f�,��"?�n�Q�AU�JmcY9J&oɭ�-v�Y��mþ0��z/�k���t�)/�:�x�%A/���֞�C.�=��\����"d�9W��x[7Fn'���\a2\6�6|FXi�y�:/M��!n��L[�6D@C4i��ۇ�?Y��nc��Lq�H�D����*��a�� �~R�D/�x%#��j��
~Z�B6�m��/�����6��*�+�[�kG��#;�2v "��=�	�Fo�P�s��r�n�5����ԃ0��)��eHYNk���Ɍ���i/TsO�$��j��*�D���,ԣI�jޥ�Z�ȸ����5Zq�H\ơEg�{�nH����i����݄���$�2�|�.�9�*1u������a��:����ȭօ ���Vv�;?	�_�����`�Z+����q��דN��a]܎	K�]4{��jw�(W�5�� ��LOF���v�^��w�����p����@牚KA�5,�!�í�7�,:DQ�jV�g�gb�4ĭ})�+��>J�u.KGV'��^駫�h]��n~��KqrG>�� �+M ��{|~����/^�[�Z��_TnX�4�;�sT�4���ZC�P,�J��o7G�~��뭱��� �|.l��̫�л�[(������u�~ycC�D|At4z֛|����Үi�]�\m�=j���e����+�x��y�6b��?`���sA�]���j�6p�S1��w*����KA�g�	Rv}��}�$�8�^㱈
�	�낔ֵ篩U{}V~��
��`1�}hF�;���e0�0˲�h�D���5Tf��W�'H�9-�͆���X,(�8�a�5���"���d��m����O���KN��sUQ���j��5kT�6̱h#M��:�U:{E��>T�<xj	���F}�<�֗���O[*����礋�U�>w�(�x_ug4�%*I�j����O�B�md�G�r��~���LD���8P(���=p쿔\h�җ��fҫՂ�ڎ���b��N���኶��W� �� �s�P�r~0���L��_���HB� ��6 jN�2��n�!��I��i9X��>���gd�1@�2 [뽔�����YD����h4�� Kj^0O\G]�ؾ��_�@�{��� iK���_��&o�~��@�Mn@Ϋ�9�����ت�j��k�#�u�_�I��2�Jo
��|xI���y�茪,�y�0}������ r%�Yc�䆷EC�Ƶ��ո9�#�����?|��&���7����]�LZ��g�Q��Fz�Č�;q&�Źl3��!c(�/A4 �A��?�+�d��E�ނDk㮡���n��V�k=)���`���'_~�~�T}L�^��ql��a�	(d�(^��L4����:ޤ`�,�f E�Z���T���N�,��+7r�4�.z ����=A���y����X�/�ڗ5���q7�<)/�u��>�Ls��oN�]e
{��t������[�|����FN�=�
d���M�@�}���@��GH$���E�d<��&��CR��p��a+��b�r ���W����P�%M4C�eqK����I���Eo��$�ɕ4�0X�ĕcv���r/�%���f���m ���J�sz�MM��V�X��0g1o���k/���?rx7y�"8�}>l��5�T��@0�\\�t�$����g�>K�r�ib��p%r�Y}���m��=�-It�<�RR0崙"7�pɷA�-Wz]Y>������璧Y��5��n��e愽�V��@h'pҍau��T1 <7VA�:R�_��y;�P1�~.��r!�⳽�+���"Ce~���ф��� ��իcV0�����Q�Ϥu�\�I�m����2;��'�km���m�X����N}��E+�P��0��\0�y)����ٚO��akE��7�X���A�׳9��!��b�2e�JVx�=0�i֯����0{uYc'�t�Y�k�1����~3��^����݃82ؿ�ɞ/�h������a!bg�W��Z��E����ۺCw�	J�|�;\��L�E�����"[���ƶS�J�c�G���${vUʯd�J���9����u���0|&6�z���9�-�<��ƥ�����i�b8h�N-�/?���ha
Ns�֌�����YS�JC^_ߏ��j��O?/w��:[ �()��xڣ�bޮ�i����:V��xJ%�SL����sn�!��'��ç�E��'�f�1Y����>���6N��c��2 '��J}ɿ}\.C+1q�,��
N�Q I��u���Q �B�����:�Z�U�����c��u���B/��eW��q�,�IM�"����7E��lA衖�VN'%Sp�ԙӬ�pK�$���O,���2�f*i���w�q��L&��7\ �:/$��CC<%sA���N�[����|���z�[{�w�h��t5�ܙ��t���<�' n|��̖��Y�a;_�gS�5�O�%u���~�ČB��&M_����cLy���fmR��'��D9��	����E5�6��Ii��+U>
��v(��P�1{�e4��?���b���x��E9`_q�QmV�6�mv$3�ŋL��#o�r[t�BQ�Gٱ�� Q�M��)	F@��|p�d[ � ��r|N�����h�6���ssg8�e�]5���+�B5���P[_c��DK����i��2<�*:Dr!SBm��x�\h������ٺ��3�����'h*x(;P�oN�LZp8̙��+%���ϴ�uM\�)�Y�ns��;��|��ω���T`�1ZӒ�����_Q�ֺv~;��E��'��$@G������x�I6�0�+ེ���,G����kW3��0����nO���%LZ4u%�(�32A%���3퓙oױ�������D�������k�s�0[f�g!@�ixv_B�䒦�\����+��Z���r�-1��֔�����Pnړ�bI͕a&���?e�͗�Y'S\��-.ˠ"�ʌD~B�;��;�<E��Q�5���&.���`��Ə5=���mz%(�N�,�
7�M'���?}�� Ɨ�in�iA��wz� Q{�;�c�cSO��I	��;;�Ǥ�r���8���9SR?5����.-�u`��+�0s���`�W(8��s5<ˬ���zs���@�Q��5F�O�+�!��A�Q��5%��Q���6��:�%U�ή������f%x��5�X�\y2W�x��-|���R��٦�*�+��/�VΦ��L�x@��T��i�ij�l]��N �$���[�h/�z���H{Ѐ��#P�S�	Үw�.��Y�U/G6<�������_�bp��2�z��'�\��-XO�a|��$Y9M8
	��`щ���x8��A��E2���`f#
�XjTu]K�쟓�����6� �B�����Ь�{P�	E�Sf.�=���_�>��;�c���Js��-�zi��1�TM��v�G����� �7NU�ͺ��M��E&��}�7ω����9���R�7�T��fF�sJ[W���TKY�(�"��-$�P""�\���k���!~u}i��P��c�hF?uEAm�ת��#��B_��������z+ÂR�����e"��-eT�u�v�ҧ���:QJ�,��Z!w�����7�n���y4�)f0�Kf��󸱇ޔ���FQ��IdQ��V��iyJ�q��dT�����?��d�f�lA_���o��{�Ӟ���j��⒡R�	�,��:��4M���=s���N��+GjXR��'���,�S�*�]N�d�����;W����q�[3�wv�Ȭ��H�a8��E�{ԅ�/�
��4R掆ʁ��9W���bR
����8������f��u����v�jx6���2��Qk���� �ڗ�~�"������H*<�6r���É�3$�B�14�c��M+#�p�J3Nfع�W������/�Q�z��k�ҟ�8c�Zl����s� 6�@�Ӑ��oQ��3�d|S�_K�#w�
���u3$��g��f�0}u����k��ꝇ�>�
b���9�<��m(�> �#�ū�
o����PX�=�=s�O�p�[ڿz�Yi���6̎83Xh8/��|g{�n�{���9~6Ya�u҈ĦӃ�(;�|��=�8 ��.),�c�����Ȝ���>��@�MX,F�E,^ �Y9��1K�x�I�3hn����v�U�}>��5��
2{k���o����¸��v�z�̌����ՔIf� w ��xz ���������%C߁N�ߝ�1�Q�<�6��d ����� Y��xoQD%��S��)���e�lp�@�h�u������R�
J*#� �[~ʎ"��Z�"��:���́�D䫆^vxʁ�F�t��@���x�O���g͈Zѻ�+�K(��Kxѷ/أՅ�4J�e�@?.�ȇ|�G|��������L��{�\��HkU���#���a����k��7yZ�XG2܌��;X�FqO5.��ȗ~Q�)����p��~t��O>#oe��(����jw���$����O2t�T��	�֧ؼ�B�2$`�xlD���už�h�1>��2�?B�W���-C�^L�m����K	�@t���p�D��?0┡bc��{���Qú����.����#��3�H���������&H?������������[��U.aA&=6��m���	�Q.�+�F$�A�Xq/��ď����	��#�B7��)�0GRv˗u���Dr��52���1cyq���+�>��`�ccC�zul��l_xz�#8|���4R��.>��۽���j�ľ@��#�D�����gB�WFɷ�ݠERp��4t���D��8��`[�Z	��[g��.�p�����@ؖ��Kv��i���E��}����[�,���h~7/�����hM�lY^_�����~�n�ޥ�ԎZ��
����Yp�p∟�SSZ�4������A��������PO-A��i��%��n+�$��m%&��������_�� �*�����/�\3��GGsI�\�Mf2ѥ�Yc~2 s�R~�3NB��g-s�$jcE����#V�p��Ӝ��ǋq0����j
k`-�k
]8��ü;���d$�73ࡸo�Ԙ��l�6�M�	���J}#߾�%򞼄��E+�RSZ���f7��-�� (b����ћ�We��I]�Hti��^���6[�~͢�X{�K#V��촀y&P�2e,����JT^8 Q?�ˣ�a��Bb�	�[�K���W�%N�Q�ߐ��pNc���2���n�6�X��K��	�����R�BÞ��ˏ,�S�{���r8��H|U�S�q�($�@����#�L�C���9��	�]*�4j;g
(� s�����Srϰ��AZ��d��aų�ŋ��)��?~�I泠��!1�8�aN���6��i��_c�`��ꥱEE���	��i�c�H͉cFތ$ Ldf���?�*w��e�!/�MU0��{!�w�8��lf'�fw��J̑�6�]\l�:	d'S
�
)���{��83�Y){�6�@ǫY���u�6�g�:Ȓ ¶��~ד�5шʑ#���8]u���:�����g�ly��4� r� ����Xk����w_���]-E6��c����c�k�uXG��"�nn�@������*㗘%)��X�+���'{%�f@�,��7��)�e���T�y���DhL۵�ݠCҵ7�ƛ�m*�КbX��}�+� 0�9!u�{��{����7_D�n�	�c��`�uS������`��JU�҆h-�� �
K��V��4�qmV��*3�;;�%������[�{X꟡gq��f��
���\f�C���  x(Lq��z����}��o#����TI���!�>s\v�����p	�DD�Va�5 �H`�,�aSD\���\L��o�q�^{Z�ESn��K�Î>��x(W�:�W�I&�0K���,������S` ׫�q�3�5EP4���[�
JI�O����[�@.���xp>#����#y���U����%�wQ�;�oM�>�̎d�i�F@��:Yx�M�@iT��h?3��5̵��|�-�6����QHX�}���ێ�a:�O
�b2��u*�1Bo�$:1a�h�^c���3�i�� v�aNo}�/��0�q���W�	�0����i�����V��?X����W:�K"�4�>�t�
LeCd���އ��oP7+M�-�>���9�P�)<�{�+ �"�-�[�-z/�L�y�=����'���vE��S�������;�,�g���e5�׈I��s2��J��3[�(K.9
R���5�6*�p�ͦ;Q�l^�׍��h˕?���A��,��vY� _��H؞_]��'�C��(C��E��2#���[���oj��!��"��y����ي�(�y6�b�R�Z[��!E��|�n^ݶ�X���bpQ�Ё�<10;��`���֒�����5�b�z�r���)�\t�D��@t��f��b|�,�0e:]��\�	AF�o;|Ga�F�;�)T7,�ǼҀ��n0��V�:�ȄSYe5�䝕 鯐aɎ�zN$[�� ���IU�ji� ��'�)����`W�r�1�A=p�'6IW�s�O���<���%�Q|�-[%R}κ_'�"�aJ�@�R!�������_�':�n벊?���ǽP�Eh?��{��D�|Ç��Ou��B�5T���o�4�+���~)��'8l�M�*{ǉ$T�QZ��a�=LD�����.�Ո|7��Օ!�:�qA����n��W��*��C��z�[��� K�7bv}k:s:�"��ӣ�A��u���LjZ�O�±@.�CT%��.���ۈ~�!����J5��خ7�
FSJ�yR˲��pg��pBD�?��Q/��.��MǄ�4�T��L���Y��b���dt���d�C5��`@�	x�	���Mp_��.�Q���}X���\a�ը���qR �y[��Ѩ"���O[��#˴����P韢	��ߐ]�h����w��
�N5mL�eU��4���&�Z� �p���*s���`�Q���U'H��k��-��s�T���w�by�4�o�d��h�v��ŅG9�M���-��Fc�43������wMs9u�ֽ_H�bJT%���$� �m���m?siP1l���ʊ���ݐ���Xـ񭾞@�k�Jؖ��:�-���Q�zm3{/�nJ�=Z�Y+�4P��x��cK�
�爄�؟��h���,�}�`/
���#���f��L��^E�=x�9��Qg�bKc���G�c50��M�u���5��%q�8�$�a�UV����A/�V��HW"L6�fȶi��]����U�� !E�l1^#Θ��q�fvF{em��ҏ�(����!:�}�z 1d7�N;E6Ϲ�����s
���RR)�U=4>W��@=K.GG��B*�fC"⮦�4n%�/4b��G�\������].E}s�|W�PR����A��fa�#HVK��j:������9�����7ܧI�(����˪��օ �ܹQ�h��T+��j�n��n�
<?�e�Y��5���d�lS�2;�h�_�}���X �m�8�tĴ���"�jz:�	������;��ZX��fao��u������E���X�ZR������[�	��k���I�-���5V,�2 �{�ӎ�#^"a�e���f��1˕��K�)�E������A����W*��MY�!�O��1�ǽ%׶�܌}���,�k�Rg�K��s9\3ۦeOr�@|̮<�V�s�E��	�NYjе�����>C�?E3��r*^��F�+���u-T���]�����o�w����8�l���׷�4cR1���a�k|�q0�����p�!e�4!���!~Ø�]z,+�-�1b�SC=��	A�#:˖9�&f��<�?�Y�SL:�w�~��a�*�S��~~���)1�#�	`��ڽ4&Lg���ݾ($"/����	��_���������؜ٿ7�'u4P��I;�ۦ�\��+��^�7�����u�o�`���� ?8g�Y`f�{�k�Wl����a�Y^�Y�kz3F%���eЮ9^CܢN��I�4f҃��xN�T?|����lӔ�i��V��no��_���	#Iփ����x-c("�^�#��&[�MR���?�H��S��us�D��.��,]�� ��X��u�
�+gBdd}���.@D8���7�����_=�M��:~#�ذf�;��dn:o
�j[����7u7E���_���щa׶J���{=�d#�׊U�}�W�㒹�zV�a��*���v0B"!�q·�Y �	����k�{�ۻ�(�S���f|�d�bd�P�������;��.�ܐ{?���}rN#��f�,}[F/�b�Q��3�6xX7Q5K��!�+(���XFg �X���!�	�G�`�n�*:g���#�;�Ʈ=�
#���Ddl�-#0��w����@�1;n��Z�	2����;wv����n�e�0�v���Jj�l�$t3g�T̨�0�g����1�Ԍ(�~~���n#��,�	���Z���ǀ)�O��=3'O�R���a����&�����Ҟ���OQ�?���*zʹ�W�v/�+��pL���ۚ�*7Z�M�R�F
f2�RS�$��W�8��^0���,QPD���D��I�Ҫ
��շu^65�э��Þtk�5�?>�>͑I�n��Z�w	nl�]Tg�f�45jk��!݄�����M��J�Җ1�HW�E�me]T~���B��0e�-���M�;�a�Q$p�`؇.�[�yTb�ʋ�'���>���#�*Ykͷ��,I�)H-D� |K'NoU�-��ct]C�d��<���ܧ�}M~��n_��-�j|��$O��rM0c����p�N��a/�s�@�{�}7N���'�8��"ӞR�#X�K�S�"�߮Vmx�DS�'r3�~'Uͮ��Q����;�S�V�NoK|�mV�\��DL�@sz��oaF�� a��7x�.�^ӌ��Jf^$V�r0$�'YJB�2�m.��Nl�=�3DRc:I���E�e�{&�g8'a?g��ӱ=��!u����_�w����B5P���)�ӽ�,��c���k�^��s�S�IzI���+Gk��8`a���F��%>/�p,��>Q��'>�(ڬ�*�.#S��������&鐬Kࠀ�Ş/��9�Rp�(��˚k����&�/-}���A�T�0���m���^坲���'���y|fz�%Pʯ��������f0z�~�{�K�P�m�����R�%�~ÒSZrJ��vwDh�u3�e����kce��·��y��֛���8?���[7o��a
�C~�I���=,��S^D�v,�Z9�r�1DL�jDY@>�H��|�"�㰫��8t�%٭�W� 87(��ʦAw3��l�[�܊&==i�U�oć�k�I�|]
���q�����ĝ�16W�H������9�>��5L�����pEX?��U���A�(0��-�z�Ƃ�A�a��n��R�kA�'Cyq�`j�h���H��1]��L���+:�ςu��Q;A��G���
#�i�-e"��G�W���&:�[Pb}����nB���7v��&c�i5�*!7:�u4�!�Ěu,ՏI�*�s��'<�+�>8��H�uS�H,_ſ��:��kFW���<y��/�w�<_�ţ�t��-\���uG0e1�v��"l�^�Fmҋ�w��.y��{����M�6�[�}�5��m�Y��'�5]��u����|�>���#��O�D��7�32���9���H�$�wD0�Z�;�3������,Z��c����o�����*�:\�d�ɉ�p9^�?�.,f�Tl�r=\��H�����,��&��񌩛	g����@U�ΉV���,b�UVظ�0��;����&�<O�����6���J���ms�4��y�g�ҟ��2����4e&����H������S�_��(����
�Z��'��^$�>���s���:}?��^op�m�"��7�Sn��.FUD�VI%��1Bj��^���e= �鲘ȟ���>ʒ�q��>A >	����]��?��%�/� ���]W��hMk���`��QC�x�A@��WdC��g�n�Y3��\�d��k��+5��{M��M	�����J�i��8G�oIM�ke�M�Jb��#q��⶚h�O$c�� ����n	�k��|6��M��C�֬���yn��Ȭ�[7�KU.\��nm��7B�#	���3Q�!걡"F�Iɴ@�j�*'��5�u|�)�I�L k���(^�U��-�#+��W���*��ࠆ� �<��v8b�����xû�7�tc������t��|4�+�1HAC������x�r�P��w���ZW �#vD��꼪4A�%�V4�U�y�B �����r��-ޑ~=��&]���iY6j�T��&'���Hf_m��/�G���!+������g�Ig�]Q��B�q����eٻ�@3��l*��H[�$ZMoc���C��ZL�������C��x�3��r�r�)��I?�sn�x}���i�E{���&������s+�Z�)��� c��;���)��3*L�-!�m�sS*ڽ�����I��\ͬy�� T���7c�`˹X^AUb��sx`���|I)�M�"��y���ǒ�>�h�#?^͑n�h����d -�R�W���)��W9�Ea����.�Ӵ׭l����Y���/#��c�pE��L���A/��"9���`Y&]�}�	���:�)3�^��^ ݰ �v��3s�Ϯ�"�\� G�]J}K���F%U[{?�֛�KO�@�ٗ�vS��� �IZKj���n\g��g�zc�^���cS��mI!�	�؀7}�ݤ���Xh�����_]0���٨����?�,G4tE���bx0�5����S#F�|޹A5��_N�	���^�{i��xM*6��U�<��x��1�(�g-Z�A��_��`I��1/�ڗL}*ܰ�H�:��8��Auq����s��a/HD��q���zW��B`S[�Ak0��T_���t��D[ڧ~���������>)	����Lv8'�x[�C��������.~�������&���{]+&�a?nF,��6�H�Y���Sy���CXyY��#�RvU��@b'4�'h��� H��?�g����&�<�볈�!lv�l��	 ����IX�At��z�J��M��ӂ�u2�[`)����/@tK���5·]�!@�� �a#}W^9�F�_G9w�y��}����ެ�S�CQ�r������*����R-K�PA��^����Li��%���Ґ$-\��b}�(��BRD��ݗ�j{bVq��{���f)"\��iܯ�ߵZ(���) ۹2�F��Q���0�$� �sI	���]��h�F%c�C�w�񆛥�����zL���u��wWU�����7�6����,�=g�6\�v�e�+Dמ�
Nn��0lb��8fsNOc���k�X�X�J?u�R�Dt�~͈���@�f6]Ӵ�v��Լ�'w��DL�G֗2��2�W~H<���|�O��{+?���T����\�}��e�;�<�G��-{E6�{��0����7R�'��$s+�����l���b�-B�y�P�W�0)=���G�G��J��3�Ժ�ht�k!��y_V=������=;�MR����~1��_z(Γ���h��� Li�Y	x�a�[���i$��]βO�s;�\��7����DY!Z�@W��W
M�H3���9;w0�~�ܭ�M"��ڠ�x	��G-��_�,sc?���u
����ʳio����Q7�� )����E�S�K�Rnc���$�?
�����	5�˂h7�����t��9?S����}sĺ}VQ��C��Ph]����c%|NAjChB.o`�z�e�����oG*�^�}S1`����(�!�j�MP�x�kw��aWf��>�!�*%z�kS�����~��3?�4F�{H��p͊SyNb��	ݭ��gs]��BsSSz� ��X�'��܀`�[�� �(H9{k�@�{aYds4��k��K	��3n��R5�`��*:,�7����S�&���.��������9Z�f��ҬE���9΃��(pvr�V���b�9������C'�»P�2�hfTӣ*��@��W�����D����*��� J��Q�XT�Mtś�9K���K{Վ�W��+w�P�J���y[{(�^]����� ��+P8ØzkCw����%�q.��|o��`�[�􇈭V�߅ls$|N��re�;?�1��Q�L��ѯ��Jt��r��J�P�
"R)���gxj�1Q�����P�o��(s%.Y��㮙��][�(��vDǊ�p^}��a���h�X4ڥ��f�='a\7���$����͖Jh����u�J��}"��y������F�c��l�uc��i��z"W�&5��;q\R�j^�=��Iג�9����Uī��z&�2���T��~qF�w����#Q0����Bnp�HsB1z�$�0�I�z�O�G��<��У�l��֍) T����H�u�\�J����������֓Dw�5�y�r�`�P����g�#Ɩ0D�KY!�x�����3�'"."�p���7<��_kB�İ:�����܀�3^5�>,�496���_yrL����)ͼ�T��uW4�W��"5��H�xd���6��,G���yA��T�u���~�D9�}Ո���>�����[WN�!A|q�}��ɷ��s;�(<��t9��xr �"��0g�1n�:l�DM"�k�3T�����;�������;a����{f��3�������i�6Ȑ���U��z�ǃ�PG	#�tx���G%R��)@\���kƼ�h{稵�c�`7SSP��^E�9�(�HW3��[�E�r���9l��*��٬�vY�n@1�A���N�fgfTސ[��Y,��W�{��1f ��&`��c=��е؈��#߬8����O��8�?I�M}�k�����}��X��^[>�z���2�ŭ���֍F����ϓ�Q�ti�ȴ�2�kL̚�Fa��2�DqG�i���kV�?����U����l��h�Vзs�N��R�]kѬ<���M���\�֦�-3<�}~��-�$y�J''��l�����K*C9�d�f	'u��7Jff����'N��k��bW֫��$�$d� ��;<�ᖳ�v.���Pm�fv�mQ������r�aj�t�b�=y�SQ��wz��c{MtN��8	jb�'qܒDN{�J�Q�� ���������Gt���0���.M�	��|5�W�HM�\�=�.vF�JN;Ѭ���9�0 ��v}�_�~��g���d�z5����2d�x�����^Z��苰[2/�0��td����ZM2M�ޭY�ַNlL�l]α�NO6��P���̵���Jt����L:$���^u9e,�p�Z�H�l�-�
�$F?���r����i�QޗD7����S�/��g~ ��_ �����h<�)�#b͎&=��gj��:��M=����S皨Yj&�`���%8�{�+�YK�"�2��;"rq��Oq���� ��uW������+2e$1}�#�2�7���ш�h����7�U��"P�7�E<����/Z_A�L��q��CC�ov?RIӇm�"R
D��!Jq�u�I��9\�w)=����A����6vx%��I.��z&(�`�<H*��%N�(���XntW�@��N��f��� ��2Z&�]�"�c������2?��������{iȇ���#����Ξ�&U|s��&@�~c�	<��$�hs�����|��R�R�B
|Y9��p�Y���E<]y�$���>�F�����,I*��{�yt�i1�B��q�R���b��`���%���F��4mF����:���?75��y,c�ԟ�bF��͇X�1i����!!�/���ހ˅�3(:L����,�mں��E���I�?`�ߟu%�3�,�{�������m��iV�R�y�	���~X4f�n&���+��f����Y���V�GM*��h��l9�� �鷟���	S�+�d�Z�[��6���N��h��Y�f]'v68����գʳ�`�W��G�xL���;\e��BoHC:���"P������F@����<4�U�I�a(�5J����E<�s~�Q+CU�˻3��X���.1������bAgj�?��9�|�K�@
9}�'k~*회�w���S���can
 �!�s�.L�4�23Ќ����2����e�BPSh��Y_4M���Z���]s�rSڷ�sڐ�~u��O�E�ґ��3 �2��"�z��F���ERm^Q.��E�DL=fzG�6��O��͵�&]��L`�Җq"��*M+���z��v<�����̅5w����\ � N���A��l���,|������@����]�r�)��A�;�w�n3Upp��=+�d�H�LS(j'9��z�?z��V��[+\D��Ց�o�j,B�I��v�g���W)\�i�9K��Ks-����/΂����SC�Z�p�hY�o{�q���I^�a�5+�����i�(�o/�#j�]@ �Ζq��@gЯ!��`}ᎸA������b?�`�c��NF8=��p�����y(�˴������>œw�1|�f��/)�;��%J��Ⱀ\��"~ec�o�OJ��w�G���Or�h̻o��Anǣ�(���$��q$�ܔ�}��U�4�J�O�ǭ�E[��~.`
f�7�*J\�U���4�L�^�Omker��:'PSt�Wv����#P��'��	�]��	A�R>=�SM��5��`�N]!L3>����:Xa%q��_
Qk�!�{�P9������?������H6����a���4�5�Z�!*��n1}>�����ߙo��������ɰ �Tq��ZO肱����ɂ��c�N�ӱ��Z���j_����rXӤQ��dT%�j�"{;�'�#�4��b[L�/k2b~�=֨9��2�]^ZUQ��(?�vrj�/0���Y��䐝�����-���^��O�A݇ª}�P�y}ѽ~$&$�M���ꚺ� �3g�=[�&Cr��W�R�4[�����~`�-'�N�Jd�vn-HL��ou���~&�z֛��:��8��G�Er�2��K�3N�����7�rN43��A=�#"L�s��ٝld�?~��������TZ�����ш���HS����ɉʙ����+q��?�U��@q��Q�t�b�]� ���?\�휝��(�+/�q�m�}�B��_G?��+%��V"�~lK����M�U ��� Q�õ�<׵��&��T�7�[��_#�O�����t�rY"�'�ƞ�k�0b���|�e��LRDV��s��%$SE���pV|�l��X�H�b.0���2�U �:)�<=ܛѤ9�U��%�g���&g��������D�^wj�Xƨ9��d[^7��i��^?9����3,�X����`���%-տD�Y��&�^����(j�[3��԰]�/�O|��᧙ #O��>a����NO=1
!�9
r��'v��=1�m��5������X�l���:�G�F�5��t�
�눏�v�X�����	�Df�ަ�^��[2�#<.)2c�b`�_LJ�o$A�SZ�/ן�:��}�E�2��+6h64�N�e}y6��IrP����`q>h��bK���H)�?���j(���ECu��4��?��@����쀑9C��t=������/o9s@#β|�Z�-��7�����$�%r��`����U��Ѿ�[�:;�� t�W��R�cm�ް���~M�;k�$�����Y���U�����Uyxb�
���uq�_ �W�4r)$GV�'�	nFq��� QgIC�Z)y�gc-�r����/��X���ߋPݦ]s��[�2� ,ec?�!��%�kR�f!�I�:L:��	%E���Z�$���(-��P� ��x��C�(E��P�8�R� sV�C���-��(ʋ�Y��C�d�^�ٖ?��ސ���cP,�I�����%e��8��~��O�Qg��@�����6�FS!n��V�g~��@��J�!|�:c\�N�G�G�T7)P��WMh����iqw���aU�e�k`eu��đ��PK� ��U�m�I�	C.g��[�rb�~���qN������e>v���S���5�Wiiq��:3 ��4��	�<�,Nf+C^i��e�Tv�#Ԙ5:xtvh�� o �Σ�Ki������(���!W��s���N���o@����-�j����gU�'��GF�AzcO����?����i���ٓ&��1�&l�4���y��&�6�(�I�ڒ�+1�Վ���6���v�Y�S~��n�e����n�H��rzK0.ɔ�@-aQ�� y'�7���S.�|�o�8}?�߯o�[�f��$�w�n�_�'��T0��Q@�4�p��-d��qS]�V�q�0�}�!�DK0[�DS&Kk��W�@���g�|}V9o��x��:�;@p~/K���!\ڳ�����-�{�B�-��j�,s;�>^���/^�_��*�.�$+�ʳHW�Ak='���y��a�T��®<2�����]ɬ��`t�΀�'o��j)S�HWq&��)�`�{e����jP��?������Rڞd�k��M"�P{���ڥ�һn�^YE�h'��h������s9+0	����cCj��)3�;&\ww���� <��EV��v9m���ȟ} J���s�z��D�� �X H�q���V�T��6�a��� k��b�sxG�h��~s/Zr\x�l>�Է�����Y���H� n�q��J�ъ]� Q$�F~P5�ά����H�������XE�e<M@�OzϽc�&r|�qO�Ji¬�r#V�����b��G²� X�5I\���g���W˵�2�RE��H�n�����K�Ou?�`��}��)�Z�P֧o/[�]B��j҈��كs�me�d�n��Ńa�h܇C�"=�U���Kw��9,O~r�O��~���G̜�#�&�(0�VMD����jb�p� ��hMG��E�d�>%�N� D��S�͹k �QH.8�0͔�B�o��8���
��҂�%Eo��J�ςh�{�x3ͮ�?-.նkȃ=�� 	���gQ��TmH�fI�K�O��xt`�oT��;5�t.��g���$�.�Բ�	�R��9"��x�q|�;���v� �α�\J��L�0�>d�+��qi{'�*q��ի��h�o	��>���g߷~�E��w3`�\�fҍ�j���6����!�@g�I�ˌ�Sc�UIoή�!Sv	ue\��u���&ʑ�>��f"��Q�?ޑ��̧Be�s5�ɘ6����u���ԧ1y��� fOc��Q������(�®��R=���X��� YW�D�,[��L����fn���;��@@>���gp�ƶW�
��=��L\��y�l�*|��_�a����M3}�f��S�il�1�0T�͏\���_5a�o?�ܑ���w��H�߷z��,C'�#7�dNW� ��c�9P1�K%)�1.�hk4��-b"L:QF�����M��)0��<�� �r��4�I����C�q��(<�PB&��ff�o���k�6�
������j1�xJW�"�,�}��$�Ίy`!�}�/Pc���<��!�%�X[��x3fݍ(�+����������_�@�yB�D�Rl�w�1Y?���d�
,�j�uJ�����,���i���{o��4[�HvK��΍�x���4���+�?��*ѳ�ؖ5�!r�%�ЍԬjW��H,�W��I
+�Y�����*���B�7)���,��ɭߣ>w14�oQ��ۦ�v8�_���8K�\(I_.\�/�o&�M�`�y��<:�~S5J\%|��8�L@W@S	n�c�9�M�0eP��J5Ht�ރ�: ��h�~zO��򂁸�B&�>���2�T�:�S����*S��1զ�糷���z\�SP�������䔳a�?�� �vw\��W��4��$x�8h��`�f%O�$�M��D�,Y����B�3�#����n�TK�y�_ZjM�q���(���/��� ����	��Ѻ��t_-�3#�GW#��XGH��7�LoH�k�`[���;M�d�ޓ/�{���G�2:��U<�<i ˘cW���LM���0�L��(�
E���Aֶw�����!]��D�O���Ht�$����ۖ��O�Y����.N��n2��'�'D��*gW�m`Lā�(�`OR��V:��'������y�\Sg�֢�pư{L�dE =��4��(�+{�q݌�t��r�]g�7̞��~kꙈ������5ː#�CG��g卥,HI}�~o��L�c�u+q]�I��]����G0���>����kf�ǌqI�=�n���A~��ٕ��h&\�.a(i�ɛ?�f���1�%��Ø�|3��u��I�s:��"��YxY��oQǼ��낕1�W�Ӊ��S�Q�2�$��[f�
M_k�>bOM��Sя&!W�ӏ#���i�7�d��"[��F��&�MK/w=Q�m[zo�_j��O]����> �хeu�#�H�:ZÓ�)�;�Vݧ%M����Xh�yD��9D���荍�����iw&\� IWZ�yf��m�6WA��4��C9h\[F��En0���hkc�����\���ƺ���8�M�o���0�M��En[��Zq�p�1&�Y]�Ԕ�ZF�N���-���oX}ó�h� �$m��6{��҂�m�TͮI���{��z�:%U[E�|L��k�oM�!��p��@8��VsX&��,�����'��	O�ױ쎦�ED��N��Ud�ٱÇ��S��#Y�Z1���;l׼�pCCf�����kōw�2�[p�iV�#$tͣ����5�8m�~�'UA�����d#5�v�`"�8�
c�dB�8��È�#���.�u�f� �����
>/D��_���<�q����ß�ݵ}��(��1Z慉���g���
"�OvxH�����NVL=fz<n�e6e�kQŠeU"T<����91��ǿ���[��_;�ᚺ�{��(J�-��F�[]���@�U�-�_�x�,�7��r�����&~܌`����V.:� �t1
�E�%���6\f��a[Շ"���A_�D*��dz�_e%�s�:n���Ra��w��F/zⲈ����zy�wj+A��:O��$�-��iܜ(y1����������s��d��}T-����x
�]R�^x<�V"��k��9����Np>��-��)��.E����X�l�w���]�.����=�Y�~ٖ�m�A��|@�w]�ʶ@Y_�GL������w�B��2/Фu�ya��6Zu,�~%�e�	Vʻ��F,^��t
�ޑ���M�彗�oX��s�K*hU�G��(�d��E�f+T����En��Tf�gc�};�3��\�h���~mY�\�0��iC���)�`hHL�񘹎/�>.,��e��G��>q��}�ۼ����t����0K�B�m�c1"����Y��µ3�"�V'��JUs�s�n�|(x-�n��SM����>%��_���pѽ�7%�A����Y�u�9����;ﵯ/*c���9��Ey匞��%�R�m>������捃�I�T�r�ӟ3��Z;�����7�/�����}���v�׎�RԄ��2��(���}��.T�Q�Ya!������;���_Y˞��;nP�� S3����k��o,B���1
*s��ۈS�!li$�	o�� �T�:tK���h�E��9��֊��k<;#��6?�G|]E@��ˤ���`=��L���v�/m�^����/7�U���k�t��cB.��q^��fR�¤i�[9�z�"��*��v̧^�\�jО{}�gn�R��_�S[5���y���Rr��[��-rQ�/vRҤs^��WVw#K<�"�Y�)��^��Y5����/u�ݚ����G��K:P?o`�Z5V�,��ˎ ���&ɵ�dX���鬟�C�uf�a�z��2r��1�����Z��%Kca�Kh�@��%��
1X��ӏ|8�h�s�7��a$x^/b�-!�����J���3��|�5x�5Z�^ّUF��3��F�Q�d�<]ܨ@?�> ~�����t�`�P ���=U��	(C�%�-u�5�ROq�|���a���I��2!��l�=�/Ǔ�����	�ՙGie��\��b���[�}d���Gܯp����4Do��D�}��"����ZKȭv�VfHHb��#ʬ	���	1hJ1⍵�o���e����"El�䢟�\����&AU��L��]��[��e���=�+�oZ���YǪ�_iź�L4ihg�q�DD�� �C�� ���#K����A��5@@t�OUU�/�8/u�?D��u�.G�@f�i���:|���w��˨�/�K��$2$�@��lp�KUU�t�������GDA�h��rh�7
!�t�W00��K���]Ŋ�n��u���,�JF޿�Z�n�^&���BrS+���6�h��y�H��ގ�-1
Bm�Q��kU�Ex�$X�� ��T�{��~J������'"^�*)}�=M�7=�ޞ�|�aNF2!���^z=%QH(5�q� ������H\�-����H��/�v�`��x��=�����A.-�J��bei\h�>E�~C*BM���?="�ށ W����r���u�(�	m:��ʹ�^s��:����5���&7���cs>D�	�{#⻈��x���v���?�x�6���-�w�3�Z��W���	��b�� #�s�{ ��	'��H�3�L��u!l�qܒ�}O(��&V"�o!,{��b}x~R5��͹�kZ��#�%����˄���t�ibo��te������?��)1�JY�KƩ��.Uϯ�:��az�<��Oi{���H��w_w=./�� ��l�&�e_�� VR5G���9��s(Kȯ����� �e~�x�B�&�eݸ�3�_mH;]�/q�Qa�%X;��+SEc��ݬ���Dq)����h� ���cE8PE
f8��=_8����Dcz��>��]��OR@�tފ�)���sW�HH6���'��Zx�G5nk�,!lT��g��?�I�:�%*e��+.�r��!ZX),? VI���dk�D�TU^GB�mSQ��4Q��-�� {�eCT����[h�M��v�u2��Z�I3�1�U1V}���H&n���c������ݙ����^r
�}A���ݰ��p���$(�,���Ǥ���{hR����kiө�ʅ��0"?,�s�㑏$l8K3Z@L��{(38�ƥ�
"����WJ�.�1��
�Y��P1�F�:�@YQ�����s�x�WyJzl��2�xz<�P�/���,�m�&����o�?�Q�"U�&eB�E%l��\�z �i�qkeм#:E�c�Ry�)���V}9�g�Ҍ'Ax��!���$�>ݙ/�Ǹ��D+���40z�?����JU�}=�;���Di�O�&�>ͪ"4��FzJ锆#aQ&Ӷ�B����e0�O����XE���b��B� 5u�KH�i�Shf5���+��Lm;�N�	U�^�²a�q��׷x�~�xĂ�o�I�c@�4���Vv��/7�&M������Du���
�����f����s��B��<P������QF�����۪�\�� ��P�.�*���kҠ%�����]wo������x
���ݎ!��QNAe�l�Q'Z����(@�O��󠋺G�
����v��J������� 8�V�<�&DR�EA
5IE�od�Yx<}CPY��7n��OhIH�A���!��#��w3$�I )�m��G&{�Q����`%^~݃ڈ"5P�B�0~c��1"�7��d�4E#VF�[d�4wW��<��z��H���~	���sךQT�,���p;�yMf�*ωK�gC$&Ҏr+C�#���q{wE9�CZ���	�*��}�L����h����1بIs<˿��ao���Y����'Ey����<r~U��R�$C���|^?l|Y��5������h�g�j����ʬ.^s�_����*��5������
�C�5DK�ހrv�^�� �;���n/�Y��>خ��.`�6.y���C��璝�U*Hۼ0~�G�g+3#����N�P s��7�ͨ��w�@�\'<?n���ώʨ��̿Wc-<	��k��g�j��Z�H�N��yEzuO���aܽ��Q�k�ki��Â.B���rO��p�lݲ��.`�0�;@M��](��G��,T��K�a^�@O�M��1��lG���8#Р��%���]o,,L$֣	������:�.H��GÉ��ҟ?�qԤ�r#!��B�p�9���M�id�H��{0b�KT�"�r�=@�f�ZM����bl�?5V:��b�޼x��C���7��ef^������A͚��s} ��~^눈b�h��.�ʿ���#hLZm����{�ϿR� �dSw��u�3Z�|IZ%~z�~��$(S��fշ��h�3υio
M��9?�`��=C8����
�����-(\�<m�5��#����_r�}2��yxRzƦ�fm?UV,���O�u>����)>w�,�s)�ec;a�}����_�+{�����}ZA�9V���o��n�d]�A�n�+�5A�6�,���p) �S�{�V:ct��_S&`#���Pk�?��3a��W���K�Sc�!e���/�c��^@�OhJ<:y��@d�0��~�`�����S�V�=?�(�~&�֚e��Vn��mDXS���Ôד�ګ�?אC��t[�M{l���)e�8���,��Csb�l�� w0���/�u;�ʁ�/�t�d�R�@f������D���8.<�Z~;+<�;T�t����҇<��/� h;����ט�Ǉ�Y�W ��6����$j��O�/�[$�������O���8m�D���'`��j��	�߫�=i�ŧ��7���Y#����_C+�j�JV!$q��uLg�[�5KQ=p{L����RV�0�������2j��줮M�ěz�>508{�D
��U0o��'	b�Qh��oH.2i�l����e4����K�ё��b�Y�IhA#�(�`����ª�Ƹ`+��t�������iOa3���z��
�V�1�i��r&�аo���s��'^B���΀*�&��:�!.kM�� �	�4 4��V�(�u���V�l�j����<SΈ	�rq��Xmʶ�n�~M�������l8�rʹ �qs�֣J�mO�x�s�'^쒴���<��1���L
F��6q}��eԨ*x/�.F}�h�_7ښ�Μ;6�g�=g �@!5��^\$\|�%��W����|z��0*��P=nJ���k�1k��$$�!{��^)z��7]���1�՜��}�������+���c��R��yF c7ba��Jִ��� �t�P&� ���\���&I��ғ�2�l
퉑��j1a�=���1W��,�?�����(C�C��n@�FA�9��Ԥ��5�I�bN��k�?P�E��$�����	iJ��c��Ʈ�5J��uQ��ӂ�'9I�̪"��X����p����lx�����Bu�~���LTJ�PLa����s��	:�s�$L���������)g9
��Ճ�� Pr�C�7�:�W���w��O������8� '����tP�����o�=Ѹ8Dbq��z���C[Cی�c�X~:4"Q
?V���i��(�����8�V!��k��5�Q���[vE�U6�\�|H�������5-��ƫ�?�(�&aX^��3m���I�:�&ю��V�7Lj��x\^�Yl��!۾`�O���0}J4�z:�[d�|����蹿�$�ݰ4g�W�T7υ.'.�k�����)��� p�9�OM7�Yj��\���7��\:��b�2�U���ӿb���hѴ�������ܒl�\�[�XL�@��MŢR���h{�C�D�׉�5#e�$t /�4Mn�?���~^�~՘3QS�[�g��_Ӧ"�J�=�b)e"���$Sn����������e��Ё�hV�2�C(_���Wt�p�׹��r�`PS���@��� ;l��0
��Ft��sU� /[�U2���H�1������ܝ�f��3������퓽�=hw\{�A�Ԩ	)A|}��.Ȋn�d@�O*��Ѩ�͡z󱏣��6Y�U�>�cΕ�q�����s�п�jhy?���F	2�$[͸/��5I�L�fm%Sx�)�Đ�HmÃ�����t����M�TTؒw�o��"���ܛS�W_$ؾ��ɖ/J4n���g��:��ow@٬��tS����i����<��C=��nf�a��|%,��Mn�f����,����5��Kgaj&A��l���%�T�-?斗5�*��|35 ���A{GjdӵU ghO��8���"�D�2N�n��砜�s�~��q�bO�oU�a`�r%�eG���5G�Yw��ޏ%큽H�x��̝�B{>�����i4��ZI��V���O��ѭv���{0��������VNG���y{�(�/=��Gav�N�vc���i�><�P(.X�2e-�Q��%���b���ce�=ð"QT��{�`��r�L���fu>�m�W���̲���؏��R�0@$"�����E��5��m�@��9�D��ϸFF\>k3����GS����P�L��	��9ÒX�(E�r�ֽ��3��҃��,�Z��h)]�T�+�w�C2�O$�-�g���-a�ˉ��� H;���&�"س�*�7�ҷ��M��CiyX�J�$��7>�����2ω�o�f�CD]6�OX�9�޼	�3œ��4\�$%�v���-���}�X��Q&��U�����>+p'�fy�S!�5���]�,�\��xnYdG)�pqvz~Pv�%ĭ,~�-�w+��~�%ի�� kR��Yv���A����\��g9���;&�ZE�3����Ĝp�k�e|���$;����K��IkV��:�Sy⛜��)�~����q[ڑ��8�����&���|,�n��>�X��SGwg�Fr����I�X�~O
�O�8yK�l�zoIxHK�_���ѐ�k�YQ@�åɻ�ć�a��R��|��Yy�E�3���~-�)(�����".�w�b5��h�0�}�@Q�Q��Q��1���k���Z����Ҵ��U��>��\�4�Jxjx��Ē�������T[I�R��V��6E�8���(�r�B�Jr���-*�D��7U��1���O����~������G:Ԓ;j���W�l۹Eu�� ҙ�K�<�^J�_�P� �J�]v���V��d�B���>;cv��H�j���UN�!����29�G�(5�dvx|��>=����)�k���y)�Ɯ>\ %�p2�oq���[*�{J4@S����-$}Jo��Л{������3dֽd��ꩶh����aE�\J��M�T+��!��(�F�N�]H��;W��{�a��~���Q7�?�����aɺ��հF��\
���f�<����t.~qvl7��6�ڞ8�R;�+'��5�gR���C�"*�I玾�S��v��׳= �Ef!dC���<�ʞl�=EϞܰZmԯvkb�t��m[�wqu�;긮�̌�0�iE��D�M?+:�M4�kV�Ebs�	W�J��
K�br���3Zr�,�)Z�3�Rb�e����K��M�I��BɬC�'�CH���>F3��&�4��qУ���a��x���_(�@��7�k��C�6��z��ٶ��^���<G�Sz�:?��p�� �4��UZ8�f���q���&d��^�F���>�˷I���>(�o�z����i�����ݼG���)�P�<�kP˹���~37,ج?N�)�s�<�f� �
��a��fH�mW�";�}�(O�����VBH78� ֦kQ��nۤ��o��F���e�< �:AsB�C��Ř�{��Ά�_u,���_����_q���|{�|e&�k���n5FL����Muw��M�oZY>4٤4M9|�V2)�dZ�h�bٶ/� -�?-�T�V?$/-TP��i�F��c��3[>x�ͱi2�F�}פ�6��L��!�D����~/�w&!(��+�����]�5q�M"�A�3�Os���k+��-�^A3ہRh��R�6<�=�,j�H��l<���Q���SĿbY�UG�q�IpF�d|yD� ]Ac��],�*ق�$z56�lQ"�+p�#�ԍC�y�^BL�*�  ߍ"��]�B�hX�j*"6?���!�
vew�nrO�:��)���,v[6�cM��r�a�]�C��<p�q̠��g�-��Od�����b��k��'�-�����F�$����'I��Y0�w�iY�#����r\U�8�;�Fs
�4S�׳�O��@��U��\�&��ZOK���|N�3�X���Z�2�F'����D&���j����@�{�����l��O�܈���~X���_�� ?uR\�]D%��1/�OϛB9zATq�����ܠ�jNl?�;�ʚxJt��~KU�oi���wY��H P�7P߫��z ���%����'!YZ=y�����.�D5�?cy0����'u��կ�J}W���i�E�
ٕ��^�L~Q�8ɴ�o�Ӄ)B���P��aI1�V�$��U Z�
ZCv�߷�Og�)�?�i�>���������Ь�m�,nz�nVd3�%�^��o�`ۗ(P���E�����:�8	
�Y���٠�s�yDG�_���{�' �,&�+�n$�%z���6ן�꽊/�o�jM�E�-P�f}N��\�.����UW�Q5������ @Ú��CG5�E�5Y�RR���Z���;��夅�����I �I�gıN�j�s�^ޱ�;��o%`G�xs�?7�V30H�M
�z��05)���f2�^�c)N��=�ɡmZ���N/ci��_�^����-����N�g�H�$h�U���_��3#��f�^y�w�l󽯲ꗷI��]�J�L�~*������#�h�!ϓ�Q:��[�.S�o�}g��58��\���9�sRt|s��	G�������1�k#a��P�ٹq�<���"�������%$0����C{$jyk���!����� ��z�i��M�����h�{�#A���i	�~�hZ�	��w�Q����rC�4���b�:�m	���F�N�~�j��i!@mD��y����g����f
��)�=5AU�O(�ʕ��iך���]��������BN�T��`��hJ��{8��"��.��_��R�u��i��B�\�h~�5��]�ϰK��P�C������H��Fd�?(d "���F���t'`����~����Fh�V+��8K�㫙fb��8��潓���K�)�w���p����h"�m�T��v%��4�S�Ӎa8�A�/R���D���$6�f/'6�P�)q�I`�����Zƺ:?���+�-e_M6�
�(�c�2�g��3l�^VZ	�*n��Z�?��sS�p��_#	��k8�O�҉�E�&��Jd� �}a5_�s�d��+�	���/�	m�%X���ӘP4#���yC|s��YRH�f�DW ��HLVN�����qmzC��!̥�Σc�,�ō����0���1��4�f"��N%��"�ӼC���(k�����^��5�5�e�Z�C�?�	O%'6�H�>ĭ����;�N�m����U�͛6)�~h�
3^��{IY��1��牺͓z$QVO�^9�\��@���&K��e�a�m�h��J ']vn�s,���'�N8�3 m���l�Ng�Bȫ��C��ג`�!I H�Zg�+3],�A��xC�3�#��)N���B{�#�Pɿ����3����ϲ��'���1 |��XO�?B��1*��	�N��Q$Uo�O)5ﹰ�%&@�=|�V���q5+��OI%���W�*aYK=$y��?P�&����A�k�{��ŉQ�h��tJ9o��vP��!���X�`p��.�pB�HĞh�=07��4+<7NĠ�鶻v@���`��������,��}����[t*M�d�OŌ�,�|r�G�v=�M�y}�,y1��oGeh.��E�����AA��0O�����n��)_����o�y&%��`h���~���+�
;�r*��Ѓ��
�����K/2ɳ�i7�2η����o���v�q�i;:G	WZ+��x�.h�$�dCZ�x���O2�$�o��1Af5��G�Y�ec���d��O^2S�[x[��v��
������4�����'�V�7	9ѫ2�ժ��p'��ꫡ�����`&j7{:�nRƗY0Ʉ[���m��1��]x�J��_9���V���S]t5�O�"=r(�!�C����^"#�u�� <�$�X��M����@����@x�8ҨHF�D��ZUl31� �W�~��*!�H��bDSM��1@��>C_�!�(�Jf� ����M�]�6N�z^�$���:�.+�^u�	Aj-9gW��"�J+Z��T������q�L*$VK������>L1�ط�J��e���� �6{��P[��EU��ֵ�:zz}vL����P�nY�k��,�.�+�7��}��[:�)�����$�q%?zs���B��vK �J�g.��]�y��b��ѳ�@���JJ�F*���H"���*t�a�D3oA.%KR�;��~��3��a1*�v�V�&Ejs^R�bA6�y����U��{�έ�$ �m^Kh�#�)
���'�Eeҳ^�A�H�!�$KP����_<�Ag�%V����j���K�}ĵ�g!K�M�7�f��G���Y�g�-7D�������|E}��ɶ�Ӹ��sis��$	�MB�US�pߟr��x�8o���E��Ү!���̣�~N���x�/΁�B�.�����J!$�%�};&�D���o[A)�>'҂Q�f6�8wh��G�}�e�g��F�I%����i�wO�ݴ"���آS|��ڬ[�[ɘ��tB|����)ߘLU���S�g���d�j.W8�˥T�z%w�?3Y��s�N�\�B�x���B�� ^����dN�D�M�+ⷎ��	]�����?Ȑ�#���`~�Z�n��մ�{WIp�[��V҄�g`�t�Y�m:��b�J�L���>l}�D�m��p���S&b���.�[�oTl|�iVFe�K�w�Q��Y;�4�!���ͤ%��+�&)��x�5j��jL��a��$��Q��|Ѫ����*;�U���s�Qb�_O{�7W���f�f��hQ���`cd���D���]��5�j|Q �\�(t�z�'����.w���a5)�)��C%@v����<'�ȭ0�����G}�Yg��{�acc��D���1�*���3_g~[۽m%]@=F�T������Q>)W(�|0U2ÔQpt�c��jOl�ܴ���h�\&��8W�2��y}t��M{�����\X9\��ha�s���Sf��y+d}Gh,�޿)ĉ:�C�?{|9T�s����!d'?3CQN�YtH��Z�O�<�UP�N��q
B	p�p�7\��4¶&�q�~،�z�5�V�ܻASo��vCV���ծ,�mo����lS���zF��jG�#�Y@YhS7��T�'�V�����[��e=S���%[�hL%ύ�L᯶%��A�OVb�"�c�bjj�}�����	"���@v{��$�{58��m� ���� ����4����!ӧ|�(cwE�I�`�=����|~���Pw]������\]N�
Cg���&��3��dْ��/��g�I���:�rGC��� ���P�5��t#1�G���_6/�[F�J��c���G#���`nڸOu��;b��.O�I"�՛���בB	4$���{O*���glh�z�
#y�gZt�ţ8�/o�\.������9�'^�Cxv�*i`/��6�^��й�Կ����`m/]Y��΂Dn�vq�Q�*[��,Ǳ`�o_��-�5N��)`ge1�W؊� ���͏(���7�A�����BZP�ު:a�z(<!3'��,���%E#:]ʳ@5ن�s���:���3vH�/iK~j��ھc���6����I�	H�@!i.N�� <���J���v5~^��r��Z�Fr��Q�X~�4qP�	�N�7�/&�k��Z	�ȩ�F�ao-��ϝ]���1K~�W�t NI�τ�5"���P�}�#b9c\����
�S�B=^�Gqz��M"s�K�X�p�Y:�<IQ���.b�΋�԰��K�B3tG�PT�'�aȀ���?���2Zpz 6ׁ/�֖��M?u�%�;�q3tt{�����G<�t����c �IÐ ��e�g��/�ukW�>8 kӋ}KtD��0���!p�2����f��д-N�\�����`c��4	����1�9�H��>�ʡ,���i�+���DI�P8���`�5��3񇟄��`U&
�j��y��+`꣚{�2O�O��m��e!�7�t� ;Z@��͟?����	#�e�gV�G�I�6��=��Cr�\��fG�s{7o���>��Z��F���0)7ǥn#<B�`ܤ���G�b��E�K}�l�8�Z����3o~�/z�	LΙb�QP��r�`�4�E����=�K�ם�_e��j��w[+�l��J����J�RON��E�������%�-�i��o�z�I���������Z�z�="��A���u���Bv�A���)xG�A�0����@��17�tntW��/T<����˰����0Δ�G�O��TT���^�9w���J(2h@'�ζ$��R�:^qs<���rQ_gJw*��NE���)�h��b�dU���ﰤ�o����� �/�|�3����[��@����ՠ���ni�B���B���\O����2���w�B�ư��]D�j�� ��\vh�X$ء��þ��z�.�Ǹ
�-�:�U�ΦE==RV�3�����Z#����wa`{��q�&��E���O���{h��5��_N��%�X=���j�qX�Ӧ|�����L�~�P�Dh����8�x�-6>�Hw-�E[����afe���	
6Y�_c>��~.K�~"[45:�XY�R�5��'u�]D:94vR���{��e�״�#RB	X�ۢ�S�$C-�wVj"����ӆ���M1|����:��+?5y9�����s�l��g'�����E��o��oW�/#��r�Xqٲ+?K`�.�T|��q��	�$�ښ���,@Y~����/z�����4凩*e	Q;3p�Q_�+��L[��8�~��P�W��h��2�⚘�f^0\dY'kq��%U����m�fG�'4����_��K��/�|�cwb<hsؾ^��j�:���d3�rGe׀�*��z68�M�'&�oe� ��l��������ȹ�]�E$��YS��`�t 7�̄C���n1+�L;��!.���PuHޠ̄n�5�}LQ���~��[j$�};�wA����=�_^�����ر����9����<�/m
�^\�YA�-܈#R����ܫo>�]U��K�c���9��h`s�H
��X/i����Q�6�G��c�Y^+U�+Ql���0�2�*�� i���s���L��G��#8�Y#S��o}Db�1R����+�Ֆ���C��4������La�[�6{�)>�tn�O�S�����t�_"�����˗B'�\�������������WY2H&԰�]�p��=/�rJ�D�� ��EQk��
jE� �p`�J_�}_h�UW���wS��N���ʎ��ݺPn�L��$���˪��<p�}�#R��\u�ܒ\��v	��s�?�޷��@����5��}�mSW��b~Q�t9;ń�+�s׌�Y�R�?54���o~��M{/�+F'�F���<=�$�Z(����-�x�Vm�c�^�L�m�)Ⱥ�D�����p�XN�F!ݻ���T� z�L��Ù�O @-Wg�R��GǦ�$~
<B5����HvFC�� ���\,��pv�=�\��z�0u�@0B+�[;����z�:��oh�� ����#��I���ߧ�CbMPW(MB��[�M����_B~ŭ_D@�uˬ�i�f�/obdl2=�{fQ3���$E�o�F�-�v\p �����R/W�Sit�2���QD�����?G��B�^�b�d��*3�ų&�ڵz<aC��S�F�Oi%�O?y���&��6�2�5����`^_�s�\��b��ϻl�S҂
���m5Ӈ�����ᇡR��'i��Ц1�s{���~1��s�G^,Z�����[����Ʒ�W�	�29Z�3;�3�9&�~-#KO.�Ղ�&�X���I�:�J~�f��$y����ه��U��������I[YrǺ��.8���.R����ԗD����f��20���\��e�j���.%O<S�έG^��&3cY�k���U�� p�sԲe�E����25����(�7D�O�1�Jc�m'�]�X���JqŰ�?�����4��fh��~���GR�dd����L��N	ܹ������=�׼~�a��V�-�5�#ӸNi`�?wѧ?��./s����@޹ؽ����g~��o.���1Ö��>�
�_��.�.D���)�2s}��T�;�@c*���q��6F��ܬ�D���y$��a!��,���|��VP�����;��v�p4��w&�-�ehM�b=$f#� ��5��d����L�.[l�!U�S�s�|���j��C��ǆ��;� 1��u&LO�TWb�Y�K%��b�D�h*躙��~��^���Jw:I�_T%�ٔ�����G9d���j�����>�d0�y�G Wj��������Re�&��\��4O���	}=_�&��?+�@��2�����I�|V�����/��}��m�v�C��a�j@է ��Q�A���>�VC��ڇ'�@�p����p��C�#T��MF,[�:K@�����XxTM��RR�z>n�V���WK��6���^4Ԟ�okX[�1�:oF})�x� 0���or���aaU��x1/�I�LL�-�[.3Nl_���z���k����8�E8'g��������2��m̶QRۧ��u�����/7�=gGF�Y�P��7�T���ǥ������/E�vo�A{��w5`�/[�*�`4>�^_�3�H~�E�A�"�����~���s�q�,/�����$hhig��?�#���˂^���Bz+-��;p�?� ʥ��lU�\jW�w����I]|�b��T��s<0�gHՕkXR�x*���}�]���̼mgA6%g�)5C�!�ہ%�x��|4��������D�3��Cx�*b����-�F\h�ne��F��2\%j>���g�q��8�A�W�(���>���i_pH����t�-u
�Az>`�`c�{8��4����h~)�32/Q�E��u��G����ybm<�Z/=x^S��F`�x�$}��������J�+�C��I4'<�ۻ�� �&P ~����;����@�4��Y��.H&r�!��F0X�y�r����p>i�T�q�j�d��g?��Ю�&Z�N���5gZ��U,&2���f��@�sS��"��_ư�V��@]E=qg�$������%r�,s�^?���$�V@�KZ���Y!X�������u��d뼦����訡 ��s�w��=�n��//���p`�Y���9�_����� W_ֈ�]�2�!��M*� ����KE�P��TDB1���u{�:�0����p/���<����Y�R�YՅ�	k6z���"BQw�>̆�3~L�(������&۴$^t	o�m�V²y��k�*}ȹ�ɃM�A��ڍH���g�,_�r�{����VG�Ae]>%�]��6�l�e�+So3��#E_�X>{���H�L+�(Zi�A�0,�p���b�rn�	�[�˹?��D@@�C������+ǥ��j�Ǟ��4��Ǎ�a:ؾ�J�I$�5&��"y@�bG�݅�Xy+N�(�!�g�ۯLܘ,i� t�������	t�Z�l�}���s]������G����8`~'���R b�lʑ� ��Ja���s����K_�&1z�_)���"�=���Ѳ��_$�Mz�S.�$'�6�������C��7�!T(�T�y��T%��rc�+����Ӛ��M�?���f�cE�D����d	�����8���'K�0�Z�$��i��圦m_VK&�-1q�~�9�#Z�&������K9X>Y��Ǥ!;����|�ǰW���EH�H������^G[��K�N�vΗ�]��>5kh:20���Nr��֭98��ta��	Y5-Z������u�&A�}[*��Ϙ*���5vZ�#;h�#�����x���S��$�<G�!��/Ţ�ܯ3Ъ3��yw�Ub����c�c-���v�J���h�K o�X�󍩢�6�̻��_.�T8��$��&o�;'������.O�������%ϕQvgOK���M�S�{�t� ��'����ޫ9V8� ձ�ڣ`��Od�o�
;�X��g�	�
m����#����:�{�P�󗝍���t�����y*��О2�
sQ0�Z��QGxu/q�4'W�7�_�q�u_bwo_q��.�ϐ#�,$zf�J�hБ��!�2.N���'�
�.���YIHZ�|ZS,?U%2��6l8�4��i��������L��Î���
� B��:�_e��&�c�CI4L��q<�}�hU۽r�L����R��vd5G��аg�\��)U�0d��^�:�a����pÀ�����t�Z��ݬܙo��
�p�d��	ɯ�@XB��C6 K �@�uʛ-���?Q2�u���@�.W���˫�����~��(�6fH	-I�Q#
n���a:�
J�6��@_F��p=gNp��}��H�v��h,�V*����T6���2gv�r�IC�ʜ7��R�v�ݽy�����*�o! ~.I�����3�<Q�ۂ���g�Z/S�9��D��z�bl#���Цtq����s���'��0�3 M<qT8�7���b�`��@;�ex���-v�@Le~�4�mU8���<'�f��kL��R�6�rPt�|F�P>�\a�S�������1=�i�Z�2���C�YL�?�ײ��1�Ƥ��q�2?{S��s�k(���+\�4�I{�-�z��i��9]���9D�=�.ϕ���0��;2����� <�b��QU�l���O��Nu��������4�Q������(
T�y��� F��}�.13�z"ED�GS�h�ǘ��f����-G�T�������X��y��\�kn�t|ek��/�k߯:*����:��,�,��S)��e�Ndɞ]pEn�}�-�#��A�=?師=f��Q���e�Ր�ۊ����������+���^K �O�BI"ߩ9^���2��X��a��⦒����J%C):��abG��l$���G���P�v�X˵��G�_(�@�/J�.�K�����{�I�8���c:�c�2$&����\�WZ].M]jL	�|d]��Nc!؄?r �2��2������N��mExgO�������ۧ��e(M��py���F��]5M���4X\{�� M����t�wF�x�m'!P�F����#��O���E����0�<�<�W���5�l��M��JϘ�.�3�g���{p���)�|Q��i T�<ot~v,�c�Vײr$c��A�����+y���ge�<x?��*�r+y�Tҹ�p�]%���@�i��h�a�5������X������A��|�)�����=w�∗Y��K2]Z`Lh���~;u���_��}�M�w�<�1�tSAKl�N �Dq
E�]�|����0~��t�ᒶ��Z��q�9�^b[�w�/��з���F� ��Gd�n�d<�R�5q���j5d-MFU�锌�M}����֍�Y��p��:^A{3�\`۪���֞c��Ȕ��|��g�,�]�p�K�����F��\�}�y�t���oI�	%Y�y�ŕ���Ѯ�xO������\�'��F�x�1���N��=�wj	���0����;'��w�H|����7�����o�%���� �֎U�5�E�vkʹ����v'A���6ʏTe�T!0%,n�2�Ѱ!���Q�(����ɀUaU����d9�Bh\��|���\|���LK��aՈӝ�gs1�bb�a��`_��z��i`�}�����r�>��Y�K`hk-r��Ԟ��<~���2걘S���ܲ����u�����jg�dT/g�v�wE����J��H���St����K�[��� ~(����A�=����[H'��"�{n��	�q|Gh%��� �xZS8�ү���G��G#����r���LM����Ƈ��:iY`��/Ql�2oxk9#a�Z�.�bJ�3H�@�����w٬��E.��}6N�Ȅ�ϒ�B,�F�e�׾�=�@�V|��.����ǥ�,���6��H�EH�rɛE��7ha��/ ̯�k�U��������ٌ�6H����?�� g�������$��|��r�6U�!M�L������@�n|���P�y���:��$Lw��~?�wB3VD$�8��ߒ�EZN,,��X���?�Z�w�I��Ԋu������K�*s^wL��m5[�b�L	O����fg�B�z��ɇ��q���@08R�]�g�*b����f�j:,V�8_[SN�o���1{���A�%¨��Ռ�,J��Ap��X�R��P#B3���6�y��gi�s��ϓ�D���ƭb���6椉on��:2�'c�b�.����r�fYV>Ȼۂw%�vm?�J"\R#�����_xNQh����;��A��Qy,&����9xp�&���z��3��-�Pt�cc���Hh}�(lW�G�;�|�lK%��Ը{d)<<�I��#pR��[S|��Sk����x�./$&ݱ��'R %���FR��4/(�:�)i�j��<��8�q:��U��	��4���
��F����?C��U��sr=v�K�t�
ߪ/�����$���5;*ṛ�Gs4��~�L��2n�֑����Qʪ�OBQ��5�2-o1ξ$�l!�ܴ´�v ��6�Zϑ����b)�%)u�\w�iX�Y����
�����7.'�}<��l�`�t^�e�,dN;妷=�X�!1Q�� �(�a*�9tj{&d���+ŐgRDw�	`�Z.�*��Z|�I�ٿ�̦���sѯKH`���b�ߊ��X��k���S�[EH�i"��H���iU��k>;f�=pIz�����̇^Qj��=!E����������B��4Ȭ1qP{~��W"�qZ^�S��Y�z$w<���H7�O!��sƀ����������"3��IA|��A�|�]5�R'�쑯yI#T�`D���d�o�e�Q��,�aJ��`fa����h_�;?k��y�Et�gq�C�|�2f��&gZ�v�F�&��b��jQY��w�XĹ�@'�����aE�{Z���9��?�|yȳ� O��[�}�5��%y�J� �v�5o��1�-jCyѪ���+�����_5��f
��i��ß���=��=m	VnLz��uy�ӽF�	v
������3�0��>��V��������c%����-9��=�M���*J[�c5��l�'.f��)Pa�B)-l���9N>���a}���T�u��M�$U&��"����ߗM��	�:���eA���a�T��kX��O�UBc,+$רu�!ԧ�ىgL@��ĳh�Ჹ�����,�뮘3����W�X�<���7ԁ����\��E2���L�E_PA��xW�7���R�sߨ��t����/�4��Yg?w��2������M����Ic ��R��.�PR����O��M�-�D^�k�<��׉�����k�3��w84�j��7���/FVe(�ߘ�sMA���N`�,Д_�7 5,��[�	�F|�R���s�8�Ok�K�5������9s 1�Q���::*7�5r�2k-���]=��_�\cuoO�;O.��y6a��au0����ϡߵ�a[.;7	,�AC>�O�d##h~,�+2�`���j���z˄����MT2
����y0{�]h;����
��X/��{
����7���$��!�+�g��]7����ÊھOA!=�R.�}2����
�Fr�n¯t�_uD�>�Z>�u��P��o9��C�.�N��;�����օ�`Q���Z+�yY���B�";���Ҙ��ZC��%ʃe�]�����u��NQK�Q�N��<?,��Ϧ��k][j�p�ϝ������'���� wȒ�X��iB^��|m�/�B�w��U
�\ƶ�l�\�'�k�P��|{;q+�Ę��
����N�nVaA��.�J�ٱ�����u7�d���/}��̿�b�s��� ���bB�@�Z�����q�����4ɏ-jU�}�ޕm4ukĽ)a���;��cp̡]�Ԉ��(O@(��y�B��4�d">(kQ��4�Pa.����!�{L%|��j[�Pj�Ao��PF�&c�3���-?x=+ЇI�5!+��:@7lXCN);���zA��s&��wT�9���{.%e�S�&��ꨱa�{uB�R���.�$���fDD�E���ƪS�4_��Ej~̣�B�3Z�D$���$����3�o/�#ڶ�ቅ�ccgHˌ��\��9����ީ�����/n7���M�:�¾�oW�=��ܧ�6g�36��A��GZ�,�>t��'猙*w��Ӓ04�!��[��� �p�(1�%��_
��x����3��԰���R-�~�����5�dK����+�n'ˈ��b�quAVk�
�k�n���e��єZE�`�*�Z?��z��Y>����N���L��im.n����������F�J,�h��a%����};Z�����o���ռ`�$��R���!���`t��ʏ�-��Ȩg�:y�,x�S�M5h�3��x��Ch�@��4�6%X��nѣlƮ*P�DLj���?M�wp�t��`o�X5��s��> $o�=d��W|���,�dk�)���9�����ʑ�/m�@��Zr��s�AT����)0�����Q%{:���:�W~>������I�9�揗ѳ���t=�n�3`���������נCH�.��|w��A��L�C8�[9k/��ݮ��ܺn�1M[�YA�,F}� �p��`6v�~�#��{��Y4G��[���l�8������$�&��q�ן~g�HJ��`)\a�gk��'[��6m�4I}T�E�<G�,VƗ���o\�b�E�5!m��}U�.H��K�M�����S�hVKS����;z�2煍� �к����6AE}������6l .�/�MK2�(��8��+�Ff��?�"�9M�O��$�T���!�7�]����&o
�o�Ѣ�NJ��.���ЂAsQ�S���s�DYc,e��������]G�K?����Q�n?}q��c�C�^�E@,(�8���Hʈ�m$fP�_���6�B=��(�R����i>���;Ɵ��ѫǀ�J1����L�Y� dkK�������}Mww�(������³���=6�}Z�����7$Ec�i�+ZQo]�xo���K<8�ʺtP��sEɘ��o��í7{�gO��f��U�'p�΀�&���Ty,i���Y�X�����
{Q�>���}H�L�ᕏRܝ\�
0����]�I�I�p�Y�e�W��(`Ǳ}�h:1�郘��W*C�1�[T�hhMe�a�3�۽B�8�7�}
r,~y]`�[���W��I��@�憚+�ŵ����
��T� Z�=�%ʌ���aܦ�����
+�w��3��P�^l�,���r��g� $X��,g#+k�Q�̢Z��U{�]��$ܐ���A#����։��R�Q�?��W���NP�/���-�I�l��%�nD�o6\�ù��_@�Oƭ���D�jc;Ϙ{�� $d����v%M�nƕҽ�'o��jWA�`2�􆃜�
Ŷ�Bf�<���9d�̀�!(�e�gnx2�E����,���o��٪]���^�Į'���y�CrmǱ��:R�n���q�a¶<�[l��f�H�M,	��yp<TGD��[2g�0�(Cf�d')�A�� ����u�ޫ�m�F��)�ܗ��anB#0���U5���3�`eI<��	��z��cXfOy6��9\��p-�@�=�X���';��M�������dJ���pK�F�����5�g��/�{�[l�$�*n�a��רl������K}!X�<[��϶l��	�Ѵr����N�D(�ޘ _^V�*�B�,�V�+U�,_����w�I���|�,1�:�����h��g���eA�Ϊ���� ���+lY��D���^&���G�4�ɱ/7}>kɷ�@mG%��/�n3T�0�2�
�{E��n�ɽv�e1dL�x���3E�7��6>}B��}�f��}�����/d�w��I��%Z�ԣ)w܁1�Ŗo�W�~`�GӪ�zC�dp�
�$m�T���a�-�Ƞ����ƫHXT�� ��� 5��Ղ���0�fkI��xk�,�*�:���� Sr� ilOۿ���Xf�5���b���
�7�@�]<�	�CA3��E}���	#�Z��e��������u,����12��6�0u��h���us�3b֚$>�����Q!Z8��HΕ���Ǔ;�
Nd�K�Vg��?�/�ߊ��Ko�:[0s��ܦF�C�����m���5�oI4�,eXh*<h$����-Z���QW�/R>sF���6�cpJ\�^�e*)��Z9'ř�`:}9G餾a��&�h�t��0���_[)��Ya��>�؆�lΘ�P������
��ª���>�a[[�TUq�˥Q�M�#:?߯I�J��]b"2)��j�f�~�2F�^nz���Ǘ=#l���b��壯i�,\�1�� 9ԇB$ ' و�����[�r�����E�
��������m������ޑ���Z�_b!B*��ze���ؽg�NL�F��'z���H��<�g���rG��(�	��#C�%�"�IĊv�����<x�Ϻ�䞲a;�>��-z�P/)B�M�$YQ5�^��nF^l�m����(�u�T�K/��Fo�韉Ju�^|� ��M=�+����A�欻+~��6;v����>�}N����i�\��1[�@w?�m���	�QH��wbk�ڡ��i���0\�I<�ǜ�*�`��L`6�x�SB�!�DB��6å�Mu�E�������	�x��2��qH�H��I�Be��<�UR8�����+�8�G0]VՒW6�K�i�Ic⃞�P���U�e��dD��lʧ�������9g�ۇ�p ��D�
9^j�����nMﲴ��T`���&���r�<2��JW�'��$��\]i��kޕUe�	�OA�"k�'�)���yն=��̅�R(O���	#�R!v8�L�!b�>�M�δ[<�P���!������������b��Q����?�h�q�B�� J���}�
��ș��O%��6:_��W�ͅ~���xG4�s����V���H�(�+/ >j䜔�L�ֻ�*ii����H�Ud���ȢBZ���Z��:S[?�v+��A@Ͼ&�"m��a,���DW��F:=/�	�Բ��0h��BT�&��ROrnZ���U 3��"@���y��Ý��
]���l�"�?��.I�N�*�L������K���ͨ�TG��.\�%mRgL�i8r�"k���_����$��
��>�У������}\��V;�(��S��拃��}�e�Ө鵮K�?$�fЈ �2kX�����y��m"u����怒��s)$v��Y/'���tm��Q�����oYە�����u�+J,z!z��h���h��d��!M�E����4���� I��?��Q�ji��!	���|-����a'i����%�*�eu��$�k(C�B���c3y,��@�}稯2�0zC �EЬݠ�#QiJ�E�usҐE����]r�0p�M\0�^J��r��c�KG�����E����cI�Dɣ�߄�1l+�]Xy7q�9IhE"�{%n��A$;����Ć�fi?M����?B���D�!����̥Z�K�焤@܅�|_�[{�H�>H��e/�`��g�6�i�����r�b�:-��ނ7B�J�V�J���JlX��*J=�Ŭ~�>u����zOT �>;N�禼�'��������vi~�|d�?��1�K��ԕ���k��J���3���}T�f��=L��d5/Ύ����{���ө�qE�{k�8��M��9N�F��wC?j�e���_�l���L�2:vĐ: � ���6�N	�ul�Qo�t�K#�1oo�ə��Uh�v��/v$��d]S��h��o�^w�������t)Q�Ӭ���Q����	��p�T��;G��pѨ�j<qꭚ�Mf[8x�b�ҁ�y�ޘ�mJ���OEh!�pN}���zp���2>��j�!!�):*���]CͩNG�������y/+>E�B��1Y�.���i=��;^���L#c+�TN�|�q*r��Y���:V�74���2v�ɹ�,���xtd-m�2�MHa�3���u��D���6%��i~h�.2�M"��`�ղېɡ�Ύ��4�b��L�q�ܒ�za�Mǧ�tIŸ{`�؝`�\���x[?�E�=Q��v������d�-a�ȇ�X�����b���ϵ���3mN���� ���<C\��]�т#�n�eљ�c�� ��C�Yɖ��U�uN��v��	5jj����f5���kN��K�l=�Q�tz�����[���A��mr;?�N8+c,M�|YA1a(8(���ؓ�{E�+=\ǛW�|:�)���}�M�P���o�@z��
�f^3τD|��vw��va��l���8\��(N���^�U9U���pLo�L�g��� )B�#�y�O�Xҕ�ڋ`?�0��c�"P����BD�o���8��{���T�/�ȗ+{ �7ak�Y't �sJ����a����g�6���_��
����x8�zƶi�"�qqe�E�+�sd� 3p"����P�R���8�/@��i_��[�d���r����οb���	���	�*�*�i�xz`qa߬����b[��WH�Y���.��7��4���\�:��F�%V�'N�>��q�W4l߫<�VB���N������w�M�=��d;��f0�Gd�����o�C�7��֤��B�۾��@fgi����½����vv��G��k���D�f�9a�.z4>�Q�n������@n��ˁeD H��JE�s���02�x���K���r���n�*�9m;������Y��*?�P�)ᆔ_���-t���g���у<�yKN�<^�N�G#h�Ҥc�	��x��*=��v���}$B
���w�K/�n�b2/�$�|��H��2�'<�xB��, ��УM��U�^Ib��n�2Kn��dbr�w��"�2�Š�{UF {?a��3O�A�-��/	�ޜtc��m��8B@��1K�f>���~��7��H�dc�x�]����?y�+�X�~4�O�w��;I?A�>�6N�i�?4d�)6ʀ+2���#�zU2�jL������|0MW���eO�Z�p�G�^h�j����~�b�Pi�jK�藆�V��$�[��4�,T���d����xTܵ��4s\sR�Ev��x�>��<��|\3M�z��d�\��k��_�Ἵ:t�7 @��wc���N&����n�E<���SQ��ST���m[]t�d�-�*`B�r>�F�ǝ����uA	��̏��#�$�_�b�:6��Z�����MH����蟤J�k����$S�2�դ��K��Mj�P��%�>s~����Rg��BN:L!�6!��g<OU���G�!�=%�1e����o�-�����I�(���399�������jYB���)SJ[Q's�)�9,^��͑1��\�r��F��X��X}�߬���P�����f�p<م�z� u�Si��e~o���#�9S1+DNh�X�%��"�r��\S0��A���:�;���sְ~��L�����)���=drM�A1Eԁ�~H�N�ܤ���:ݨf)�CmDAY��[���z���߿��<���>�/���U�� �Y���[|��n`����F��vq��:�a<��p6�㊹dt�čɼ&��-��L�/S���Yo���m��܃$0^O�R&u�.����_�-�S����ת�.�����J,�8�6�/�x;A�#Zs"���� �K� '��@���Y�8V��e�@ES��H~ c'��i�!疾�I��ź9R.�#���3dp������\߽����R SӖA���ɓA��SG�>�b�&i`���]���7�G��R�'�O0�]�UR"\}Wzm�{d�W��TN�+D�uM��'2�yy+r�$���?Z���A S(җ��1���Oi{�~�:H��8'�jg�x6�Q�X��fBTN��s%�xaz�A�� �%޿�$��5S����TC:V�O���U�cړ���]<%!d���i�0(�d����kꓚW�����X���`ۙӃ
�(�-ޮP�FB�{��"�:ܼ��O&kO.�O��S�6��ɵ�wJ�&��Z{h�����֥�y�e�I̯K��f�w�*ȫ��j�0Zk�TPz���iʣ��y��y��6i�px�xQgʘ){����ӏ��J\[�) �j/t�8�YD��׎�_5����(m�"��ٔ)���l��� D^��D��b��oI���
���D�o9�mw���tǙ�K��b�LG��\�\]�������Oů ��Ʉ��!14�,��I㩶���$�<�rv䴡���'#�l�"�R��`��ŚQ52	N.::�];B�[`#�2r{��ač��ڵB�h���ۻD�����F<^Ѕ玝�dY�YK$�	wcW@L����Wo��y�d6��1P�C��?z���jc)��iV3���H� �k�ج&�U���S�v�S��]=�	��:� ��#�����1q��E��C<�>�Skk�8�v�1���1��W�D���B/��l�"t10�2Ƣ��#��:24�X`f�S�j�����B�~]���*�Ҳ�M91� �8^���p,k��r�A��\sCx%����ۻʵ���6���*0 ������6�7sʹ����$����1/�%X�$:FDM��!�4�\FF���	�[��<��ȴ��묉	�(g��KK;��.�߽1�}4�s��wY8j(�-�Q��������y��������Iܷ����D��^_�KEg�s�1`��:/���:O�6T/��V4�+Z�2���_e/|��EK���AY.�>���Ò��a1%x *Z�p��UAZz���`z�t:�"6�0m�h&�,aMV�?� �G�,9*RC�1���K  wm�DXoCa�z||���m���&����N:�ZlޯTZH'Z)�/_�����roͬɱ�lH�3rc���5��Ϲ���+���)}��P�>�G� �8~뢔�](�Hj��ڴ��I4�=�gnԪ/&@c�>svN� ,�-)gk1Sq�T��AIgU��;�{fr@��C��,{w�'�w�h
W8�!J���<�����Qg��	T������l��=�'��)��v���1&�g�|Ĩ�,:t������cL�S��B���`)�ڛE�Ξ�;8(m�k�r���*��E֬a+b����DMN��j�����Q�o����|͸��[8�Ys2fU����6s%Q�5pD����x��k�cm����W@��
����D>j����ח13,&'WFn,(�y�{q�*�ϒ��m0)Q/}z\����t���/`]vL_�7hyUQC�Ŏu��Ğ����/UDK�������������d"��yk��9}�%~.��	/ _�J*H@�k�N\�� �N�c/*�8��ky�nbl�O���#�wC��H4W>�X-;r&z��Z˸�J���Y���j�p2��s���r y�XzC�=?޶$M�o]�HF� �/�kPu}�� jd��;�[�k��g����O�}n�'� ���f��p�i�"�;4��/@��g��CEN��eu���ď�ʈ�~��G���w�(�tl{�S��sw��.�o�����S��Qd�EO�(8�L����Da������L��aځ�?-KzR�뀬u��n�p�Y\��ҙ�.a�32&ߌ!�AC��%%�]]_W�����-%�A�~�n��0��uA�+;�1k}�`�=W�%���Q��ԋm��7!���gƹEb��-,⫷��Q�_�ÌV�EV�s�	R��rr�Q��G��d����W0��꧁�j�Yn���t�!YG��W�x)��5֡���3(��.��ا�t�#�?�]�����}�Ug)K���BhG56�8v��5#Q�	�O�<#�-½�;�ȿY7,&��H���y��n�п�+���=�L_�@����|��f���:|��^�/?*� ���Fb��4X�/;��A���Y���v<E��2Cl�����;x�2�C��a}м����H�Ki#��ޕ(���bB�*h���Y��˱0�����
m^AkwL�X��u�"_}���F�:!Yi�Ώ�KL������o�M,������*��]5cU`Y�Vv`����<�||�$��7���&b�yA������V%T�!&̦�o�5������'M��"x"��1���8K&E;��>����\WاW�\�&�fX� x�	āJ>Xg��c�Q� x�ۘ��GwO��6t�jD�Iq���'��f�)S��u�l��t��!�ӥh-�|/|X�$�����ܾ�]�"�mV��z��DW���q w�<Y�h����B��T������ޘ�F�@��jX��I������@�������6�΂��Y1>U���z�~��s6K�����|�u+�i=i�W\I�<8�k7��5�p�8Z�懑Z���}N�ӄl��iZ�Q�,�O��BB,<�ju{.�}`�rZa4���9QH�5GR�H��4� �揮�4��f`0bZ�D7�q��b.�i���w�����bjOY�?17Α�Aæ��H��������L��w���|�����!��v~ruŇ�B�����{�-�\!�fZa�j]���򉋚�x���H�t�����A���r�OZ���X^�K�����]wW�^��$v�v�SϜ-���ɇf���Ăz&�jҹ��?�!���O��.�K�V���jҲ�'㚔N��e�>kx����YZ9I�vP �l��w�Y��"�����x!�3 2K��*o�%K\f�G=�-%��G9X���tm1E��n2=�-��dJ>1�;�$ǖLAEzO)ˋ:������X�r����0�@�Ӏ���_��iy:�GwI�-��:fR�5�r6��0�&�}+��ǢW���O��IA�������T1���퐌� :��y�����M�˄ҝz˵J�ӹ�����[伊b�U���iz~���eoD8�;r�0Ń�1I˚|~�~��ΝɕWWOC�oe[V���u����3��	D������7F��o/���cD���7�S/�/�
kI�;�S��t��N7բ����cz�h�:�%2��� U�B��_�?�$�@T�>��{��n,�ђ |�N���gJ�W��}�c��)
���պ���R{'�Ձg�aÉ�d[f�{!�t�D�P=���r�XyOs~Q��
L9I�x�<��Z���%��X*i�OGu�i����	+��l��RfU���ê؈�=h)du�7po��DU�\̴=-!�|z<c�)\o[a+�Կ�ˡ�g��I��
J����"�]vo�:�we��,��:��V~��L,������d/�H�箤�%�9�7��u���r���t���em�/���͍�����G��
u��0-�,|�C�Z�|K�3����Y`���-f^�8�h�Zg��t�:xP�(Hck����a=���xi*���(�$�9%����-i�R���aeDSgl��,|���㢓�*\��M��>"��E�R�D�,|.�b����SΚ���SD�3h7�Q��X�P9�^�[�Ks�o}������]p�}�dD����]�q�?Qk����9����<~ŧ�>(d��U�L�&�f���;�c�m>a��Vj׀���QJP���`�oQW$�w��E��mz^����M���fP��j�qmu��ׇx����Q�#ʜg����˴�Q���`��z�<�����5�C���r����7�F�ڄ��D�2��QS�h��^�]�q��o9!��(�U�vp.re�M��)�p���w�c� �\ߌ����*�J�i��ps� �^
���'tR������ �"��n&'���2�vqn^��^���ʗ��  +����Y�)X��_��|R$�,LW-����o�E�;񎙬B�s�Tю��O�)�B�G�h;BM=u�v�����iYy�o��d�����Xa1]��+j@�q�?��G�TvA��@�˃I}M���{�[ �F
<��%�F���-�ӣĔpGj�:�<&�;���MO>����0���b�3w�/�h@��SH��k
ĿYEK*��Ɂ	s�V���.-�k�!�I�
!MYȽ-������"�t�k�c��=}7�,�
aS�t�{�hh��8,~�;�76+��`O����%��f��Lߴ�G�Td-*��ZPS����#}fKO9�â�Vn��,{Rx���^�TP�(~跛`��yp\)��}x�� ��
VX4^*���c2��b��}=b��#a[;�X����({�����rc�SjT�O��tڗ�s����y;�,��z�|!��dQ�q���Ɯ�Q{�YL��0T@�3|���u�ݥ�g��v�R^4�o�����(��>(h�o�7�ط�8i���������kn�$����yo{Sֽ�$�t�94lNV6��
iT�3�9�U �a1�� �J:�w�0:���߀c�� A�����	�94��D ٔ��C�^��Pl��D�`@��XY,5G	5��'k�J�A��Ƥ���'!�06L ��:r�X��* ���R)�_�P�%Ϋ�T)���l�����fuՉjC�W��2�����;��ҫ4�A��0]"��p��a��OZ�^�t�̢����;���Ɓ1�Mǩy��:���2�0d~�
�r��ׁ<<9�`�T^U`��� �!�~}^L�W2#P���A�DPҥ�kE�}�e8h���cTy��|�
�%�H�t�^n߱�Z�����>�-lJ�) X�&[�LL<�F�cst1�)�T̽��U��6�@o]�S��m�Eƒ(;?K��А;���Wgr���L��-W'j�J�:2M�ar"��R�269��CLKG&��Ǫ�)�������ZF��`���~�%�+��D9nM�za�����6�(��S�l[�G��]@�"z�չ��	䧤���DT��)�T=_BXd����Au�hf�7��<G��&	�X��a�^r[2��4K�f|L��/���Ԫ�y��a�#����F�#��"�����X(ƌQ���3t��=Ϸ��dIR��9��	�G*�O���� lP�}��^r��lg�G۽"NE$���vs���1Z.�Y�K�%���y{��Ur�e �Nœ>�'���V��%�$Dc������==Hg���������[����b�Һ��}}�ě;-�P��2/{�I��n�v�ؘ�2N��v�Wi{v��bY.O����ː�s$�烒��)��h3��t�I�Yyȧ��+*T"���/
��#e�?~s��]�ΐۍ9sr���y���5��+Du��U�>��Ŝ[��GZY"uS��݋z�1݄+ g��e���P~N�|0>6(:�ns^��UW�9���ͧ�MM�G�y�1��G��K3ѳ�r�lBT��͝�Q��'���n����P*�������
��j[s)`ٱ\��?������E��a�C�"u���;G�D~�*֪��%��l�����p>Ү�p��n��
g�ѷv�/}V�d5�T<��� ;�;I!R�6Ǡ��C�K컢j����>�4�:��TO������O�d	7I�w�[�HAXw@�Z_J]^c��"9�#޸��˩C+�'��Y�c������~��;��+�H�ĸ�{M�*-ƨ���H�z�VM��(����<��,w>=N;(���W�� �^�r:ml�6R����7͂e����9�bsL�r74�+,Ł�dg3�y^ �ͳ�S�ܹP��u�����v0�<d6�x9i�U��|_E�P|�I����֛Lp�"�������<�0��}����y7G�3�_D�����Ɛ��)T5{g�|�����Yעe��J�bDY�#r����<2@`u�=�&Rj�4�|���Hù�%�������M"��q�/i�~��2�7���v��d�k����[�2"��qD��ڹד����@cΎ�A���
?�fe���P8h�$K\�����!�yD��u�O��(�L�����'n�@�����S/���1[ݗ&�s��z�`j4"�e^�m��e������U���>�������~+��Jy#q�U�#���!-"�c�綅k�fP��bw�8����w7�2�9@D3C�,k�C�?��+�P��IqW����ⶲ�YZtK빋Af���o}߀ԧ�ǃ&�^����ܽ�-��NF���a�bW-���a����ḯ�z�8�*���$@�����؉�����ó�`t��כ������ns����;DA7m�BrC
��2���4j䂝nj];��� L�p��d�*"���F�~]�p�3�ZO��<�2��_pB�q�*ԏ��;�A ������&g_m�c�x'e�$C�y�*�)P,s'zi�od)u�1cc,�''��t���){�1hL�2N������R�M��\��-� [�W}�Dn�5׸[O�om��ZÍ�*�M���˃)�
�����˱reaYhO'�#u������oӸ ��꒯��?���uG�0i)��2�t9I�R�Wç�E����������/�D �ɛ���G��5��6�
�1��L~a�f�ѝ��+`#�G����eW����k��GN���*�!�l�"�[/��>��c f/C����� #��蟥ʵg2 �2`�u/��$R̖��p�R����'.��x&b>��S�e��3hp�� .�Q��� ���T�a���SL�r�w���"���0
�Y	�hCteZ�^�f�CT�9�$L��soLi���
���|� ���3f*�� 1sآ���ϏBs��)��}l�������hW/�&�"	=2d;�kL�+Te;�e��Z���g��9�e�El����uOǵ,P�� �w���#w�(G��ZN�΢���9��M����/}�
iag�VFt�
�K���^�ǩ��B<[�Dض�^Ҧ5x��	�J�u8c�p���|�X'��Ts]�����:���	�â�	��ֻ�X�w0L�mjK2�y�b�w��\���	*�h:����f��T�F��O|���F��YD�6�LϜ�w��C�
���N�{1�&��t��Gb��������>�������bv��7`�¦$?L��xC���!� ��Fu4�߬l��kF���m	��_/��j����_ť8�`o��<t��J�wP���o�5k?�����}��FJ�yz�������%��T%��?�O�6Q���i�mZ�O�虹��lW��e��nF`sO����#��'bj$zz�t��5�w���F�w#���ɵRV�#ڬ �0���1��`��l���xJ"�<	D�w��y3WQ�)��ۈ����]�+�ؾ��g�+�W�iԪoRC�\Ħ}�u��*���my�#)�d>NB��>�d$�X�$���K͞}�"�]��L�B�U��XO
P7�DPA
?�`=�:���yfp�&�;�:�,��*ϟ��$N��M��=���o���()f�#6�4�ٔQ���M*?�tA��"/v1COQ�4�zm���ĪT����:ˏ0ȥ�.u$����{�)���"�&!D����_՗���#l�	��3޴쎮	�
�����5��D;�C%�"����F�H�	��N��$^T�GM�i�2.Mr������GO�9ҳm�H�e�����v!��Ҽ�<Ԕ)�T��� �,�yw�}�����%H+9��S49k�r�.�C�z �ת��&S���9�؊�;�}��+��N`�Κ$���WR�1d�^2����C�*=��I)�j҃��
Y�R��**u�%���|������VZ�p�Z��V5��[ӚDQ����D_;�so��qNmgs-�Q�$���P;��-E��{�e)U��۹�xZ��,m 5r���B֮z�)��^�A鼖!�ބ��BRmg��h����JcF�l K�^��Ĕ�j3�ߑka�௰|��q��Aƨ:d����5�l�4���*"2�ST��D��MOl�	�B6��"�O "Q8����z�^F#m��bO���<^�Z������$\~�r1L��V�("ԁ��[Y'I=y'_�w����h�I_�ߩ^\2�XP9O&�Mwy��E%;L��|%���*�e�[/�)ג�l�����(A�!����Y��U�|����١���x��Bf����.�#�v�w>myPتI��u�jW�NBM���ǵl��,�G�yif"���ޙq��
�L���v�������d����)$�@`j�Gϸ�^6�p"�g�-�~�yg��ks[�2�~��,fv���ݕ����i����Ht�;�X�B��ʴ�Mٮ^��V�6/O���������Y����H���Gs?�q���
[AÏ��Q���>��h�؏Ce�j�[�]�~A%ks=�z�$��i���}3N�{��}jl2�2d�~��Q�� �Փ� |1�E^��K�ҧ	��2YG�{�m\ ��^r��άPTH���v�@��E�"	� #o��Wd��;2w_DfSK�bN���zs���Z�P�o�V��z�H�f����׃Kpn���PF�p�º��	�毠3�.@�pL��`Ͼ�s��wL���c�4U�6;��}��EZ�@�GW���ws���G^Ⱥ���E�j�S��������=��/|����e&/�d�"��ʆ?�k�B��bt��Vj�9y�=6:
��D����[�tF<ZAi� }�>7��m�a���L�"��o�Jʩ�/o��w@]�L�GW�yw��r���]�U�`d���D#�	�Z������h���ҿCf
��~v޵k���dVt�0����j� f'$�\e�y!��_�D���0i3�{pԯ�W�3#/L���l���n����K��%�a.�������C�28�hև!+���Z�!��lH=�dy�R���������zin���/��!#b�vL��ۛO��ڽ�8?I�ռ�AgQ�3J\��s�	K�Ǽ��ET3D��u�z�!��|++8}E2�0 �?#,��������:�?	囨�%�ߦ�1\z;�,����qo��ԑf�e<�ޛn�����8Q
i�ߐ�kk��jk~O�'��c/ӥ���xj���h�sæ� �⾐���aj�[Bڋ�"��Y�J���f��8����Բf'�RdH0�e�~��+�:qM��ɵ&��~��d|#�"!=�l6��,��J��14����9m�!�|g#�J��.ޭ`3�ֺ�a��-q���VnD4���8���M�k�|m���^fRǾ�*p��X��ǩ�5匳���������ЩO�Q�sjf΂����2�B{V%��!�3Ь��)s��@v-���4�[ [���N9::�s���4�$����tL1����ѯ=X0nl��0`o<����-T3|a��9UJ���[��pT����5���,䋗��$��oz��F��U����`�j+ߙj�*,
��u/��?� ��Y nav����2[�Q��g8���l�$S��y���T�7DY-sy<�iՑg1���N�-����&V	k�e	ϥc��/i%�*��p����yV���}^���:�O=��'t�����60���o�b��a�f��]w����4n ,L�� �ʍ}����F	�[z�QVs�.�ZS1#޷n+i"%/��Z�<�f�z�`E���6�ՠD����W<�����˅7~-�Z�����BhM�W Y8�(�f�m� ��"7 ��	�Wx�I�Dfݦ�su�ݹSF�����~�:d=����Tx|���&�g|l󡛓)�H�"�9^t��Z�]�Z5<�P�s~b��i���G�e/�9R�Z�oS���l��N"���'wyW<{h����Hx��k��ၹ��X��5��\���*
�!t�E ��d-�e�,�-�,�|j\��V��c}�L���3]d�?Q̪��U
#@,˵nڦ=����=Pj2�]o� Pq�Vr:S�O�$�L�t��0��2�Xj���So�_�%��2v$��5������y��3�kU-(HoP���7X����	D�*e71&!�����>��q|�:��e2T9n�5�iv��.�G˥�D5dq�ƣ��X(�g-kd:����+4Σ����c2�K\{Mr}�� b�]H��*�u,�'(e�f��_�3���׎;��q�S�̊I%2�"5�t��&4W��;>W-�oa{�׆s	l^�W:mLn�C(	7��A��oL��rV	��)�׷H#V��0&RM�o;ݦ]_}��j)�^2���w�6��`#��Z|Vjg��Z-�E�~15����Y�!A���T�C�t����}p˒�9T.���f	W�0�$�������z����kPL4z3.�=y�J|+"�)es��.'�;1�q�Q�9F-���-Z��M�Gk����X��"`����z�D4��Ds�i/�(ukC�-��&�t�כ���%]M?�m{~��k(}�*���v�F�v���M6i:D�H�*�-D7���o��	v=��_�0tZ����uuN\�����}�Xr&j�M%�6j��l�E���
{x��Q��N:N��D�����4f���+?6�-D�3&{p���ʮ+�:so'���;�  I��.<��	y�,I� ^1�}M�0A�����$�C+2Z\�*���.&���P�r,6?��B&�u���.Su�����v����me�_���a�B�e��� ��5��_��:�X�L��6n�,�ΰ��$���$�/0�ä��3����яӫi
�*o��D�g�/��1��I<�G-��o�������i���F��Q� ����If	���M��;F-��͖
���9��K�7g��s�R���=�X��&�Y� �g�Q��͍������|�8�t�G+�9��O-Q˸�|������en��R�O�
���s!T5\4��T�h±�4x���[�A�%ց���¸�L@��e����ܞK�c�T~���H흷&J���^qՁv#�us�s�f���"��^w��I~����A�q�U�����Ȃ�:V�����>U3�,&��}�˝�4�U!_���Þ�����#>���>*��x���k�(�JߛmQ�4����u�G���8�"�4��^�Zs�[�.�*��ֈظ�A���n"|��=��5H�W�%i4�N����\Զp�8�A]�WV��u��b���B��]mm ޴!��p�g{�2xhH;�X�؍���Xg�[��]� 4O���bF�����3X|�e
���xvS17\�; k{S~��GԦ5Cak��SFՊL��TE��0�"�~_�ZC}9��`<qۦU��a�[�MF�\(�겉3�	�Ơ��En X���/0��h%<�k�9�a��X���S�L�%��͠�'}���e3��6���nt���J*�e�e���\W�Aw��5'�
�y�n�Ʌ�B`�� w�Jg��9Ǖa��ju��/�G�q��Ub�a5�����t}��u�o�fq&�*F���WBݕ�o�D;r�<B
����Hy4�w�7�]Qt'����,��+g��>�.���e��Ƹ�Sh�!��&�K��톄G�5v��BTewi��q�U�
0=a5ko/�/�]1Z���E�8T�k��S�U�{����&GCL�&ʨ.jWTh;A���K��|4��	b��p��M���l*+����10t8��䕾��O�AĶ6LE�|�y��\h��O@Q+V`��&��)z�IIgk�|L���D��g��.{L�h�ˏ `��3=�,�i�{-��HE��8B��5�0�FZ>;s(�ď�r�ᤐ'�+(mp1�E6�I�rV6��@d��%�#rs:��f��i��bU
�����#��X"_P�8�/�kk�u<Xn5�$�yS��yw�-K>�u��RDu'���WR�5e����7�]-�v����Ѻf{��5gVjz�/�X��� �Q=�so�,`�1	@����yn���=>-�W�Ɒ�h�V�cj�U*�@�X��m��^�P.�ږ+ZN�j�p�F���ib�ҿ� K�E��#v����N��uD31S���4�B���CT���]�� �
��wf/#���]����et_��q�I�y��Ȁ�8���P_B�V��"yv=�Y&w�nM��"4�e��"t���j����Q�aj]�!�sGEKN0>�ؾ� ޝ���a[b���w�1���_��}t�"7�z�_j�;4�0B���I��K}'����bl'��8&�~!�E��4��O�g(����D�ˬ���G&��%����˜��mC�,ځ��!m������Q3�m
�hc���r^P���5�����S?h�F�=��>�J�5**[X-�~��bO���нη����J�:�f��zH�o1�DX�?M�E��_e X���ɮm�P���3	�����<�ˁU�Ѣ�w��Q{u`�K�-�Ef��,�� 6�-V�s[pH_dA�8�_�0ڮ�y1jǫydε��?�z!�4��p?���ny�@��VIb�:ﱭ��^����[����@�(�p�V�j�G(C�ܟV9R �l�e���������F-��ܫY5��H�uO��(��d+Jǹ#�'ۈ��a�ȹS��`,�d����@��+`�3� !��e�;�}6��8�"�����C�^�.=u:�2�j�A���1�#2gtE1,�<�	����{�Xs$�hN�Ck'�� ��)7�c���g|��t�u6�"0�%��׺Úy��>OPUd�u���ij��ۈ_�q���_���T��l���/��� �56��J[<9&~�3��yK�Nt��l<�%�n�kR)��$F�"�_��,�
G�7���_3En�`S�8�R�\^AD�0�h^Ğ�gl:EAY�����\��J!m�a'�`���>�7����/ut�Y��b�_J�����F"�.�mN{���@���va�-���qA�\���Hg�1� Y��t��%	�w��Ì�C"<+�y	�i��
s�@*-���vq���tI�ɴ+�� ���˛�G�8^�2jiB̀1 s�� ����Pq
����B}�qG~�M���*�H��ּ��x[ah8G��ٞ�+h�!V-��ˏE,3.>�lo����h��4�Mԧ� T^�0 ���u�g��ԫC?��1���P��|^���E�@�ה?K�sY����N�6�����D�������~���/�HȆ�<��7��c<J7��e��ĉJ.�W�!� ��~Ō�Th{$�5L�bCK�E:9l�CcK�}zH��Yc��l��@Qվ��T�Q:�#/1`�Ӫǈ�\#k�ks3��|���d��gI*��Q�G��	��7�P��V��
��mY�p`�[��:P��R�0���G��'ޢ�8���V�Y��ET�I1����� ���\q�g��G����l{l�_��`�����|�Z�!\�
{;���j{qʋY���¤��>����It�T4L�#*~`�\/$C	&�lt"ܙu䡿����ha0�S�r'�6[�X�!4}��N��R o�c�W��XV!a�Ң��1t>�͚L��Of�u�6�eg\��O�����@�`-a�g�g��^p⏪�K�mYc�G�-�k"���=�+�Q�F��84;��H<�3���v�f��vT#9�z�����T,W~<�^B�����[���O]t9P��K�%����4�6+�(7BC�4l-���A�v�"�L�����(�07K��nv|�� "5Fe���\�P�&Q��t�@��!�U,t��7%/��K�uz5B�������e���l�(0�;gΔ{eoa�B���5�J��}7��L���sfs����ʮ�XI�"�Z��A�tX���Clj��T�CI���-,V��\y��ZOq"����a�B����\�T�Ã�\��9x�2�+��7L:c敞��i���Z9�?�i3�����ڬ�+� ���,$ Ym�9�o|[G����-.��k;�#���'ګ`��"�4�9�O&�|��{T;x��e��7(� �\+�G�s���N�hd�SXoTwȔ�e�*�L�����xWyI�Ǩ ����H���cKݳ���!Hh��v�_���?黎�j_"rl�EF���ޅT�#CtU �q�>���jJ� ϽUV$�
�mq�츓f|zM�/�.?��Wk"{h�~����R��S��jm�1���ίW�E���B�����\_��Ez:�R[�M7�,�Y�����W{�f��PQ���ŉ+֑6����K��`f1ݿ,{Iu���ĉG����\$�8#�֏�{X7e\�ϭ�6��ci��������lwA��d���S�$u`'��e��>g��������S �b��9f�t;�do�u���f�0˛�	�%y��J]�%쬂y���X+��/-�S�mN�/��M 2�q�p��b������J�/h����]
���B'�s����r��A��I��ֲ�*��I�����^e�r����aL|ǝ�D�!��.�ow�2��B�ʦ���_p�����^�~�4�,aâV�$r�J"a�d�
�����Ҵ)���x�&�'Z�f!���ąS�8�	��6���Iz�tzn�?M������ݧ!�ơ�.�ϧY�Ha�۸���j���C�d�+��ե�%!�l�ς�:�M��q�2i��≎SR��~i� �`!�3�9]����SLqk�Df#��'���aԯ�W��O+<
�d��`A�Z���8 �,�H��vlR��J�^��3�w!��FW�����C����)[s��:!�����Ň�^5�y'��7d�>�))��7! F%}��GD�)��1 -���C���F��+�ކ�jt�a���0~�鐌�`6�1��]P!��:S��gJ��7o��x<�[T1��/�bBT��ξh˦������luE�P��=%�bP�v�\f�݈v+�Qh�4�� �3S�� ��p�~-T���Pl%���}�DT� ���y�N��O�[g����º��N�>����h�C��ɸ}GC�M)c�>�G������G���ҀfS�i�2�J	,�Q�P�k��=��V�O�B�6T�?�>˷9����,���ܯ��mk���\��\|��m�=����z��dw5~S�/�W=�9+\��G�7�o��-$���L)�r/��F�Ҭ�=��ā�`̢Zl/2^��E�p��ɀ�/u��1��Y�kOg#���\s�Q�x�No"�桡���\�&6�8;��B#Ϗd�к�|���ڻ�Vߤߏ^J��2�%��w�1<gD���B�~CU�z=�
�1�z�z�L��(Jmp��Ɠ�8��p�v��֎(�ﯶ��1G�_�
�	P�;ʘ��p�K�
3�؉T~�
"�!KC�g�2��Fx]�1#|A���� 6�\P����������`3��q��BFe�1u�̅\$É�B��b��,�i�plx85o1�ȑk}�/U!�I ���K�I��q��y��z���q`���j�{q��hh�P&�ӍƉ��W����WUK�>d/`���W��V���������+�Wm[�g
�+d����󚄜�i���~��R����_ɩX��J�qlwt�lT���l����+^g��%�|Q�]�K\�x��J�`}�$w3@`r��$�<��B7~�9�j����a��Q
M��t�x�u��	���e6�6)�/ZcP����a�ڏ\5��鳫W;�R���� ��w͚�
7��H�*!`�GG�����B��g��h��%V���y�v����\���0��k{n� X��=�:�D�9F��kDf~��J�w�zx⬥��a!��[I��\��سu�\c�������g��c�C/��1L���� :����W�@��K�r����mL� ��im)APm都+2Q��s�6�=��X_�v/&U��{�k�\�U�8:��z�V��T���AS�b�?<~��C�)��VƩ)�k8��8��{�j�ů�ahY�;���O<�;�K�D-�'�,(%>d�"��OƄNqa�4f�E���� �����ֳ����Q�U�rѴ)X@O@�M�7�Ai�N��a���B��PR-���Ɔ��7���Z.PFZpce�H3q�M02HT0���o��O1��葅a����O��Tˮ��p�9�&����@`9�(������B{r}|�PGl(	��픡6V�k��M�{���eo�6m��˷�Ӷ\�Py�ڎ��5d�}ꯤkXx9�|��4ȼh�ǐ�8c��t��OCN�zI �T,�?K��ƪ��549F��u},B$��E]��e�"��i\��%a�&
�
��#���g����һ�������z��6 @�ڔ��N��F1�{@��K��F+m��G�����3���X� W��V�r�Pw�%���Z��5��[s�c	@)�{��h�t'p�h��-���Isr���(�e_���Ӱl'1��Q�_��,��^"�4��}b�|h����%V��m�qH�+>9Fx�S�M�� Yղ��3C)-��2���@車 ��iCb���\bjo����)��f3��i�������p�V>���`m��? ��5}��׳�pw�+A�5�Q%��/ǵ<���u�٣�8��ߑ%�� �a�}G�k�l�%[=��p��
)��ӄOw�kr{N���j�::�W�xvk�+�#�l@%O�hw/�$�&��3n����D�p�����%�K6�6�_�qB�^��TTn7�s�"�=%-���	��8_(��9ʈ��֧]�����kG���ف�����Q����}�hߋ�������1�~[P71NMk[Q��J#�`�ȥ;��&�Z\�^����~�ϰ�(e|t
��h��c��s�<�3NZ��X_�U4P�e��B��<5�p��ҭ�*��fBI: Gı�j�����p:ڽ|2l̄��w� Vb��IJ��/�3�s)�n'1����*p�Og�zn�f��4��瓜�i��|Cs�?�j�|/Z��w��e���j��{�4W���-�r�6R�;
0��;'$Mw%��X�����5���(ubg��K,v�Bz��X{h���Ӡ��9��n0P�ȸ/.� &x��Z��&,/��X�O��S�˴���Sr�5��@Ę�a�y��{?��?_+�}�T�v��C�d�9$7)_�
<�����C�9�Q���S`U�����2�����u}�:��H݀�l0.*s0}���9��V0��!�m��S��𝛚�B�m����aDy?�^�\B`iG✤qA^���{x�W���IC}�F�l���N:�%�$>�`y����z★.ܧM޶:Y��qўS��)�ƺH�A7�S�?��'y-�����&�yտX���\�Gb������s���3C}X�_�6q����p�`!SV:I͍��N��M�㉄����W!Mtah�˥M�0�uRJ�x������5TPm�=�ȝ�\�cT���]H�I����Xr[�(�Y=�<9!�U���	�B�ዉBS܈)��+�d}��>2�#H"v���׌�{�җs|g����Z�v=���:6�$��hm��O@��W?���Śd�fEQ��Y>�8دߺ��D�e�8�\F�6�!1'�A WB��^�iLv!єbOrs�T^�{�Fj�8iP�Q��&�l�B��K���L���U�����ԄC�:�s%���f�[Og��k��Vl'T��3>+儓��Ԟ���="W�Ȗ#<��IyH1j�?On�Ɍ�3U�M�������"#}���>�yH9_��5^��7��|o�� �mI�v�֬�p�F��j��8xw(���B�N��@󠻂��?��z���F��� �A�z�Tk*$���*F�0���>�I�U	�f�J��$؈Y!�8M��'@��A��_𑋼�g��E�̓�ɫKG�T�0�UAD{���"y�����N�b�j���_t\�S� tgJ,+��X垧7��3���V0�C�2oX4�2���W� 4:�p� m��d���@]���LwƋc�S�Sv�#I��Y���7Fx��,�!l^_�ʿ�OnP
�T���k�f<��o���*�!�>S
�u�V5���)�?+Zǝ�2n��=N�LV�!�o�h.�H�	����`�A�bG����Fj�dLцPE�;e;�c��.�d���=}u��"��+	�UB���aU}驄>�5DR����B���D�� a�Y�ED;X�ӟ�-��H7���w��3�B!=���c*�/��2���¥�l'M�A�<x&���R��D�Ķ���&Lt��̧�(�Z_dA�\�X{�(�����}�8�����Tj9>G�[%�Ae���m��4��o��e�m�M�ZL	�����.���_)2�������v����/��AB�=���F�ש�g�,_�!A���ĘND�9���g�-�+Q 2���mpH.�dp~i��qpI�����p���K����1W�����Ŕ+�ߑgk4$+c��h��7��vI~��8�}�l�N8�!��~�<�!����Y�|6��;��e�Eo�٩(Yr1梛G���g��ޫ���_��C�O��	�BUYi��@����צM(�h¹<�֞�-Ly��Kp��=�L�C��yH��$����9�v����&�O���]	-�*.߿j�0��{���g{�A��z<�����UzF��y��2�*�^����W8�=��D�g6�2����*�7��0z˔�s��*�(�$���-�(��YR�$���1n�f-����)�;�)]���7��nɃ�=���(�]�8�1{���+�Tm�$�g����;��뒋 �U��
1�i�������LB�A��Ӝ3�y���,�R�X
�R���cw�̨�P�$I頊9q��kb6�{
F���na�.��~�������'���@V���5�i�E�[w����}{9;��n�
6Cޙ9+����g�����9�e���@�<��:z�<Ƽd�͙����ٗ'U��$�(mEݬ"�Dk5m&��_�\L�qg�;��E,gi�~@�{.FI�j�'l�'H�}�s�h��ޖn z9k�>��X���@��ӝ}~"���9�R�~�^��&�3�����K�Ω*P�Ð��wʘ�hY+�/���n?��R�CG�p��=cS�oܘ9�����c�� T��}�4
�|��ڣ_�q����F�'C�Raq����k�`*W:�
D���9 yH>8����y�Hl���!+l�&����p���l$I��30EIq������7h�qF�j�S�D�����J���"~�L8;��i� �����fٸ�i�/�i��t<�9��,���q y;������'��������sDwo!.x}1��������^!`N�`eq�hء�B���ک�����#b�1s���@�z�*xX�ז�fq|�u����
I��069vō�R�v2��b��=%ZM���QQ����kX�٘�%��n�K�Lh2�W��dO���uhE�)MӍ1{��y��/���З�6Y��P~�k�O<�<؊`)�^��_[`p=+�	�X�"�E=�î�1~�z:]��z�5�I������I�mW,u�GA;�1x��*T��v ��\:O����J�?�uq�ˋ����oWl�������ﱳf�,�K���r�'1��7��Y\Ϡ�)���ȃ������T��4_h��5�o�Q%�l(��U?�Y����C�<�N�f*7�����'x 4_R��?��ýv-r�����)�3#�a��F׬�ƽ���;W�m��<���
Q�y�'�5��� �t��D�d�X�k��G|w�6�1`�G-?���o#�K�
y�m4t��B��/����X�Hy<���}� �tJ(L��
�TmN�#xD����C؄gK��˺���QQ-�g���x��6���7F��庵�O�mR}��	h0�Q>��_���Zo�QD8��`���2�o�!B����P���&ASah���H��g�V$��tF���� ��-����<�_~���5W�t���}U܌]z�([�vD��
\��eB���������i�Ӧ=��4aI�1�q��x�$�R�� L��:�W\����K��[��ϑ`o>\,钨���xH�mލ��O�kv:%~{WH_�k}U�k�~�e�(a>���N	��l�q�c�����!cs�lfA�X��j=ޑ5���c���>U���=F�cM����nnV�Q49��!�:)FW��"�2�띱۽A��{3˃�p�"=AG�א;|ٝ�gW�L���x����W�������υ��Q��i��u��g�%�[Y(�-HA�I&��m�t���)#6�ܢ�`i^�{C��M6Kl�[M���X���:�?�tog��8�ũ%�-%��s\g?g ��ePS�w��#�%�&I��eI<����pluSG�f:)�w6��}����,��_0Qa ���m�y8Y�7J#��6^ ������%'�_@�4����$M#�Z�\`�0n���/�a������2a�M+�� ��Xw�p;�8��OjGc���;��p�.yV�ga�2�mK�����&����ͩ�����&p�S�ґ��&�Ot��cn3L���EW9�w�.�V|D�}�ԣuw�gp#e>�m�C��[�Ǚin}�7Y���'�e^�����C������c��tBcQ��h3H�1��'��3��ܫa�8�NG�����,�|�';��c�y\��(�`��reN���C>L
��#�6�8i���3*z��Vł)�-S2[���=��<�Wj!�%K���uQ�\p�K"˿�/��(`u
��.�1C��7ռ�+<.��A�u|Ҁ�#��\ɮ��j�B��j��@����~�AU�D2� �馏l�w�"��c��؂c��[p���DQ[1����,�����)�?�Z�[�,�LD���$�w<ۙ��!�}N5�5ӊՂ����/�Ƒx�^��X�����S�6�e:�9&�<��4�A� ��8Xg�W����|�����%�*���H��7	�����w�����A�:SQ���_�V�E���d���n�+�$�ly�P0��t�ᎤI�8���6&q"U��k��^f:���7XssC��@4^b49�S<�&���NTEt F+����Ѳ}9ˑM�?���nz���:�<ः7�9I/�i"���uC6K�e��2�b���"�i�[�͞�*[z7S'�=�c���/^`t�,	pTc��}����$6��]���ի�J<���sEߏ�74��q:c"VTE<��/�!-��~��L3T��Z^��n|Bw>!v�ɓ�7E"CP��7~둠�f�}�)�*�xC}�����#����%o��7�Mm2|�n��Ě%�Fuj�R�t��j��Q�;L�W��0�"Fs�����a�a��/"D��������o_L�5q���@pQXp��ĥ%�_DsK����q�xCژQ`OK:�e�8���n
�ۖ�Qm���hQBɭP�"l�[T|���g|��=�c�.�R�8����|Z�4�S�Ҭ��8��� �I��8���&�v��"��Q��ag��qX���r˴���[���4!m��q�E��FB�9Y%�y��J�L���!!�kO1@xr�4^��j	d����~�pD*4�f�H"K4���3H�����K�=*�~z׆����Og��Y`�F%��Z�7#HH�|z<5��������,[�Sϱr���}�e��d2��c�5�&gaaP�!0q��ّ�C!9�HH��B���m�_�e�VA���ղ�E.k�x�;��{�t[*�`�:��|�͸u�!���
�:�I�'��������37@���b�ʿ�t���'��!�
����c����GqI[�~ .��6��C����TSZ��# ���R�����M�Q�����n���p��(E�N�a�MK!*�
&8n��;t���Z`�E۬���d񠼜(	�|�ܮ���1Q����I8�_��8�_:���p��|_k�Qf[�D������!�ٴ��P�T���Gj��6TEW�d��+�;���U.S8>�j[�Cn�G��?b�#��C=����V�f���Hq����F��\e?:W���uB�F���%����a8�I�2��6�{�2��� A�q�e��/=`F�b.}^��/��@𞲉��s��/ݫ���U��wo��y5.I��(���'����KD#�K	�,.xS�||��PU d�3���`"�W*�f�������&��[���;`sŨ`)�$C�sB_��/s^ͭ�Jff�X�&����)&/�@.U���(%�������!�l�v^le��C�o���%���]����`nt�^�`������[�ǫʔ$o�C������&�ˠ�'��Pq��$���T���d�t^鑩L\�/D�K��| pGMZ2)���]d�O��1RY�q�3�!��v2� u��6�0��(���*��ɠD��k��X�>]�RY���4EZ��������Q������F ��M1Uhb�H��� =�]z]�w�9���F,��")�(���mT���}�
)����T����8�q���J3��y^=����i�J�'pY���b�qؓ�N��<g�:�y@]���{�p��;,�+*���[e-۫��;SWݜ#'B�&���}3��
�����2Ǎ@�����&�6��Y�`�T��m���=�j�~���v��#���QO����fɳ��|r��pM�u�3B���bw�>F
c�na�v��.�� �g���*Y�tdk��`�#��<��KMc�C�џ��2=���Ș$��[nr(�2~�U�}ۨl��x��Q0�����9�Iq�\�j���@��*`l-���P�n�1����:��ȉp� roa5�F?��*��$KНy`}Ż%y�?�o���/;���r�ͫYp�7<�ϗ|X.���_07��,&5肣1쵞B��3�MM^Nh���O �&����(5
H>����3u)<�|��z˚$8���Q!_P�m)kQ
@I���Kݐd�\l�t@f�O��
��O/.솽v4��	>�q�s�����N@(���j�FI��Q�p��t�IXaW��'�ĺUh�1V_�<�h�⃡���'0��8fBE4�9(��G���� ��Yo�I0���ֺ�[^��|������*������z���#F#�����e��_-�5c{k�ʏ�cr���QI�j�Wؘ�U��CĖ8b���R�u
�W����l;�� vp����f�-��͊ﲠ�i+�&?y�:�~��ڬi��]�4�-q���Qi��!�eT��� ��ԕ�d�t�.%��N��"y�����g|w�01��;I~69��7T̝�<��([^�^�����~;����F�BU�;xXML^�K�@bF�8D����&{|M!��2�0~��CO�![��T�1��7|��Z��g�$5�k(��ɮ�[`�c��=�ܹ�����)��[&���T`�k�+�;���^�����4��`J_N
3�4xn�׷q��Zq��^�h"�<V��e�?�N2�hK~D���e���l���X㌥�7O��-�{��a�Q1��[��sJ&:�]JV���
��*G��_�ȋ�_�:�?��S���]�sD���N�����/�3tb�A���"�|9���WQe8�j̀���*s�JG���dc�V��-!��d(iߕ��Kl
~���jSV�4��~S���'te��2������Pk��Xu�2����#�]s���ڴ���o���iBA��
����1��D$���9s�d��������)��N�����G�'7�˭;�0��L����MF�1p{K>�P�0��2�v�|K��_r�%sn֌���ۺd.�c��Fo�: �v+r�q���V�pwjc�cO��Xݢ�1� �s�Ԃl�C�ʸP�>1�Uj��(�s(�,EFlPD>�6�/���ޥ��Lq�r��uU�g�4�~�ƽF�ѓB�z�JCž���.�Kl�	y�Q�_e�W��P]#��a�c�un�����T�bN�E$0�<�,JßS4p�^��/��E���ʀlg%��C8pFC@%�M���p,{�<�W
�X����jS���e�lX��/|)����{�����Ǜ3�F��j�h@a���ݓj��h&JѸ@��l�b�@:��]A[t���E�6W��\�5�GI�0��O�����CZS({�Q�G�㍄�:�M+Rֳ�aM�×J��1��*�c��u�jV��i!J�D�l��<[�J`T������Ns]1� d��.�t&��*,�Ke�}j�p�
п����B؃�Pp�'2���н��?^˦&1�.OKo@�x�������Eq��ϫ�\�z־�����5�wjc������0��0��$@{��`<����+������4��(i
t��G|��Ț@�A�ܜz30�1^=����x@f�+fֳ���=�N�i�"��*A�2/)6��9��;u��ܼ�Om�]E�ig� \��U6t�I�J�Ľe�V���e.t˩�����A�������W�S|��m��9sr�L��6�&�Mb�VH���\����(0�D:P�J�b]�M�o�?y�`�9h�mJ\�_��P�'�|o	����ܥ%����y`|ylR,d��oc|H�'�&V��QNy�C#�Zt��l���R��������bgt���x���������x�V�!��4��w�/�� �>�ղ��3K�\3u��wf��
��@���W�Q=C΁E�ၾj��i{�����U��A,�ܛř���b����@[ޢ���Պ�2ܠ�-��xϐ��k\��?$�JZ5�U!�r����<� >E,�N���j�d`tXt��GDACH��@d��0�c��ew��yW���SKK|�����=�FwD��&eH.%it��*�kfO�Xp�\W޿u��Kx;ˆ���ړE ��GO�!�1=��[��%1EX̞����+�U���w_����Z7)�C��ɯ�[�0|��1�6�.d� q�{�_Dl�F� *�!�i��zmXh�3�n����V��rPF���	i�2���~����q��`����S�cn��{����5A�^���3#�p���V4^�$;)zo^�A���A�"�O=�w���Su26�E�1~4P��b���J���zt��l}NQ\��Hki��0W�@q"�M�X�W�^S�r'�A�P���m
�K��c.E��I�VB5�8�<�"�9�4%����5������0`.;�_>�e��iO�1�>�%�,�y��PIq�)Ѝ�
��?��*O^� �]NoP�{�f@���Ą]Ԑ�Y'<K��Q�͇<�qNJ[����cc��آ�a���u��'�,P>��&\5�n�ᵡ.{����%]��l@3E�i0s��Ѿ��',jg �b-������{�$���C�D"{3{���e�p� �6	XI������{)`�V��;i���$Ԡ���'`�����0_~�֎�6pAؑ� ,kX���� /-��/$�gJ�ԋE�P"���01Rj���E,>�����x`*��������ζ�K,9a�	Pw`�欷�v z�j[�Uf�?�L�]�HX��՚3%�\ ,���7���ʸBe�"�i�+��b�O@4GP��ѣ���G�j՜ O#��*�#����PbrreNb����K͏�]a���X0#����F�slc�\´q^݌hmK����	�=�q�}��
wh"k����Ώ:���'���?�� ���T:�I�"Y �@3B76�Mٚ�y��A�Ľt S0��tB�Bۧʣ+ � ���\��5������ܟ��o�ץI� Z�����}J���O�!(��Z�H��IS�\���<�T�W��`hrX���ė�~�%�B�\~�,a�*u�~w�A>O�����\�j`9��dVJ�,|:��!;m�>W�>���A�O�@=��y��wwx� �"��'��K��Ŀ��ʰW�M��vo's�S����+K����������,��Yz7�����r��`�O+r�i��6v��Om%��^
C��8�m.���<���1>Ͽ�_m�UK�:�甊&8�!+>"�N��	�Q#��B�س�q�t�M���o�B�h���p��%O=��Q	��y.Ww4�1��V��W�l'R[��4�P��;߫�_�*��,�E}���9O�8G`��ꬴ��^���{ㅣ��d�X`iu�����2eC�����OU�ی��ړ�-�u���橰2�co����wjYP;U2��z5�%�o��]G.�ďu����Z\`x~u�J=o�}6�ڋ:~CS�Zi���9Eȝ�����Շ����j�D���!\�F�ϺEy1-���ؾ��]��5 �ܔ�{���O�K�� �$�����H1�%����uG��m��6�J��S�3��A/z���mbf�'m`��w%�?��`^�z�bv�&K�_O�3ޖ�t͓)��~WVi��(�Q�3�?���
�B"
Pv�mB���.��U-�l1H�>�@�R��J.�c	��d��whٱ����v�;���l�F��g"|}�$Y[���%��6Z�Ԭg�uD�
��F-��d<�c❛�V�7��j�I�D>T��B2Uf�!�Yr���/�����ff�T��]��Lŉx�Y���l�%L�pQ��;�i`�§v�$�ʆ���9/���nR���#s�y�d�;���୓�$��s���	ӡ`1�y�-�P����gq��;U$�|�OaEd�/���<�<_F��
����@�$FL)D	J�p���>DD�^���j3��3r�U�!a����]���a�.�!�%/�e���D�n"�"���	�G��[;qw<�J�ÿ�w-�����b���ɋ�]����դ%�E׽��.G^�
�1� %5u~��J@��l�^ם�&ch���A�U�ZUgH��ӫɬ��6�����}� �M��#�z���EEI����\ܱBk>\\5|V��vFi����}e5����#�nF~c�E������q�]d�����@;��v޵���08��Ԁ�ݭ�N#�nV�i��*�ݻ�9��`G�Ϝ�z1te��TJCF�c1�{���C/+�fλ:C���'����ޠ������T<N�\�J�.���(K�$�z4�)����z�tb#!�Cj8
�6G&�k�=��������0�9�,��w&'�������z��u"n,b�l�Ze@��:c�K���������<Q�~{u2�?��5%^g��A�!�&ܾV)�ڏߪ.�m�����m=�k �#j��$�=ֈ���=#��L�z��2]$h�/�-�J3ɯWʘQ����";Ӗ��>$oǖ�8C�������_F�VHy�P[�C�_�+�#)�fz�v�Ċ�uX��!�+��A\gq�| �0�Xi)a��0* ��#P��B0]��Ƴ���x��I���V�A�����O����&wMK��}�����ع�͟��"�N!���h�kG���9 	������n޼�5#�u|�#�d� NM�,U�&�&���5I���A
"�3�
��R4�!��*}o��R]�����q�'l���]�CW�2�ŤX9��t�iS{F�8�2�!R��ŉ�8{+2k��:2�^}��n`��c���a�nKTd�`1h�����q���iH�����9��Ny6��+c�]7x'}׻)\T����XҾZ��o�9�ȹIW�J��nc�^��>8~�2w���vɍ������h)c(�:={�W���C�DLA�0�0��9�0?��<2ͤJpm���D���z�c���)�˖�šԬ:�Z7�@ %�Ʀ�^�IZ�pZ��Av��y��_!����vV���W.$ ��x����cÀ�ל�`��e ����|�H����LŒR ��=��=�t��
ό6ϡ�h�F΢G"b�9��˿y��1��S�4.��q \�ĬB@�V�����N�?u��!@����D��-�+^���wE�����9*�fl�CG!��g}:����Ks�i2ߓǫ����h?��1�������$'g�	��7�o!֧�=)���Mx����8��"�}�g�3n7Ϋ�[����8��.I�v�2�5a%Z��z��(�7
�Z;��7�0�Dq������O���ͯ�v����/�/��X�3u��/4�:���>Po�$q�^�<�7�'�K1̢�؟��@X��4�&�>9/�a�U�Rl��5����hS�����V+����"$6���p9,��g1c�Kb�!(形#jL�
���\�ߞ��/�A)~Y���fU��j����tݍ$X�?�*&x �֎q��˒�<ZZ��e;���P_��h��}I{y���<fLVM�F�U{�)�N��=Xǘ����hoд���`��y3����ca@%��Ƞ��/��+�$;�����j|9 6_�&7���bg�?��7 �b���p��H�w9v�܅`�y�<���fD�����p��߇ԕ��*��$�N�g��=�Dc��6RI<��Wj��쌺�C��3#`2��2-���W����z�eY�	:g�-������h���c���ri;xO	��P��/��T��^�n,�@z�~���N@��s���3V���U�Ö�<*^Ĩ������U����(�m��W\���	�Y%) 6���8{Ak��0�7���di�gʅ�w4���4%/�X�A���B�|�?��R�ֻD5v��K.�z��P?=/�Y/8C6D���P"؄�	#ߋ��zRipm�2ܶɌ"�kE�TV_��㈕��>AG�׹<?��0ou�|]�\�ʒ���%^�&�Mx�wu�?	�ml�����Űz�t���r�v��0�uf7��'���@9�yB@Z��a�
?g�[�s1Md��*��'y[�e�>�V��q�:՛�l
�f���k%�@�e��*��"�%Y
��ܒ���Y��@WN�K�3%d�b=�W%7�IZQ"�l �gg|����s���!���4`��{��Ff�染�
[���>^J1�
G0[W����	���V#qj�R�\����Jel=��/��Y��  i���C��L|��}z����n���W�
��[��&�v�&��������BbbO�.��s�΅���N[�7���b�TP�}>0��r�/Y�s�	�MOx?�>�KԔS�J�1稰m�d8`1�~{�mA�n kn��!1̈�Uk����,cz�*L��s���yJ��G؎/g���m�u�{�P܉Z�TQTܴ���]�T}/K�i*�W�E�����N&�@SU �pI�Wl �g���`.���y����>ᨏ�q�	���}�<q�^��T������ȁ��X�[l�ɑ(r�)��01�T�lc4K*T��@-	�_N���$�R-mV�|M���b'=��{?�1e��JQCrf�*%!h��	�b��ݢG����V;��҉F�����ʬˎ0�"���%+4|�G$���.����
�����n��e����AɁ%���FEϲ��-m9����$('�)m���b{��ƶa��^���>���(]k���	!�?;P~����@7m���@�1��L9��Y��Ks���g�l�h$ �qm݊�ee<�2�����v���`:�z�WʸL� $�jA�\�-�7bz�XlyN�D�׳���W�Z�N�h���˧9.��-D~��Eߓ���%��c%�ˢ���G���û�b���'7 mN�;%g�U�hz��{O����ߒ�	�J�+�~;}�^�l�h����|���XӘ�[�j���^U��UHx aK��'0@��Q�g��]�%��ZQ5�z5	#8��L>>Ti�C�R�RvZP�ίG�W9�$���>8$�ґ��Hj��R�~F�e��`����|�+�������إ��� 3E`Mg����@��W:ƍ֕S��HC߸��rWtTE�4�B��4�H�����#�M�3�K� ,˫�M��8�$��	 ��D�}{	Bm�	���^E�k�~(n����x�4�
�fЁFs��ǧ\淎#�{=� R������HK��4������N��}W�������Z�Q�*3<�L˳Q?N�ѝ�;��I 8<V���\����������� �䫸SH��IQ0 5A>xQ���Qt�)u�uJ��˩���﨓NU�y����P��\g%+���F�y��})�2Җ�d�Wa܋o)z�"bP��aU��Ҍ�mj�5������'�G��x��-�ȡmf� [�#F�WX��A4f��!�����&�)/��^gy��j;��l�(��<��M��A��,�`�2�Y�U[8����D|�ǤC�F�/�Gtܪ˴1����3�'s�nQ]ja��I0��A�_�N�r����2��[�SOE���C�ٔ�+�$�#���Dt���_]���IBh$RB͟t�KZ;��`���|�{��+d�_0�َI�z,ۓWe\[�|h�+��RG�bn5��;؝��h%�7�սP�n�Nۿ��s�UP�B	<NZ���IP���s�^��H.�f�8�dL�z���8��a.*a��Ew�.��k��p���|D���	�0㵽N�kN��S�2j�=���3�s�E�n��:�"�C��(�&���jq},s����[b����l B��RKW�Lj]���5�Z��z�̭��6�{��dq�#"d3_�X|@<&��ski�oK�+��A�e#A@,#�U)�I���y�"���ê�� ��Mp�J���A�N��RV��n�L)���\���?���c�����0��/<{c+'U��KuXe�7��`������(�HV�S���	���� ���j ��ynC`��`f�����)hO�w�� �-|F�ޖ��N�����̴fQ�1�����8�堦e�s/=�G*]y�멨]?}b�n��0˹Z�qwwՈI!�k��$���fK����6�ܚ��qUkl�꙳�ѕ�P��.�� dZ��Ұ��z񓇎����� ��,g����̿��Tb��=�e;7 7��k3��$#N�]aV&0��p]�^�j�硴`��Q�5�9�H8��y�a�I�S����A?GLF�>u�^���)�l�`���� �q`G�q��)�6�	/A����S��S;���,���������ڵR����/���{��̓ ����خ�"L+7�{�řR� bp��aE퉩��d�d5dv�s��Q�6�8��-�D���>c��O��MtX��.ؗEu�� �}�-�&(h��q�1䴨�j��B�Ɇ�����@��BD���^�_��,'X���.8��/�&N;O�7�IA������&�&oV��%�9�{�*�)Mt-:�Z�3GN�n��=4Hv/�p,��(���^�-ے׵�5=�߿5��"3�՝�/J:@��ʇ��=�7�+|S5j�5/�JtD�U��.4�<�R�F������d36 h{�H	0�Ϭ��\<�bS�蠎��� ˚�L~��wm�4X�WtΝ� 1�௜{t*kk�<�,M;�W�n }Xj&ύ)~��I�ܕ���e`MP�x{��� �ԕ�Ko�z��zZ�{p���A�6G�/1O���7����n^��@3{�E;q����F��Y*�E
"�+�B��wW.���Cz/i����G�Xbm���p2���!��M��wW t`۬��0�_�w�ԇ�7�#w�b��w�,�AD���V�'��b�J����w��[M��x,t�`��}�+���8�$�qׯ��4I��:�����1H�w��q����(��8l�!8)���ex���D�1��L,�Z�C���?0s. �5Ώ��~n��A^�B���!x-4]�j*ں�Vn�f��vr�5|��:I)����6�4Q���M��O�i�v�S�A͛~����ˁ�/ow=J�������_�rǀ��70q��@���_}FPA�1�B�������F�b^#�H'����C�Kn����j�Ζ/������)���@��ȧ��\�1��Sr����f�ZX+8�z<���Bt)�������V�g[v�f���%NҼ�I�f����?�0��uCH�#����B�U2��'ֿ{r敪���1F��ŋ�qRd��� ��` ĵ�uk�U6k@͈��Xy�D/�O�F5���&}5�7LCv1�L�1�^�޴4>`ϋIje��.�KVq�^i�����4�-����8�������h ��(���A�۝�b�r�0��Mw!&x��-��]N1��dia��j�]G2,RN�d��)ܴBF�`�����΀�г���]��;a���u9$z\R�?�F�R�xpq���c���sT4W����Q�1�F���I�2~�v�)��������"3��z'�����av��/;IF��T%,�&V����72�̖�	ޣ�����QmC�P�Ftݡ�-[yEŅseb���P!G��)pV,-�0�ߚ���C�l�o 뤰�-���#C+H��`l/�����.Ɋ��f��K5��.�2�b����h1Z�v~i.���^��|w�N�uT����V��&����b|�)����+[��q��+�ݕ*�	O�@��:��
����Dݜ���>3������s$N�bH��͚�:�u�׌�����/��>���TFT	��`�CtڡP�
A�$��L��H�Įr�IR�w1�L�mg�=k�n�(!��^�z�eo��ٮ3o���I�U�6͋(<+b�vi��X 	���,�o�T������;D�8�xm1���*�'EOV��&UVoի�ܠ,�!,'�߱�1�qOqWP�1��mF�'�=?����	raP5=�1��w�����a@���J2^#�V����Vv��vL	�浖\?Q���+�o�VO�*�JHG������6_�1"��V�Sfq[�.C$ڲהZ�Β!b�����\��l��"i`����&����X��Ksǡa!B���~�-pu��&��M5^�UE�V��P��ťc����t]�	�2�Ɣ�� ߏ���r�H!���[.~2�ط�vl�ܸ#�#x��4�<e�Ӥu!�Z��~h�`���  �Ca'@S,��B�$',;ּ|��jC���䀑Ĉ�����:��j��"^w=	}��X�G�GdK�HxR���l"�".����qy�̷? Eh��H���-����1C�~r���Y�;e�C��xyq%��d���Ε���P�,��
�����{���i@�$i�u3��B��(>}����j$R"�� �,�(��[ �E�����4�6�X�I��6`���%ܯ�q���H�K�����y}#窏'�l^�a�w�!5�u���	��������b��(�5fb ����/(ER;�*��&�v�GBJ�w ^N�G�-=��oD�z�]غ����:n��˲����eѠ֞P�ه�2� %*61����R0LI�:]P�h���v�c
d�Z=L���6�5����ޛ��kY:��Eۗ��K����X����H�L4`&��J.0붖����8��9)�G}-eÂ��2[^��M;�b/����F�ұ��6%6m�{���}��ݖ��� ��!�[p�{�.�t=��#_���?��`9��'w~�ǃ2�?3�U��2a]R��q�v�J
�����'��_W��m���a�G��0�$U�=���h��<�6���`ݘx���q�A`��?��f���n�
TE����'�GZ7;�G����5��{a��s��!���bJ�z$2����;)�S��l��wc.0s��1�խ�ΌB@���%8�nƿ�˾��!;�. D����cc�p�f�9-N��ĳb�}��uhp��X%	(�u�����"G� J �� �tZN�kpM���I�A?T�K�*�!�������Ur��t8���n���
Q�u�5�o�)&&��G3�Aj�d��P�Ӌ��p�i]��,�̳��_��U ƍ�e[*��+�#t+�)+��������it������w��%�Eސ�>{���X�x{��ҶNSM)��|���<�(H���a^j�Z������P����
AIgw*[��I3S%Z�=�ci�Vw���|�&���M9���I�o{�fCDN�%I���\t���`�Z����S�_ �^���R�v��|Å����Q�]4���tE0HW��6�`^�V;�i C�s*���s&@�?��'�V�+=��MA�%����A��l�!M��u��(d?�D�$s���N��h�b� 0���|rL�\3�=)�e��=�;(d)���=L�xM"���Nڢ��)���a�@�g n�q�u��y�Ƹ�j;c�$9���p��|;�+$��@���4Q��>�������O��w��O������]��U�J5���7�޺!�Qgty �����hڻ$F�(o�"W<f�5ޭ�`�+g����e������͏Y��(C���'�x����'�LYP�B5'�ٚ���
�v�F�aӌ	.$�ohW��B�9l����i��OGv�	��sd���S�.Y%��>�q��@�2R*��C�錺c���N�L�Qx�t�TjQ-D�R0Z�q�+'�c�З�S�י�4��q 1J#?�*Nwt�����
v�!.n�pӠg�-�AW.2^��N�=�eieȜ~��FX�e+*7x
>�=o��SKP�����.�,my�t�KV7�d��U�('�G>���Z1	@����[�@�����rM?|�q��pTn� 0�p۲7p�>XKF�|�#����A���Γ��Ij����K}��z�o�����Qn]͏S�n�h� � $�������Y\1�(H��Õ�v�\��B8���j/p���)�hM��,<Є΀�@T�2E2�چIh�丄�ѳ��[�~ҁzzb�H�$`
Q�̻��n�SC6̌L`5�b�B���J+�_�_[VM��)x�l�V݌D��kޅUEDA{x�1�@=>�}�kX�a(?��� �A�����o�w���ǌ!�[�Tޑ�"���Bom�b�e��n�]B�B��5(�Ӽ�l�!�y�&���o1%ն���(�l���z����؆ �%�+�N��]'�/�ڕ�#�5~r��a��{����B��}�'{�������n��^ �١��{�s�QG��z9�K�< ϼ�B9�����ՁG����I���T~������8JqU�,�Ť�Iz&Sc���n�@ϣ��;O閃b��|i#����-%��8�y[�ܑ�<�=�?��N��}Sg�AӨpH1�f۱���S��󻣮�m����S��ib�Et�~���*.����Zņ=�߶�h��1N�.z��i6j�t�X��
��e��
+�p�6��B�u��%˂y-0'YS�8gv�Y��T���jO'�}�
�Jd�ݎL���݂��IS���~EC��s�Bgz���
Ѓs��I�A�t���Z����{18�*U}�^{R������m�9�r�O��b����͛j;VX�A8��|����d-�I|c�����9�L��r��da��������xn�	C�C�F�f��1��dOA!�7��s���-�E9�/�!Xc������Rs���EC���}jν�`����9��]52n�i=`Ҫ���>��u�GU��N��~��d|�U_O2q�j�Sm�|t����$��F؋�T��7��plt�M{��{��Zgl��Ϩ_E��k͔2�F:���:����E�9�P��a[�"+�L0���1�0�-���QabS"�'�K��cn$sĿ�g*��mt�F{S�xs=8��֭�[�*���~�8�R|��k8�m����
cMO8�Q����w� i�]�a
����ە���Q�Dd?���^�S���	y+C�g���<p�7z��;��*�%�B|��fL`m^Xg�39�☁�o��	�֮ �o��Ph(�>]3�c��X4=^��$�=M�{m�(����� �\}�H c��$���2YN�콤c����h�q8S��ͱcyFA�}�,V����h.!�]Ih:gpc�bueCC(����>|I\@�|�Õ���4J���rM�o%7����pm�Rډ\ɡ��>�雿B�Ԉ0�`�"tf߽}��w���2T��~dFV��D��/���pZ���N���K��� .�A\Y]ty��X�-�o؊�$3y�a;�>b�)��2د=sz�V�Sb��8E~����n�̳� ��8";d����"b�G SC������2�0c<�����]��s%(;�g�8��({}�a�Щ�jJ�=����"x-nG�ᩙ��{�׵����'Vs��ߙ�?#�-���L�ȁL$������`������T�z��΋G0s��fov3l:�&r�0h��+�{�����[r�^+��O֖�����D:ZU�f�zz�����~Qo����������H?N���5��t,��0"�	�琧m�o�F���)^[zY��!"���B����;WA�˔�c����U�. ���J�W<���APvy��A��{_3�+��c�����4C;63��J6{�ˋ�s1��9�
zb������R�ȉc��=(���[
$�%�f.�o*��5���]!sy>=�l�V|Ⱦ�OA�G'���`�щ5�k�y�|z.A�P�w���\�= r�5;��D39s\�O���Ύ����(�/����
���x��!��%�S�;.s�6zx�wx�ʯ%�V�	�_�rV��lQ�4�d��U���'Pļ�^)��Y�}s���ip\+�Pȩ������
K�ZŃ��l������vP�}0G{��@<��(8b��jUp,��BgF#�����]���,�l:2��Ж�Wj�s�/_:��z�i�VT/��e�\Rg�F�CH�O�U�Aw����E���1�Q:��(菑��Qa ��bZ�ܛ�d5s��t�A����d�	���Ю��#���atj�5��#�>9�H�dX/zM^���O�w�v(q�Sy7��jP]��fJ�����w%�w��Du�7`���5��\�8YǠ���� ��)*G(���"ATT�=���+�M��<v`a��>��r-�᝖iR�m��?�%�o�Gߛ״HM��(���X���5��C=-��+�b	A�H[��2eS#�t	�Aj[�D�/b?�(���W����ԍ�,Ȥ�^���龴�*A������dZ��K)�_{��dU���".�^���w���� �d��k�pƮn����%єޖ;9�J�i��PA��I������)�?W<O��'I�0�Zt�[�i�|τ��Lx�ṋ2�D�,lD��z&�&.�"�ſCg����b4Cd�[��X	�s�A� e�����[
Qv�*���_kȟR�C�T�z���2C`X$��-�40lR ����,_a(�*��w�~;;?ӡi*���5���K���aI�:��gD#R�,����;
�U�ػn�ݒ������������
�=犖�POnV����S&����M�fb�8;*/D��[��������s���н\17�N��3���	��BS�~�Vö$x����Qh�ƭ:b*l�=7��k�ƌ�MN�!�?zc�hZ)��/`Z�HQ�Un��2'�����Ʀ��c��i�!'iW<6�K��]���Ww�����B?�0��v�.�k�2W���3�|��؎��E�&��*u���%l<f�dy��հ�^D �:q�Ǐ��W��c��`����u�d
���NF��_IV��gL@X��K�]3�5�1��g=������F��R��	72���XYѓ�q�y��'��WP1��cn�%x^��%��ϧ�/{����_e�T�X�w4v�t���,�g�3���>0���Q�o>���8-��q�B�'���կpLU�a<G�<kN�#�Ԉ9R�̶�[�/���˭���)ث%&����Rې�q[�ۨ��:K}��a!�i\(ǽ�gW��VQ���:?�-v�J〺�_����a���f �"O������ʀ@hkŅ-�A����bM��5N�2e[��O�W�$
���j�< �����5Cf�qm�S����ra���1�8Y��{�i�����J��<�S؜��Ne�1;bbO
s��ڮZ?��Ԁdf���i�,��b�,xb��1�^�M����<�d�Z1LD�[�2^K%�����@�uU���ߊEo� M�?ܠ\���^`ܷM��BNwk����7s�9'o}��*��l�Ze<០���c�.�ʮ^�F?�ː���}m(�����M]��iQ�pOQ�s�Q��/�{�R�1��4������z-6��wRP��cz�D�:����B�bʼ#�j���� -L�Y:+�h^�3���d�܉.�I�Rah�Q'1)���9Z�1~��j�pߐm�+a��Sq�1����?��9��=�d�X�7��q>�x0}F���L�DiQu���;�/��%�Cd�s�5a�Q�X�����G� I� NO@ ��뉉�Ԩ�7I����7qF�O H�����/n��#6�	�G��T�+n�:F�]/2iã[`�s����rPڷƭ2�)�;&M��������[K�:*�K^�����k�ߥ۶�����XC3�"��[�L1�] [M;�� ,��g�L����(���e="�/���!�4w$y�D�/eħ�NJ�MR;����(��!.xE�C�`�e�F��S���jU�L8Ue��<A�7�i�_�_^94AB�G,�r���A˦�V��)�.�B^�~`H�5�DAG,1h�j��ѨC���[j[��[���ks *sh�>!=%Hg5!^	0.61�ƆB1m�v0�lIL2�.�\���3�U�6o�n"����~�8E��)����"�
\�O��C챂����1�dy������[��+6NX!�3����Ʃ�,(�1��*u8�xr�*����*~�)gqVa�c!ؑ�Qo0���BX�P���54�T�V�
)`�=qw��t-���`D�<�K%,Sn��Dh�i�-���g���*o�H8' ��>X��j#�:7�F�"�����m����*c��$S鴚�l�ff�Ϫ���=X�u����|@ )��%Ų��"^�:��sh�ENy\����Z<��Υ���P��Y��9h�R
�������$Wxus�?�ń�7Ų�R.�\��Y����c�c�p���E߫�h=CM�>e(Q���1��)�ұ1�"UF��D��l�B����C�P���F52���1�j������S�Hq��8s]�Q2��p%Y����.7a�@z� R
c�W�gs���s��Y�]�p-w��ytp��V��9�c/�SlY�`Z��% m����Gӊ�	h����"mR�(�cO�}�Ȕ�r��Q�R��AxlZ��(r^��=�,��������U$��%�\`���k{ ���iA<u��04���$*�(������Ť]kA���9�6c�@�k�$�Oan��	k�y���^��=Hx��%$$`�}p���E���:�v��\D�|*��WL����R�bɼ,����+{f,��ˈQ��pGa�O���6:�Z�����c�e"�>�v��2��v�aYyH�68jf��y�U9�����u�_�������tYs&�h��W��L��Xza������i��j��[S	KtT͌���/|o	��,d�n��h&���l��M�"�
Ք��]0�0
xq���W\r��z_���縗"��|�M������kO!��9vc���[ �t��#>8^���"�}����L���Ͱ4�Q�`�X�F�rAg]ϱ�uD���El��9c����Ij���*i�z���������aa�A����<�z����Qt�q,�Բ�#3w�F��'������*{�譕81|��x����2�nX@���~ᐔ4RXFN`�y��[���T��; ��Vcuh�/L4�J���S��D	7i����	N<�7p�rս�g�&�Ԓ>
~6�R���:.�xsD�LmMǴ?|�����������Q�OAcF����r�=ԇ�|��K�ϊ�s)$��h�t�-\bY�>�g�*��Q.4X��&�)� 
z�b,�s{{��.��i�!7��;G%̀�����l�=��w����e�[(�{C�wTiʞ���:nfݺ�-��\�x�srcw�����n��_�cF�2�T�����Ņ�B��3�S��i���Q��]��If��L�j]���+6.4���?��BzoF?�ʧ~�66��B&�8�r���m9�֬/yƉAz��؊�o`t�/^Q��s���-V=۽�������Z�6��#oY�I��ʣl�F}�U�2�{��#��w����# ���x�>rm�Y�w/O�v� %��ji��_,�a�<��M��]3z�ޚ"���o+wzӷ�X��l�[=c �\rqW��'�#�~r=������%�"�M��Ok:�������IV���{��(��eH�b�ۯdr4���Y�h��߼2�/��)p��x��6Πe�
p��T͌��H�.���+ �����iRE^�=�����|��#@��g*��գ��k9�7Ǭ[c+�q�l�~�W{��5Q�}����E�����l�6�9כx�6\!��]f����놶NQK��&��x,%�h��)�N��M�,,=uY��tsk�U���RK+6� 4]G(�͙R8�Qv��lB�˟Ck�c{y;�5�nd}���u-T�qY8pLlq�A�uASP�/��=��;�h���#�IQ6��2��ln���ql��֣�ъBq��p@��֖R[���S�7פ����:�{���No�w�����ゼ�T̩�|q)�=�^Y�o��C��IH2"fes�GJ�H���Dɚ
nd9i��C�!fT�0�v�v p8*C��z��m��Q� %��ZA�򤝪.�6tZ[�����
GS�W�˰��!��p[[��=�\��08q�Gl]�<G��G�1-��>߰�\������"�rĜTP �W�8��H?�2f ��ܧ��5����
2h��J���u3*�.�/Q��~'���@��V�޶����݃:�R�����0y)S; ���g �Y���ϭ���k�K��9$4�'�ؔ��z�0?�+�Z��ђ��#ҋ�]�D7�q�3@�J�=�"ε��,{צ����O�+�|��C�>�Ť_`�8�,v�ǵ^��l׋t�{$��������ݜz9~q�!�ɿĆ�'4y�V3���J�!�\J����G۾_��{V��>�]����~�t�jry�2�x5�B��$�1-|2n��AK#SLL�S�uxk��MgH����+�J?�"h+�>u�?����΄�������<��$3I���!�2yQ�R��K���0M �pxB)�Z^��8�=��x�G�>�hO.�g^3e��+����O��:)z}�]]So�M��*c�DY�r���.^G|e�̆�$�"�
(�S|��-��!Z�j2S� ��@�{�pǁ���u,��)���o�As��%�]+�`n�ݾ�����'��I����#���!��a�^T������UB{���,��>�9&��G�{W_eZN�w��G���*@�e�߾G�����_�E(Hґ��˂{N��p�̝vi2\7��EiX��h@�9�%���{t�\����$�wy��ǃυ�1��#���\��)�d\7�ߏq�n8��xQ����&���s{?",ޝ��k4��6�EdG��$��ŭ�Z��=���;��U5�9��O$Yg-w�|�1���@	{�����g�T��Yi3vxby[~��U�z]H��O��7b�$.�/���I�pV|:`Z���,����1������L��� ��d'�)BR�lB]��cP���i�^���b�G0���:пa���J%h�،˄����i���e�`PNe�A4톟Ϻ"�`r�B~���<N~r��:2�8�V���%$x~7��[��Tء �����Y���	��=��̖�[o�v�� ]��ۚC52�o�6ȯ�<�~�'�5���g�]�-�Eo�7�c{�'�7l�<�N�z��]_֜�7�[5�F�\ �u����	?p�g��G�.N��N�So��̖����oc���}a�N	�9���Jp�)uY����S�9��@���>E'�5y*�U'OI�1��7���E`3.��K��;o�������]U���YC���-=6���������4Vs��y~�u����������8�{n�u2�x��&<p��i�8ZK��8�+�;�Q���t�F��mPݣ	MV�(>������`z=(n�ut����A�\����1u18�ct�,�
�29~�q�!��c����;���Mt��	�85
$kB���kmR��2U�[��п�b�/��.?�HV���ک�s�Ä{�"������>X���%��UV�I9Mo��ڵ���X����+���=���dq�	6�0Z�h֙ۊf.\�x5xS��E>�c�hp�ԕc:1�(z�>��&k�jw�#�&�`a��S��D�Ge�K. o�goH�<�(��J�Ҁ\��ә��-�bR�)p��
��̈	��4*���:F_1�����|��:[���,~�W��[IT�?�q�tK:g���+���ڮ�����Ve`��=�HF�;��L֑����h�� ����+nb�zp�^O��Ԋ�����{���z�CT?QAtLMd�I��tΓ�r�ß�^J���SΤϣ���z]iz!Z�"�Q&��NT/݌���!Y^$�
�Xp��ƌ�t��3v�<�6���޴�BAW,�m%֑�M�A0Y_2�7@5d� b��nҡ�
�=���Ze+ɣv��g@M��N�A��`��J>)DH"�B^��Re�R� 96��I�坈Rq�v�b��,���,�/�]�UCޞ����z#"�4�,u�-N����7���G�ޑ����VS�T�?��x$;�>��a$��D�l(��sQpD�2�~�Fs$�j��3Z�f*M����E��M/u�P�ح؇.�ٮ�_���X�Ђ&�?d���A>)������T6��}�r߸h�Y�8�=�����		Q�h��
��1�jN��[����L�����I��pG�42d�/ֲ�D#Ӊ�R��C�#H�H�]�'�Ā�Ծ��^g�$;�W*����l��ւ�glN��X��/�m=�Jr�m~��Γ7������
�[�ɖ���:��A*nB2����o�'��@`�;77+�����^�}hT��]��u��P�$!�,�N�DX�-qW� &���wR���sB Ս�P�</M$���H�yt�Ɥ�mBS.ہ�-\	*�a-�5�,��R��'�߿k�7�C��:I��㾶�����Y'z޵��C�˸m��J��S��$�rɯJ�(.᧏KDSp�}�p�����J"0�Eu�W3��\�K�tc�+�kLɡ�O�뻭�F.�vr�Mo���<���<�'`��{��H@�޼�V?��9R�6����5�D�4^f� ��x\,W(u��b[&�� ���]��^��	�]r�<��<`Fa����O?��7�=[gt��Ǧ_l�WF�J��М���|�MA�<��9���I����<g�m��pU�r~T�-$���[��[�8.�e(���W.�z�
#8�ae5�R] ����:!��`Wd�ϋ��ǧ�Ei��%��H��Jׯ�o����6v[ٙ�uH6�!WaY�r~6���B��K8��}�JU3%�
��G�����˺T�:N�3t�=#�}�
��Q�qZp��D8Dt!OliBD��S�\W�C�@��)����" .T��:���e#��v�{��-��9�4# �8?�`״aL'�5��^�a��j-�)�����S\>iQ3���7��ށ�m�.)���tH}X��ӥ�U����v�]��K ����{�t�;\�����Ȗ,�u��S�@=�^U�{����8��OCљ�"�ςX��_VbX^�=ޯ��	�(�쩩k\7��,ጛ�s���
v�q�]�>�?�|�7�������0�ƈ��C��EU���kҳ����N�YK�Η��`�ݒo?�7�w�އɕ�]T�z&<R_d�s�/��vtL&���8��_�$���W�!�R�<�	�)=H�%T�X���F}Xc�ÆA�	�[n<�S�t _�A{_�3�[�o.ҭ,��Ms�������BW��9�w��
'ʚʺ]�u�$�����W�!lF�BRT��.�n.��w����ù�G,AU��P<1�>�i�K��z�7D�ȧn�Rf��=+N�/nV}K��B�1�*�Ϩ�Fg�^�����g����\�X���N��S��mL�����\������sBh���BZ�Z�D3 Y"h�w��&#��kyT�]���v�l�������O!&�R�i,��Y�i�p���v��b|�\e�}��=���4��%��M, i�^l���#��UQ%�"�J�&$>.��-;�.�+D�/
bÿ� #3����z��!]�r�������+��{R�Ȑ��(�j�O������.�����V�X�o�3v��ᩛ�7��Z�;}+�8�p��5��u����HD�xW�bї|��ƈZ�E6�R�U#�g�ҋ�E�e�>���,��1�tL� �h���	�<6�1OK���|�������y�����S�Ȗ���!bH�oڪ5�U�����S�5�iҜ�^}
jN����tڽe��p�`�����-�;��xpI�O����E�:�?Y)ex��R���m����9{�k-o�&n+�ƞ����2߻���
ٍmB�q�߶?�.��LDb��NQ���`r������!�f�KdB�0��r`فy��L"vu�T0��TIأb�	��<͌U�}G^�M!�س��=�R�����E3�iP�|>\�ټ3����Q�	�t��j)�n��6��P,��7��b�D_�a�s�5��ʜ �6*��m\��%�ܷQI����k�n��A��c�C�!^?nm�۲0�ay���$6�Q��GB&j��'<މ0 ��.��9в�g�?3.fWòl7֑�E�2jJr��r&,<��h�ɼ52Eؤ_�����П���n�`��&�W�p�S�̀F��r���0��۩�t"p�"~f"�r{�Ԗۛ���i��A�f�:�� ���jvZؓ�Į`�n�DD�N�������h.9Nq�3����@�1��թ�D`<}��e�>�P;���sy*S=%M+����������rB���ٳ�M��'h������?H<§�Z�Hj�ni��o�=
�Zx��!��v��cl{~�>(U+Ô�-���|�N�O�{2@��>�4q��U����r��(�/Jw��>L	'���%?^�O��ݔil˞��v��gi���s�NP�;mv5�w�S����_�5�lxP��\ִ�S��MԦ��'�"�s�*B���j�:t�߰���{�d	�������t���sG�D�b� ����ºo��Mu 0ެ>���I'Gޱy��%6�����t�5Szg�wh#��v)ԓf�#�����k�T��x��8�F�3�O��R�B�뉐�`�٤+O� q�1�h���D?	46#��$j�,#��� �׶�q�`�����}fE�3�EeK.|p���@v[,Y�븟���K����p1|m_[RAٓ���������{?o@������_~r�]g�IJ���=&'��چ���-�wjô|_��hN���T[
o�[��o�}2�=(��QA7C���L��+�N6�m�V=�
Q�Au���v�`}z<��i�V*�K�-���Fے8�N#�ن�R�GM4s�#ϭ���)�_��?2u�8�a��"�#�I8����#н4F��K��5��`�E9|���|{�׸k�y_�zX��!� �DWb�<��a��V��zL�/���s֟��ޭ�felO�8�����G���쿴w��sD%�^ ����[�:K��Pl�0�2bn�L��)Kw���́[�M���<������H����XMu�$�Lx-Z.��jf�pE�xC5�c���E�#�Iu=����M{l�n{W)W�}V�R�M�߿xLJ�ld�W�P(�lOު.<i�/\f��7�A"����>�4$c����_���,���#7v�{���5�k]��T|��0��*#5Vu���ڢ�YY2�	]�"��uܒ=�;M%��d�Tx݊n{H��M�X�t��M�A�zH��-Wd��.��H�
�_U�T	��|�B�2cC 5��''5Ӛ�_�!N-�] ��:���]�Kn�P7�N�Tl ��R�.g���ІU�Ց ��ckp8��g�97DvzF;��ܾ��KV�rހ84���d|N��'8��8;��	%��bD���"��4��P�Ό�x&��+ސ��ob$#�Aed]D��s�w�zN$mM,�E;��T�l`M6n�:�'��kW�����C��~��_性�ʚZ���c��Yj�K�U�#(�%�2��>�`+1>����l� �,2g�mn4*��Ā|n�0q�0fpG��B��z��c,�p&'Q���qW����0�&�GIooE��h����H�?=j�J����W�J�i�A�8��\���X[A� �k��Gl!�R�CqéW��@�3�%�]T��3u2Nf�2a���>ߚ8�!��AlOd��?��@K��������{<�"K��P�5���2�yx7�	�T@~���x�	OҜ�7����ަ�)pi����V�������nB��e+��3��-^��N�	��`��7M .�|7m���:A�q�������7��
�F��`TL�D��ک�H�k�MEx�G?�'Ĝ��R�K�+/��w�{��/���90�a1�w�`r�%;��bU�~]Br��ɢM	�Zo��h=-��nN���%�s��`k{���ȹ�c�f<���*��6&ޒ%����R�K�Ӣ���ym��R:��X��g�p�F�^|ɝ_�!|\Z��{u�q�;2Q��VY��yB�Z��4�F�/|���}IY����vķ	��z"޲��^\�/�x�̓CD��)�#���i�&��G���q^=E�Fۊ��R��it�Hw�8����͗T.0�fI�����dr5!7xxW�9��5���fe��8���h�Qʣ4@U�����P�1l�� W�*��0��+���͉����8:�ZX��mr���%��פ��<�JA\��Q�l��;�Xk��m���V���`�5�2R��Te8F�j��(��P�y��(p�$̾�?D�����M��i�^Tph6P�&���"�(T���o��P���]_+-!���V�t� �ӷdH�����y�k���Q��A�\�UKxs�ԴiS=�)
�=�(R��hb�j����y�T-d-�Z>4m Ê��z��J���5�=��E���+D��:������v��u��eR@X�D���ֿӯ]�ŞAY?��<�F��*�1z>�����)� JJ�x�&�|�1�ظ�?`�$�j��??�m�Ĉqk�$�I���H�	[c�sT��9W=����W#�0"���Ģ�:���S��m��A�+��F��{�7j���AsbP�H~��Z\�,Q@�ܼA���n��*�A����w���������Qr�Ϊ����Љ��(�O����za�:��~�E^����t�z3�L�>@nqDNI̔�<7���e�	s8S�k�;��/�P?��&�2���`	_W����P)&q{ɓ֘��xSob	]`B�������X�0��.�G}��5.ҹ�q�:��c�	�S��M2c��q�\)Mbؚ� � _�A,Д�[��/�a5@�4�?ton�!�W�H����Q�DL�K��/	��%�����;�&}�~L��]ˇ@c\��'�Q�a����w��5p�������B��A��=�lAˁ((��K���BȄ��dL"V푏XPxWƬ���
�vo-V�NT�L����o�tk��bO6��n�R�1�C3�BkO������Nkr�����]������z�^L_�7y'c�9�����+p��8�_[ry����H����f@Um�<s�K&����@7��������
�[�)Y=a�ɚ?d U���3h˂U$���|�3m=t "���'9�w ?����+c�({�y��jܢ���ţ	s\�����R�#QC�+�7�l����K5��v�L��·˽ذ$_S(3l�ab�u��ik��y?�1��d)�^�!I���is\`V�{r&��9�vq�X�R��c2F~m��!�ZUpi%���i��!IZ�6��#� ~�D�u��ph�k�X!Œ�����<p�h��5�:�Ċ���)���I��\=�偣���[���\1T@�K<ϻ����b����dU���AW-c�)	�D��]������Nn0��IM/��!��[���8��3����@� �h_놇t�w�un�'�r&��]ч��W�L���Sy����m;2�f�b�t��	]�b�Q�a& e�Ϲ$��A�MdӮ;궫W]��-}�0B)L+n."I�u"�	d����q�����!4qvV'��m e�5n{P���'��A-\jI�4j��0�����Ӊ�l�T�>����r�
��9�3�����J\^��1)�@0e4s�,*�[)��{H�P�i����#c��T�ׁ��y 7M�+�BR��h�dc� �9��	�s����;������r�����'���׺	������D�|����<������b4N운�ۋz�����FQRo�k<�}��$sP���	~��S	1T#���z�a�O������ҹ�l���vv���`P�[�?��ɞ�)$!ڧ-LU({h����;k�4��%�i����v���%C���Ex`�%^i�5��1ann��do�˱L2N�	�5ꋞw�͈pD�v�2ZV��f�\6��%�7V}��)�
?������6�k������?O-�)��.֋A��Å1Ce�A=��	&nY&c�7�O[+�;���;5r8x*d�o��k��N��U
����߾6-."���n��ҭOr�k��c��nQX:?V�I��D�Q)Lt�4�˶��J,��0_'=_Y�Ą��������D��R�N�+ ���I ��9�� h�_�D�.C�K��hE{����B�>F&�,k�u^���>��ץ{�p��l��vk�
��G����&�ŅP�E�ճ�}壀��i甏$�%H_Ϭt=���-7��2�MM���)术 ������os6��}�\����[���;�?�e��kE�ƥ�e�TM�7B�yդ�s��9���g9����	�97*s����Uۖ��@��,�x���q@o64d;y)���^��b6z�m�`r�cg��38��Q= У�;�M�j��d� ���c"�Q%��f�g��_�!M����'D��������˧�?�5wf��G����Y:�����)~	T�;!��mkB_��.��x�o�sE�.�Æ�:B���-��	k�~>3��RH��f���5��"8�/�祷Sb���j�~��%J<Sm�vLu��VUi��چ��2S|�y��ا����^oU�`~�g�E�+Co���!.$E��_(�Js��HM�pN[a��Er���j��O���o��Ph����/�@Nq�W=�OD� ����R�nI�N������,��g1#���b@�v!+=��>���h��j1ȋɏ�_�f`g��!`���6s<[���]R���?���6��-�l�"%^� ��\-۫��F��������=LLuCu��]��_�����j��o�o��V{-���<�A�ì��I�	A�DB0	�䴲Q�����x�9kL��ۊZz���O]����^��83K��V`�?��q�9�jಟ/R��O/>��!$��
�vZ$��	?�N�+�[��5#f�v�շ��yI��C�9�`���3ʄژg�TxW���&0�%���+P��r�R���t�E�sY�(󆏨K,�v�[hR�(��1����t�b�@O(���m���?ٽh��|4ѹ��� �R�b!V�k���*���u&����a��E8w;X���u�#�䰢O���$�O/�ߵs�cv������E�PC� ����(.��9 ���ˎ�Z �m�o���{�$�Tg�qa�({<��1G�/��x�	EV�:��B:���ш�8�iVGؚє�O��73�^�kl$8�	V�� q�:	5.=5z�A'}z��,�j���}��D����J�4�-V��ss�j�̽pGW2"p����A�+�ɣ;&g<�Tܷ+��"�'4��8?��ޚSi�oy~��K!�1�t��Y��+1-�[{�|���j�8�gy��B�=ЀL2�MS������_�k���=)�q�$�;��2p�-�A|���I��q�&�;�`��V�eX���Ѹ%�3���FL^eɫ�kf��bI��Xԇ�+��C����

b�@snb�ٯd�!%q0Zm��D�䑋��fL/_D;}s�ãBʓh6z���G%x� �S"�}�f2wb�<�}ϡ�k�l�e���Rq۬28lb*��PZ��1���l�c�a�]����φV��Q�,v���@��h�:��5�'�*��A�����4�ېz���aZ눏������Y%�hg�����J�Z�y������7[Pƙ%�уM��A ���~ ���S����)Q�}�l�}L�7����PDWK�j��Y�G��tO�L��4�_"�eǅ$mw�#�r$�,�h��7'�~��2�<�C�nx��	� g	 �؅i]�/w�j(>n���$�8R��1��I{ښ�#U�����`��CCnB� !�l66wk@V�� ��T���L�T��ĵ�=���m�@�Y�
6��n�^�p��������� �f�����d!�l.X�n�t�����z�!*�� 6A�J��ǟVM��_[*�o����j��5��]�4<UJ��38	���m�<0��a4������Ъ�`�>��.�&A�9=G%>����U��x߾�g�� 6�2��i��F������+~o��7$ڭ���^�E�,�ʒ��1�2z�?����� {�|�G)�:p�?���E���}6H"��/_��
_�㸞�)}�l�([WV�s� �/�d5Z�9��`V)�ǋ'��|���n����͑%�jf���UVss��њ����Ɗd�ݗ:r�خ`K��X�
/��B������oD��fy�1�Պ8��C2�7���U!��K �L��l��s�o�H_ T)����yɐ���v��j��O�y�+UD��_�2K�a���g|�{���	�ɢ�W�QHu$c����<
	h�b*�`輼�(4$q�"�
僁��fr�m,Q_vJ:���}!	�����߸�zMd;�\te����kǤ7N�!���H� R��'�Wm�`I4��,�u
傊v��
��Iv6��7��؄X{�L�F���=ǳM��tX=����Ii;��[��'7{�["�<�6�~���A$uԪ=�[�],�(�j3�敻�m�ı�c���_��ړNJ�������*�n�[����#��Y"ټDg��:�LgnA�<�.sd�����$e�����VV[�ϖ��V�c0�d���̣d}���"g7j��{�VU������O���,���V�;�B�X~7"���߀	_�l�.��vqV�~�]�ϡw��n���H����ܖל}As!�i��=-�;�,�sS��uSX���G�����sXh��:����]K�O(�Ke~��=L.�)��V%�qʆ㜮b��+ǴaG���gNj��� �i�D�+$�3G���m���=�66��T���t�	��b�2����0KJ�ֆ��-�C2r��K����ջ"�X7aY��7U6�]nI��AFn�A��/�L$⼠3Q|�F�b�e�����"7d������
lm�Qd.�=���̔9����T�R\>B-��v�x�R>�*�i��G.�&	ub^�����O��-��+i���Zrh
Gp��"0SH{�ov��g^] �d����y�>�~�N�<��v�V�$���.zpQ��ث�1���� ���3`E�<t�U�M��F�Ͱ��oG.
�D\���G�\�f��Cz�D�����l����{�^��nG*a�|�|��{t���o����胧��ɲ�>E��=���s���R�������b���v*�D �/Q�u��_`nA��
G[C���^A�Q��Ȇϣ�]W��J\'y��$�!L�5��>f"Z�S�������#��e�5�*[]��%4Ō�t�V>?������kF8O�����|������6:�xɜ:�Q|s��C�^�T�?��r+�B�y��S��(�9_�̣}�V8�}�"�#��&*�����P6P��g�����(j�d�,���}����&ɢ�֜�� {�'�JSG���o7y�z3dRV�.{�vE��<$v_+�Y�o��Y���ٛ��:ߖ�+l���E�+�����]y�6W�]�E�tlN�:ǫoڻ
z@G�e��20��{�*a3��%�,����k��w��|�y��%�t_�f�|�8�@�ǯ�!c g<���=J0��@�Y*��Yj��n�V� �È�&F�cB/�e~7m�*�ձ����(><1�����y��<��Y�-�Q��P�t���~Ař;��e���@���2�#�:�=�ɏo�:��@��r�+�m��э�}οrn�p�Z�E�Z�Z�_z�2���B]ָ���P��x�>��#����@�S� v/��Y�������.���c�����<��&�c �$Ÿ"s�µ�|��>>�B@����<��;{f�D[`&�.8�R����ʶ @��J�*������uؔT��(">�XJm�(t�P�'݋������U=��I� �7.Na��|Dj����g=s�]�s�[1cUgK2�Z ��l�e��
��4R,��I����Z�����p4�"���K�8�T��S��I�ݨ�t������Apu%}����{�_^�#Ul�0��* ���[&-��������ny��ao����|TΙ��C����w��'�(ۂ�����U�ԋ�+���I�e`�cS��/��J>�_�����&�q|���ÉK}"d�+ä�>Vl��H"��*�����h�˺�G�m����P<�qqG���)�ވ����eun�M2%�K	yW@m�3��b�̿[��tM��n@�����*!AX_lk�2���$$�T��67yMv�f�G�A׬��Vc�t�� �*�L���8�yYL�A�_�B�NU��fǠ$�X� ��&}�&[�����¡E~b�v�e��Ic��#�*�;ǩc�}�Ӿ��bTRa����	#�g�ו����;->���7�\��4���VmqzZ�w��\]���D��!MVbl9=}����n�!�>S�Ij�t��1S>���f&�x3(�����V!4���I��H������3���ܶ�`�����;9]��HFc����م/�7o���2�vk�ƿcd�2����f���Ȟ���*Y�dd�cnyS��q�ӡ~]7����~_UvZ�T��W(놑gJ��%E>�}>�G�x�VF*/+I�\hI��W�s��ϲ�q?tPh�k�H{�%��4[��ĉ?���S��}�?�����0���w�/�I_Miy0�qSڞ�(��j��@����`���0p^O����7�l�Ux�1����5ld��癀���'�P)0Um[�����5w��y��`��h�U�}'�$�@$�Hޓ��`��Ԅ^�]�z����z� �E ���9�zgS�.H���X���]pj��c��?��O�[�M�&�п���]��݋T�`kN��cQ�N$�U��j�LG-묬��|Zh敫	�PŞ�"�tQ$'��8}ec�l�E��"7U��_��R�A�3l=��w�����i��Q���±�*I|��>J�F�$�t�بk�D�/���o�sb��5fH�6�k�)������������о|#�π��_��Z������ǉ��\�y)'�Mu`5@$AV�3z�`����y�
�?��P� �~LH�X�6�����\�z���tdv�B2��W�X]�a$��E1�[��g�~�h
��m[�N����>8tc���1���:'�ؑ>�f�m-7dEk�w��K�,��K<�:�>��N���ˣ����.!�&����17KZ�΀[���jEs�-�0�P|����
s �� �Mj��R���? c��8�
��N7����Ҥ~Ț
����2w,�4J$&���>�umL�3���.�u��NT�-_��ywHm�QE�����	q�6�
��L��E��8�3��@�R���$<\���7�g@,L�d�F�|��@�$���!˶g0�j�rXj{E����Dg�Zz׈�����b)ʬގ��P�ev?�g�I��+�Ņ%����wXɖ\Pf��ܯ8� ��/�]zI�����;yV��cl�z|�O ,�A6<W���J�+ܡ�9�O��; y�@m&M�Y�ɖ-�6s0���|=�O�K���v�9�

7v�!�wW�S	��vz�G��'��[�F�d|�)u�B���(T&��1\��a_�t8�r��Dǥ{�c�!Ԩr�$Q���Шļ|�'b� �K7A�y��W�����g�U�;@X���n�Ҏ�BOJ�����z���t2W锪�������A�k�<
������A�=5$�$��Q����,�5.@�c`����s�C�ubh����'�(�gY�)�s���NV_��_�I&'
�$��uloH���l���q�<��}8?v.��B)�����g �o��@.DA>�E��ֳ0U��T ���G�2���οǧ���\�vW/9 ����Oku\�_tj���S��U
�L�Fk`5`�,�F�פ�b�n�l��%<�ڱ�q�Vw�U����D�D6��ӈ,��+S&����\�;�0Y2G�
���t���87�m���O��]��<�L��TY�j��������r�|��7M�5���ds���&�tMW 
���u�+j�磴Szxn�f��u�E�Vqգ��J��w��X�Yǉw��;K�ӁB�p	bd��o3͎!�pbW�i�䩲�Ȼ����}GU�Gݨ�b��zAZĀ4�xl�v��,�A\���`�ӈ�Bq����5+�g�����b�S�b�5�Q.(뭪q�ث!���?7�Y��*�bu�2��e���k,���k�h��ށ	Hw{��Qtܰ3�4�[�}�(��h�4��J��)��'ʁ��!t4����H�m��G�z>�M�$F�#�6Z�*���3'c�5��,�L+oؼ��?Qn�Q(���>a�f^e�)m�2֯�S��_�);��#k��.��?�%�T�b�0����-��KJO�e�uo���#?�E~��i��o0J1~�ז��_��A����qn*���]��Q�����"A�0 ́�{\dw�M�2����/[k
^���ǩ�b7ۻ�L��:�M�+�ށ%I�=Z�+�����Qf�Cg$��u0��4(9N鹧Q}fza���k�Hӷ�`@�7:�nXeu��bG��U��R)uz�&��7�+<���4�$�\=�����s�J0��ة�J������!佯�^aA�x���e_>�T�ұ��'�v6�#*<���� �6�=�WP��!��1���n��i�x�$>Aq�D�Rh�ӷ�V`�GY��� ���dT�LpY�ho�NCT~qr'?Tvק����J ���o��	��5�׵�,���q^�X_�j�U��9�ݴ��u�84���\��9�.��g%��J����_4�e\.��Bo����Ԅ���4�o�O���{,��=2��C�#X`iw���J"e" f3�S���h�	;�Yy �)�5��J��M]N�������d��$	��R��W*��V��]����{��XFS�2m�o��ܲ���J�+�N3��g0WNr�d�����*V�����*
p�K�Ch7�N�����ޛ���� 3��g�M�t���7��ٞ:�����
�C ��Uf�w�O�%�2�M�GY�s^RO���h��U�zX�R�Qq�/~Qyc��"�UH���M�a'��бOVKjΈAR_�[�Q`���^��4�8[p��}��7� 4�Y
;�������!���s�9�x����1�Gw�س���<{�6P���" b ��w]W�~�I��	�'�g��u�X���L$ӆ����z������q8�"�U0�ʣ�&2�"��k	�����~�������uн"����<y��l!X"��	��*���I�c�kK�a��r���� f�Ǎ )�D�$(�#�t����sR�M/I|k�����s,���>Ʃ���;2N9� )�<�o�M�1鴃����e�/@���3G ��񛵅^>��h)\�17 v�I1|�v���w��w��l�(��P�<p��{�	��M�iw^��5������v�33�43H�9`C�������H^�U|��9˰���}
���yz�tΤ�O�l�������? 'p��X̏��0��=�ۂG�?����SR� `,���]qbE��Z�Vo���m-�)�
҈����{���p4ǣވ��-���4ҭ1 ���nF8�u��6�n�#{Cȼe����� �G޼��ߢ��Z�<	3��TZ��<9U�r~���x-:Wˆp�U���}C��*~Q=Ńv��D�R\�lY�zb�aaX��ɯ,+w��q:�	@�q��ľ~�tG�����q���t�[-�9o���9�u�I/��	ê:OPx�.�t`�pMR�pI��]"��
��L��Sr��ʫ�I~q\$6R�狃L֠����c�<$�Ǟ�M3N����<��"Y�=��ǩ+�)/Zw�6o^��rZ�"�p�$l��x�n�zf�^(X���>;Ƣ`�q:��}C�/#�FQ���!���+��1yiiҖ�RՏS`]���N�r
���%x��2]tC.ߡ!Wl-�颜8ɼ@����m�K�zǟ�-��	E%��3W�`�$<���%��M5XZI�΋7.�C´%���3v�2���k��a�L�7�/0�G�^�o[��e��V������6��Iۡ�c�X�/�~��ែ��z�~���
q�|�i�!Ш
7�9;J�7+�Mv<� �A���AN�Y�z�h-��X3�FbũKl�4�����| �����'�k�|�npA ��Rg�����e�#�Y�I�n&���p$N�2`;�Uɶ>���� ɡ���a��b�<�lk������Y�Ɣ�j�����`�����'��j�C�MN�	a�Ev�x=)M(�/Z|��s ��g���dg4}���֭ڜ���VYQ"j�ҖT�I�ĭ������c5q����ϛ6������r�թO-�^]�mTx&�c:�9���Z�vY�}���z-�y��}�x�"qJ}���_h��rn9�t��]"��5'Vkr�FG������4�uL�7iT�����<	�ȗK�{};fOMB�/�s�i��D�iN�].R�����b���A�'@�yA=�f��KŢ��ү�r0\��̸�xp
�sD�W�h;�9>��@�l�ٛ�j5���>�L�)�������0��.��A��]K��z�*���O�6�����3���<,+��kFD�	��e����E>@���Arlٵ�� �c_�x��85�([{Q�i1��"Z�t��d��5��w��b�r�Z�� �ϑ�ϗˇ��s���%�T�4�ʻ�a+����b�߹B��S��%r��QZ'��%}ߑ[�)X��h!L��RJB�,��^ώ:�Tx�2;���+��� �`����u��IV�A��4��1�F�_������;��@���RX2�W7� �
�/�Y��NѨU\9��#�5�KC�Gq�ߝ7,;�EF�^�����W���mJ�"��!a:�6.ѷt"=�#��x��!�q����a��H{w�r�U>x����̿����fȯ�$�!P��_G����b���ꜹڐ�d���چ� }�X�B ��:���)���!Ů�\��q�{��.���FiO�%3�������� w����Z�N�f��Kp.�>���Ĩ��//p�h��U/	J-j���#�Ww�Y^a��b�}�9!�]DA�.݃|{��<�(�#�Z��<�1僝Y����ۮ,�ͤJ;�Kg����*��|O�&YUu�jkl��j
��b4�`Ż"�e 9�l���S�ME|^�Sf�m�^Z�on��V+��������G`Q�ɽ�|0V���B�&
�v��	ul�iC�L��.ը����2�n��]���������!��L�#�=��նYb���������6�+�=_�밸~y�3/0+:V��h��%��,쫵]'��#���F �I,����dD��3��7�;�$���]��Sp�D҆&��/���>M٨�۽�0Awy �$s�4�X�����9��!���46���C-��,��u	��3+\�z�W9!��M<�ɳP|�чa{��~��n  �ⷕ'�*=��,2餞��n�)V���%���O�zN�Sߝ�,է�h16:��ѹ�E㛁��~.n:(��(t}�h�a�Z~?5���N��l�ᄎ�#�	]���r���A��L=(I0��Wc�����5Gp2�jo����TD���=)H�r��wz*���$���KF�LE.�)/.�/��
�¥��&~��b5�6ƙT҂%"��H�
��`�^���C�ɟ��3���:V�.L�z�,X������U!|SӼq�"N��K9�px�0j;Cs����g�/��^��;3���h�@F��o�t���?fI@Eh��qs��� ��(�Q�'��uv�P�p9�4���<����!�P�؈���� =��H+5q�0T30�Ⱬ���^��0 o�@�T��=pļ��ច��j�%M��`a�SIs�7���
��:2!� ��t���"F*5i��p�d��,?8�[�D3��خ'����%4� uF��5������{�Q����sLI�v���V�8A�9���PF���F�v��Ȅ�u�L�dNz�<!�H�K1��9��M�R�}	���}����*�wS�#[T��/��g���k����&��F�
�9>(T���~��xZ��;/2�h���]��V���e'�����\�y���)m�_o@�ic�)Ԃڃ-0Ä��lX������x� rX��Ϥ�Jq�	��ڦ[C�|��NKc�C�}?� pi�W�9�=���;�-��l����K�K��pK�YY �ȁ	�G��6� 𼟢�(('x���Z�Vk�����̞i�Uv�MpꭌBؒ���<~�O"Mm��B����Ī_�i�P�W&�7[s������DQ}��v���.��mhKv*,�}��+��q' �4#�$�}�I-��5�"+�|U����}1���)vx;b��t���':�#����s@�gd���:|\�b�]Ϋu�7(�0�%>9ߖ*MN�B���$��L�P��}?sV�Q�[�].����c�e�p�^�f��{��,��b��3&N1?�m�"�"bC@k^�ȃ�DC�0<�eCx��h�b��w���K1,���1V��xw���q�i)�YjFf?U�N�It�tw�}�]V�Ь�R�D��6a��°���/^�̝�b����eGrs�)����z6t���.���p�<Ω K�w��7�}�+�4i�E�0�l�i�� #�h�'tV,6G�}uI���>u�!�o��0H��k�2\�E�\��n�'�dїgp!QRL����w�>��M���Zo9��4 �)�N�t,5����cv�i_d��肪��<gh�2N9a�B�P�?Nm�EP�,�q��閡�*�\�uޟ��I���d7�))��&����j���6׷Y;�����	�u���纐��5����?��� �O�թ�4�"`��J��pR#�{���tBC6��2h����&�� �:n�
������=���8 ��G�m^������tvN���nQ�o�SimS2�����,�Ѫ\����e���6�����jS1��/mR0S������w�ҢS�g���C��������6�#����>�5;��#�>P*2N$�y��X��%��9�@}�*7W���zph�&-��'w�ܠ"�r���'��UV�n��F1�<�8��1�I�PD�9\v��<���/&i�.��iI�!���T��%up?.��$Ș1��+B��uxqģ�O����'����a{!q-�C=��c0����a��|m�O��E��W�r����0�RM�ͻܾ�ߠx�~�$�[S�M~�/�1�cd���/�rw�;��Uz�!NX��N�jį��	Fٸ�BO5�*Ns�|.��V�m�q]Ǳ���	���*�a; ��]1c@勚����+@!�40����s׹	����C�ڋ�`"��(�l��T_�Ћ��-)�M����k �s��8̣��W��2ȹ_��V� ��2r�y�1R��r<�zc�4�����X�h���=�b/��|�l���E�з��]����?Ъ��4�1�-
��6�XqŅ�<��d�Tl�-��}�X����@��׼����"�an�ۅ�'e:�Bp�֥t�w�nK׊#�4�)�ǫ+T���yL�Z�JB��]�U����m��F���@0A��`mNG&�Rj�x�&�F��Z��*6䡘�g�{�!��q
�UTyvi��HN�"�9W1���`�4�o�̴��L}H�^�A֎2�D�.����@��z�6�{��	9�/W:1c��:C�$��coP�Q�Ÿ�a=�hT���)z/#��1マ�,X�+,����[�u��R� �Q�����#�e��Su��������``�ݓ�����Bc��
�z����� ��Ɔ{鴐�=�F���<-�Ww�KV��t�e���5Y��7S��+zC�U�� ���U�~u��nC��}%&xU�I�,�"h�ح(�v��;����:��O������T�9�GT(Mk�1�e�ɢ����n�j>�uЬ���}��$�h�b�D��7ԃ�g_��We9�y��N�>5sn��(0��9��x@��u17� v�]��n�(|u�؀SQ\1l31��)==֬��>�������l�;AE~�H���S��?8~$�g'����NO�a�O�.���*ʏK���z���\��J0�b^v�$�2�������ęb5dr���,��gkh�0)
�m�P�e,�S�l�o�����;鸥�Q$����,��E��I
�Ź�s�$��Z�@buŎ�^�GHo	I�H�=�D��r@f:.�v�Bto@t7�;퉦��O? Y�}� P����ꮹr�G�R�t�q���):C9�/T`�3��s5��NA���S�
�>�60 �?W]�fE �`j=�Y��%(����Xrk��c9��۰�&��&ŜL��!SH�`諝��c6�?�Ȕ<۔z�G���f�ά���N-�nm����gڤ%�����<:����%�m:��Ǖ���7E0����УY��C��b �k�ʇ�����L8u���t,�\���P�������CYQ^>(��	z�%9�dt"6�ǚm5��='򽫮��T�b{�X��e���@������ƍ{�o�i�w!�5TaW^Q�Gȍ���ls��e�aj(��v'i��P֙A��xmB"Yw�rr��!,H=���5��wX<Z�+�'�FјK_����=��OV�"����uw��
"���>?CS�n��뮪��(��{�qQ�@���+��$$�pIa2n�X�)�p�%@p�|
��#�X�6�#mg�p=U���Due){��*���G��Q�*����J����J�(�Rr���=�]��7� /��9P�cX{-���0%�j(��}.�s�gA���\[�#Z���H�����կڣ��c5�� S�5��d���Ez���NF�&�g��Q�&�(=�\?t/��J)ŗ���70m�)Qrܽ1�-��j��L�A����i�fO����
��i�L��֖bW/�XEt*ꤠ��K�؝�@{ynО����'Y8�~���G�ƹ�_lE��g
�¨��'�'\�ʄ2�0u�h���2�+[��o��y.����YD�]7U�ɱp�!�K�G$��A���uj�҇a�.��zOhz�L����������)Ē�︜E5��g�1�+�2�#]&�նT���pks'o8�:�D%��� X�EW֙��J Z85yT� �@��;�m�f�po粑8���DZR�)�i�ˏM�&bE�����
ת�#��GS]�b�w����C.W�1�������F�(w>AI�};��̪���	���DU�?�j��d�T�p�＾����L[m�C �&n`N��BE� ���D�zR)��C{&n�~���c��WM�:�0��.�;�0hJA�ՈV��[�JQ	�U����a��-Җ�g���P$^����� g(y���e/5ZY��H͖�0��Nɏn��"�	�}�(yjj��酭�[�+1C쮘�e�I+)N��C���E̸���w>b���/p~r �J^��Y��{!q0*rW����"����:�	�q��[��A�b�&��t���;b~�����.z���	��4h��
 1G��"E_�(|�Y< "���k�U4ׁ�"�r7�<G��Q���Yo�'��&����
\p(r�t{���p�l&廙�*��>6O�*aM�W;�d�q�z�ՠ��@-��¯pD�)�zT���Ʊ��y6��|�wٞڮ��LW���+"�z�-�*6�����,�>��K���x���2��)��Bf�kt��ь��>q���h�Ɂ�r���G�^�2Q�gQ^�dL��LT厍m�4�hR������R}����������-_��cMyu���L{�=��R�v!7����r��l�;�t�}�ڕ�Z�p"o��oT�L��`F��zԇ�R�6A��Z���
�y�9 ��m��-��;�9�CuT?��Z�l��H�/�l� �<2:폒#=S��|��γ��r3ߜ�x-H�F�!�PH�'H��;�-�;�iMES% _��v"����������O��G�<w�O�e?JLJx�q��><}(PŸ�(��\5d"NDg���z�����d�hL��D�a�f��q���g���n�v��g�/��b�6'�7�)���x,���ϫ��]�
��O�S�A,���0���	���r<�±C���!�q#s��W�9a鳕��5�8�^I�n��o�8��a��5ƺ�i��E���tz��T�;U�P���ho| x��w$a
�䀹��~x�/udt�����mޓ�s�r�M�mL}^�A�8���GHgP�82�
`5�/��Lxa�j +�ͻc���#n������P�rg��(�X��~vD7n�+$��Qk��B��|���0���rd`�����%	4a�v
��GkLQ�9Y�r ��Cz�8���'��쫟�� �vk,b���w��r��~�І�I���T�X�Jx �p�Ng�A��8M�eq�V`<�j�*� ���UA��3�����Z��H���8���CQg��S~�OO������(�`���Wc��0�FR<Il��Q�U$�#j�ϗ�U�-�ch	v��X�I`���.w�>1c��g���r=�*(ȡJ���_.�8�f/��E�����z��I[�=��"eś���&d�P�n�D��d�53u�8D;�����ݪW������b�LG��Ц�L�V�ʎܐ�=s^������ L���|�qZ$���{e�ӭ47EEu�{���0��q�demQ��Smx�'���,�����ږF�I��X�����h�>�l�w(Kה��z�=\Y�!�ef^�4�����X��Β�I9��j�Z-�}��
�Fxڭ�������)������W��lyd���fk ��L�ѣ���5�:F�3��!��)��|	�6�?<�$y���fG!`=��|��횃E�"��(�	�����3o�d�t�`j��{dy�"��9)�vݱ����	���c���ډ6�Q���'��?]gZ,�	��ȋ���8`���rZ{g@��i���s��l|93�*�D�Wy2hPH�D:�0�dE�A.�<T`�� �]Np�;r�F�֩,�7�� �h�&�Z��Z s1L����pW ��A�%:�B����5�|��.`��*�Pɤ�|�G��LJP��Qd�5��\�=g@����,�ar�{�(��x�~�/��Ҥ��.��_�	`�G#0�)5M�=�u�3���t/�̳_w�����"U&��b3�u��p�-B���B�v p��ji,�KF�$���.��om��I�\��-A����0�.fٔ���:�H�ɞZ.M�0�<�Y
�����S�2R�۔14�P8��53x�4�8s2�pmx�����D[S�W��RT?ȹf4�2�n{HB���#i�����i��3x�;ix;UG'���]� e�|ppC:;�-�E��v,z�,�|ꍘ�̝} T�I�&b��5S�z���t�]��M�A�Ɏs�X.cA�9S-��d��pMr���A����]�����`30G6j�� �n�i��b#�[y�$���@=
'^��dRL�|̰N;ߟe�zc�����Xg_c ���3��<�����D]T$�:Y���o��e�CB�$�-)�	�����]�=�GÛv�u���"��K�,��yʋNp��0a(�����/�� X|�ezh˷E!����/�e���A��U�BG�p��-X/j��i�3�c?����%2H�׉+����g+v�;?�h5'.��7S.�QƵ��_�����n�`hܚ�����eFwk�
gK<؈�T��U���I�s�U������x���#��>�<���4F���L����gD~:���~��-lf�A�u��p��؟2��M�-,��I�T��Z���'�� ;��t<�Ù5e���m�ä��u}.5��V���x��j�,�ᕪ�p(c8��pS@�6��Bf�5՚�*�C֩H	~�g�*7yu,삟2u�����b�r���-|�D,}������Z�P�=�	9I���4�z��#�}�8���f,N�i�$y�� �'�@י:&Q_-�� c�Q�z�xcΉ�7�b7R�Yo���\� �H�S�4�_�4�}|��]����;,'�2}f-�E�xJ�8��2.�[բ0�d-�h:]N��;��؋ޣ�� ��--���f���r��p����A��/�J/s�87�ݟ[�>y�m9�k���,te�+sh��W��a������Ïg�a��:dF� o"~<!��GG^b�� #�ڥ����,��y8��udl�i���ˊ{�M����҅Ɂ�S\8?���e�F��Z9&�)��V�E�u�=z�V��^��|D\E����X�kk���4�K�|s���O�����7�"&˽�����'�I���4�΋�*
&`NaEw�'��<�(��E������ֱ7Y��T'��%��6u���i��"��K�;�_}
�T8	O{-���	U�:L�AnoI�����?	:�l2,?9k�A,t�+0պ'^�7�R��x>���~�=(0+�7��ɡ펊�/_�(�{�M�ˬ�9�V�͢R	�7	��-�A�'�d_-���ri���l�@+(��[&V�C'��[$M��&��	�cK'$u_��`��s�ɽ8�ǟ�m�&�!�G��dB�Fa¬�����5j�r2�[Z��S,7[��o7�
��q{��B��?`f,s�J�X&��51.&T������&����O��t��I���0���+�q����kH��Q#��F�t`U��k�N� {�H;��7�(hDզұ>�	�'���`��!,o�}���L�:�33��ڢ!����ը�<�1Y����?L���$�	�]����r~!��e)?���y�T��&���n�N�����5�X��oyJ�ZBU5(lXrqмN�L:+r��C0j�6���	�t����n!+(�B��S]�բ�ǜeCAt���������I[W̚eZ,L@�b�0n��;f����+9�kG*���۰�}��@L�B��.�2 ���Aٵ��v�9�w�u�/��������ɦ�����^S����V��`�x-{�	�|�>�`G�n	m��\ lҼ��XHڅt ^�[�0�����dW��5�p%�l��=K�?�_�Sy*J�7��������y!߀<S��4��|	��S�<����@��
Ὄ��n3w�Bz����娂� ��^��T<|�Z$��|���.)����;m��NPq6�Z�����4���Iw������.~3���n�R|�R6�{J]ݴ0�O��ƍ{/�%Go���n{�7���Ј������?�m�Y��D����"
�m�YX�b,g�뗹��-��˷Ԟ�A�:Fh�k*����/��/��i�
A���**bW_�� ��
a}x�ƭ�/�P�����" �?�0�XpIA�k�忽�VJ3�m _;h�e���EyI��О����0d���{���\��F6͚���6Ĉ�1xH�����۔+\�& lHۛ9��'���Bke��s��������_��owlh�;pӔ�@�d��3.�A ?�m����\�g*��>*���*���K��㖫$�� ��R��ɭ�
��[�m��Č+tX���r@)�g8R���>�M�3p��4_�|%��$�ETvߙ�c`��a�$�$�:�|��ta��U` �s��:�	�����c�s�p�jѫA����ڔ��dj'*���ԡ-����ܛ@E�$���AG�!����v�6h�.�{�ń}�W���o<Ww���Ď�Cyteb��aRJ`�5p�ڸMi#��8~�:>oD"�N�W���E�������_d[�tLJ�N�ܨ�{|7�B�٨�𪈷T�ď��Y6ch$�'�i��
	����2�g.A,���A�"&a�Y��&[�}�p9�B���A�d��-:������-�����t�Ն��~l_Ϳ����EoJ.�N�O}���^>�D�Hek�7������35ud:�`��D�bU4����".��|zE��˱:$�%��͔i:9і��/ccOa�z�_H^�S�C{�.�G6���?	C��2�ڮ���T^��c�0Z�=���@)���qg�ag���61;�N }�\��G�����R��ƚbK�	\?�~.(�Aq���͑���~��+Dh��7�H�:R[�k"�t�7���]�����HP�����>Td�'�x�&$dC(�C1$l�Z�[����-��o�(�?�-��gQ0[�W��l�M]7�)���)AU�Z�=�ő*�|�qV$��B��HU����I��b��ν^���r�����n��a�1*��z���w�\�Mm��t��Q�X��U����<F`��7X>�-|b��{h9ޥ�1ս��.҆�iʓ%�ȝ?��B���]���BI92��H��$����t� HG�?R)�_��"4z^A�blH7�e'~����6�ET ��UB�����c��@3e��0��F���*���|���1R�ؿ1�ˇ[�i~7mF[�E�ԣ��R��:o�t�yrA��D���lzt�R�n���[�ݫ�U�m��#���U� ����6���7�I�����Ǡ�B�b���v淇 �$vƅ�TPQ�F2�:|��YF����%5��0��kͧ_�}-hF�����(cl������4�x�B,X{��lΤF��."����R(_�F�5H���m�����F�A��S1;��L=�w���1f�h���j%T�b�N��Iњ�w�����,�ɮ��tЌ=�"z���qu.;gT����p�O>W�����x����M�����!V�\����Fu4A�����݉�M��~w�J�*�V$��k����̐&��Ӽ8& �q}G+�,��[�W��Kk	�F��1U��+u����������DI����������K��S��@�Nn�(���G
9�ɒ�5�II_B�9��ќ��c~�5T�o�m�([�@�6���I�^��6��'��0�z��N����2�G���4�3I%d.��b����XɟX��t�Y�����%��ё����u��{nFv�3V����מ "��?�P���p�O��Q�|H��榾9�9��3�o$!�6��ci�'[&b/y��j��y[�S�WO���%�9��Tۮ-	gޱ���R��tc����0z�b�c�{8�=��BMt��dܠE|O���f��Y��L_���t�g���J:��CH��Nn���p�wO����=�&�S��?�&4�[fy�械NU�#��K�`κ=	�B�+w��I�z!=_V�+�G|��/Sk?��Bz�����<�`�6��� ��[E�kBTq
]��U�u�Q�]6Okus����o��@�V��f	�ZLvo���sAt�EP�i�}s��Z0ϫ<�7�/0�Q����趱�>��Wȏ4 ���&��*���s��:~N�ѷ�\�%�%�:��Z3� �?�_��m�����WfXN�'�%C'��Hx1Z�.ȿ�[��-�I#f�\R{O�Oo�T��^���T��-���C����ǅjWE)��bLy[�Hs�U��k»�!��X�S�[�'@d4�J��C��zlI]�V-��$BL#�&�ǐ�Z�y
'�R��,�.(�6vܻ�vs@;B�ٽC���1�TwۺŇJ�����5�e�_�P�,��|3`��\�^���j:(����'_�k$ �F�`L�,�x�g��i�tJ�~L��WC����� ���k
���X�����D�3�9ɉ�p�[=$�U�kҽ#a�鄆O`�U��b!�
���[Mf�4f�=��iz7�Z�ɥ�xR�,������ˊ	vI`h�D��ە$��c����,������3u��B�"��O�ađ[�Q�ș�jennX�v�5I��p@�8���FD�R���=��bEa��]�NՒ��6GB�5Ɨ�r�yʸiV��C�.8~�(��HfuH��Z	��"����>]{�q|��a/޶Sn��s#�N����8�I�ث;����|NF���B⺝��k��|���c i+	O|�C)��Z�U��D-�3� ~�G��[�ejR���uj�`21f�	�2{���T����/��(1��%{�`א??ri�A���ß�p�*݆{�r����n�1c��%�%<�4�_�E9�f��Qv���c��.���m����R=�?�N���r�q��ɀĉ,�L��'���YT#���@��=��2a���"��w���o��������K/b��5f�p���k���NK�Ф��d��Xs"���>���k��{�|�4F�>�ؑ�,ǧ�iF@3N�&1K���}�J�Z{�	��3�M�ߵo%� Y��)Q�w�E��)7��4e �JD}�3�$��l�K�!|4���2�wUd�3�߿'�.�m������	�� ���Ґ�!�g�m+bn�� �F���FDqW�Ҿ#y��V��ʥmc;�&��9��[��ݹbA����H�H����e��M��5��������$��N���ZU"ZX��g�S+3(�F&H�O7�g�j>G��O�c���^�E\�<��W���2��aF�u2�F��ԇ���@M�C�hCg3%���w��|�Pd� _me��T��6t;��O�^[5�3�K�8&!���zgͿ<��ϹB<
���-	��>��]�՛S�i�%6@YI��ʏ�ֿ�C���X��(/_L�_
1�oCr{^ՆƔ�9�J�@r��g��#�3dZ�m���U*1�P71E�u�|Gg�����u��9�g����ho���I�2n����J��T]�
���*���>��0�V����"��S��J@<#1x�f�I� Q^D���ou�C������ y�(nr@�2I�~l`&�a�̻�u�o��%g���M�n:��M����AE1�X�F�l��.'Ó����x8񨇋#Z��Iz"'�"�j��_0T�9�\N:G)����E_1�}/lY�Ӯ���3q@g��B�=5��r�Sd�|̌FR�4H���s�h6��������0V�%�
��v�?ga�����'	�~�P[�q���<����yt���?�𵇇�B�x�#���]�jM �H�[�0D�;�Q9(Pd�� 7}:�h����7��[!�RB�3,~�wI5I���i�l{ӥ*M�/��S��Vy[�v�pB���^N��9QN��٪���� ���E����V�)���ŏ�$�K��)Ցuʰ�f�iu�"��Ӝ缃�v"LI��TD��j�X랯u%ҺwU�����j��rnYl.��k:�bθ��,�m''x�X+)�
.Ѫ�	dEX�������H# /N��xg���c���ۏT�
��@��z�x��Ju�ǝ�-����鑨Kʑ��6@	�X��M�)i�-7��m������~M��+t������{����p
���0��Ӽ_P&�n#�7GO����=��^@�W-{>{N�#^��K�
��W��}R'C{.�j�A��5n�����1P��IQ&c|� 枇鷒%��[<c�^������'�˪F6�o�tL��b�$����N�4��m;*ê�*�G�y�_
�����8��l�[�,~u	P��>L����ՋH�ھ����'�+�
�k��6j'��%<3� I$I��sѐ��Pbb�q��erw���^�鉫.`��4٩�V�&2.K�Ԥ���h��>�{Y�|���$9�R�0�#�>��E풌D�9��І�}����/��@L4�h��~�����EEK8�F�+UA���) �5�koy�1�g��ɪ���ڧ�|����/�����R'����y���[
��P@FQ���1��;��iEƾ�d�]%�|��:݇9	�4B�;�+����*�}��X'��{����Ӯ�u�믡)�iR�k@0��!�+��}Nܮ߆B8%��-�\���i�%s)#��I\_�;���V�^���$�e�`ե���"��*��/��l_K�i?�̕�)6�4gģ�^���쨔FٞK�/���<�OT2s�)��t{l�����Y ʈ����d�eǪjp
,[�!�?\�Y�r�s"�|Ƿ(�8�F}���[F�c�Z�cc;�P�t�'����;:��+�����ѥv>G����K��9g'�Xm��K�~�\vQ<}	oM�Πŷ��ծ����PWG�+T@���b3�b���>�2�^�W*
.i0�|y0v
_�1�\���k�$F�VwW�����Sz秮�e���+�tL�F?3b�"��L%w�mD`�vO����,�	x�V� ��[i*��i���_�;�lċRg�G���AKP�{^t�Z�vf.�H<e����2���]�H|nZ�i8�Zāe	o���Y�����)i�p���9�r�ʈ>C�~�\��LT�SA�gD0��f{��/x��%'.�5@��(� ��,��N܀�k�[�*��&+��~v�Ԧ[_x�$�	t���;��{U��E�a�Q��S�"�`b��H���W�^��r��3�'j���3
�����Y��<�x8=k�z�	�[���d��:��{�����	/c��E�&��6=�4L"��ʩp���~_�p���*�ْ���:�U�Ñ���4*���`��VvU��;�'�P�O�iJE�%�9���E���H���G
�Q��D$�eݒ+���ҿ7rP�w�ڴ�ݡ²f�Ri�!n<�<�}�X�=��0�Ap�P�u͑v�ճN����*F����ށPg�"$J U>�M#���aԳ��������s�~���Q[�y�����K�m�����j�dc�K�������4	��# �kn���m;�d�1������t50�T�M�2����E�C�rr���{c�������⯌	U���W�t�S�ށ�d�~i,�X,��8��Y����-M ���+1�(*�x6*�>�W��p��-ܻ�D� s���3	p��w.v{^�J�.î3�
��cN\4a[��<s�9>A�P�TSx��&��R��G�}�'z��)h�Ss����(־91�F�»�YK��+���@�Nmm=��Ś�/i���H��3��?%t�P�.}}��C�T`=��Ft�#뻎&M���%��M�۱{�y"tRe?�i�ݬ�{UE�(�1�򠱪``*E�����e��}�����l��K�b�	��60W���Zأ��G�N���i����5�G�����U$�T1�X�&lA;�7{�U��㯮���l���@j�(��#W I�g�!!DBf�:q��`w�n�M�W�3���Ӝ�OA\��za}��E�p�H�6 :6���e�n4+����H�`��3��i���3d�R���� ������`�K�(i�����Y��xp��w%�/ �~m��j2'ddP"\�c�7@cw�wi~���^���Z)��HP'Z�W���P�r��h�a���8�XaҢ���-0m#gF����!0���I�����yFy��uQ��&�Ǎ5o��F:��C���PEi�r� �cq9qq�g��]ł�����i��=D�n�I�T����ør#�ߚ�*5�>k���w��ڞ�Q�l9��Y�M�q��cr�U�a=-'�jF
0���O0�׫h��^�N,�T!F�r@iʒ	~�1�\�ȩ������8�A�{_JO
�e���ī�f�9�5%}����lN�Y}�P�Zn����p(@��'C$5-����z�7����Ʋ+�M���ӎ�D,<�R[hn�8�JdM��u��q�-�~޶L��޷�4�������CQߠ��]�r ��=TT�
�$��jrA�Ů���Y�+ϐ�&e�+M��D�H��g3׋\�0E�6�Fb �M�7�Xk�8"�q5��H�d���Y�~ �����<L������0~�Uj�Z���y�!Xꏳ�IV�,�d���u��f��I�dguJo��D�'��h�#�\�,/D������#�f;���z��9
?�+A�����|ʤ���"�-�}���4Ra)�3D��ER�����ʌ��j���<_�ڣ�#��#	eN��ry�zf�I���Ű��.��N�)F�l���(¤ ��b"�t�P5�I�խ�,��yck^��e��	���j�zl�V�h�Qh�GX�E�"U�@�hh`B)��F�%�t֒�́�\V3U�M%�C���e���^���(�w���-Ա+�[	T,����n�G
�¬��v��@#A�MIL�zȣ3	�������l��>�,G�(��K:B�;ݭ����ϻ���_P3�����eM5�wc�\����1i0���dl��GN���Q\��W3�� +ޓ��a8��9h7��m`�R�iU[��YU�.b3�)A����0%|�x��_K�=�y*|�A����B��(���d�SY	�E�BC���o��xhtO4vj�/�:U_m����B���rS����e�-8ַ����6��KX��zq&)q�������7l��l��*���Dm��tӃ|񅮭�&۾�^�;����s<,�ٗ"o�(�|���b�	�����>L.�b�&�Px�#���)�ڻ.����0c�$�3"�qhH��� ������4W�����:PL�OS�B@�R#t��Nu���M}�Sl*kK
a$E����;_:Փ�46�؃+�Q��EO�ԇ��8k_5gl���s�_'φZ��8@"-Uv������t�E@<��W	�ޕqwM��L.Le���ƃ"������1�d.#�<t�8������F-��A'�m%o�<��<he7]m_;�d�[o�s$�?�E<�T1Q�d�E�P���y�����"�E�!���Z_pO���}����-���9Sa����>_�_�
��6嬾��`򿙾3Z0�E�O��gXxu�:�?�4qo�\)^j��&E.c�c�7s�6^B/�:5��:��o�ɞ��1�~�*�X��R����0�S)���Ӻ4ʙ�F�'X"6���\Y�^b�|~���O�=ӗAL����6<d�OguB00
��o$D�Uhl�.�ҺC�d���W�S&�	*�3�^.i�m����K���Dl�5ċs�@�e�yG��I��\�r�8�?����K�ꑨ	ӍD$�HC�4z#7hQA��20��<P>�
6��,�>C'b"=Ep�ݾ��A�y��͍P�1��C��V��%�tHp����B|�'�{�}��UA�����?�b���:t�!/�`�?�E� �)���=�Cz-iIv�,K� Z!]H���!}��pZ=�r\Ձf&�te����_�'�#C�Jj�����e�yZ �[����9O �TB�Ul��"��a,Y{5��@�p����=n�����?����)xd'<gy2-\IR�k��=����	mz�'g��sQ�R5ț��xD�K����8~�ޔw�`N���3��ӹ�y���s7&���� �O�D��_M�=��"���eé�`�;���BDbw�3b//��2¾�ϖ=�MÌ�oǖs��9�,&o$�]�g4sH������"��pt�<�7$�/��Jg��c�X~���lz\���a�����t�FQT˝23Y\�<6�S��;9��0}�U��s�v��
v�@�Z �kiY,K��]���cHpoP�UQ��#Ϳ�]�ag�V������)�g�wY}<E�H�t�Fz$�	�S=ou�Vmӽ����Ԁ�$��d5��. j$+1�$�2�S2\ �s����k�Js���9�)`j�|�p[k�8����B�A��k���"�=@_Z�v=�>��Îw.�-P��2�g�����v���@zwD(��%ds�u���A��\�ɗ6$ ���C/ǘ������OZ\����K6���઱.��\�}<�j��X��f�޸iSA���n�}pH��ed������iheݯ{H��R!�"'kZ97>`k����5�s���ȷ�|4n�{8��<6���ޡ��0���@�d�SJ��D��eO���g��O$B�t�V'\lb>E�Ym�����Q�$JZ�z&\u�����/�/��Y]������eK.,���ْ{�����mb5����t�*�l�����L5�K�q�U�>a����jd6�Ϣ�FT�$KY���Kn�Z�\.G������߻k��8M��C;FHʏ����VsԈTo(�1�W��Ҋ̼t&:-ҟ��N~�wϢ9�hd3X3d-g�K���598aOVr���͉��Tor�[����C����Ӱ�s2�pB��J��2���ֈ0v���H��/pD��x��D(�"��L�3���f��
�NV7��F�-�uڥE�'�Uw[��� J��{�zN���G�i���ip�
���R�7I(M�y�yr*�*��a)�_)=C+�i��橋Ƃ��>�WB}g��)ȼ����"�@3�aJ��wk����<A��pA���;'}�$�����TXk|tY.~qsK�y������B6�/Ddή�ˡ҅֋�]�~X�{O���sM�k#�Q'~�p��	��<d��9�WY�^�݅1Y��91Қ��A�8 ���
�T҇�0S�2�+�TKm���I�QJ�3��Z�eO?��ܭ_�	.�Z�0+��C�&r�)`���g{��p���}�N�������իUezlI�������o���E:� Y��j�����S����/'����V����=_�r6<���Z�.����!mՕ<���y����DZz��`[;���Ϟ��H?��*���e<��:�2/��8ױI�އ���U0
&�(&�G�!h�J��s9 Pe�����~&��ZL��gg��1��W>%j�[?�b;E�W�`�����f �@X������*1�k�^<�0"�Y�`U��T�ґĔW�4$N�n}q=(J�*$�n��F��gˀS��Rܻ�w�V��m����. g�#u5�d	x;��5��*��ٽ��;��&ȀR������������8/a|_B������*�^`�,o����g��^C^<��TXb��9���8�~�$th
��O���>ƫ5aX���
Z>W���v�&rK�뭆���NYd�4'؅{��=ZD�q��uY�8�8�f��f�������#k� 7�jn�������:D�%�H��A	y=�k���S�F_S!>����Y������pepʜ3r��s�����T��0ִ��2$�B��_s���DW���O}8$�8w]�I�����M���~���?��3�n�����t����ڣW�~�������d��"�'��~�j���o�R�'�l�<�v[�N`a7���Z=B��&¹B����{���2�`���ӖM���gvPJ��u�^�G��]����)Ǉ��}�"�p=7Q"�y��"P���K_ek��9��K����KX�?���&
�]���{%�d�n���a���Y�a�6�`x�I1��"���NCen�D;*�c� R��i�2��0�~�WK��+D: ]�#o����L�q_ n�Z��R'!0��r�����І����d��&��~<��*[h;�F��*3墇�9������y��`Cf�Q+��d��xs�b��
�\����?�`�+Ò��8]�p?$``b����� g��t������V��gB4����7��6?w����#�t�4�C���p"���`��p�I��ݡ��$��f��O�ի��S��o�G-!��V<A�շV+w�8�b�G�����;q{E�PԪZ����܁#�sH�($7K�$K0k�#[�M,s�0Hs�	|�+:A͏�ƆPN0�n�4�]fJN�2G�7iSǤ�xZ��H�"r y8�ͳ9D#F�Ty
�������HP��z>�4׼݇=/���[�f�:�<�1~~$qH��ߍ^�OG��% K��)q���(O��s�0F�t�u�������U&���[�"�J(��m''q���q����~��xk������	\��bq3c��PH(�Jg�g�c�A�1)�u ujrh�m�����1F9�ǟ���}^���/��ߺK��Nvkek6��>Q녗���/O�B�_�Pw[Ԍ*���0�=��?*���l��pSAS�Nj��7��w�Bn��El�T���
S�7/�ޏ��J,~W2t��S؃�bx&�"�s�́X�[�TDUH�6E�E%���b�Wϡ�,�A�OuÖv�&n����H4�����΢��`,���K'�Mh�����g��m�b(w#�DTU�e�X}�TV����\���vzᰪϫo �,J���t�k1':D>Mu	���Ig3_�-�^p�b�8������#��_�v���tD�J@��9m~�b1���u�0�?���S[�Y.6>��+��bN;%����Hά�R��b'a�	���qt�o�a��qD�e�Y�hGߏ]�z�t 
�Iy�;�1���Շ�è��BL2h�v�^��֣~��"β�O�%�q���(����;��P�����z~W�q���g$�"X[���ǽ+�6����`�%�i����r?f���@�o:p,~����&�Js�@��]��р8Q��6����Jr0%����c��
Y��Q���r�.h�Ϯ "֎��~ 7n��ҶFO�Xi\祤����xL�p��\j?��b�-uV!���lI!����bL���s@�*C������x�����Ec)X�` �m3P��<ɬ{�-�;��=�0(
����g��.����~��*��VVF�'��bO�����`/IdY(��������gPʪa�ғ�v/>�N^�Cl�vJ�UB�lI������δ��v��H��R�T�5�f�{(y������	Ӛ�do3�Luў������/ۑT��j������ >� a����8�}�� JC��<��w��S���&�.pE���~���-�.Rq;؈�����q�m��W�lLY�DJE!˒�@a�m�@,��?��������2�`������F�	]�j)F�Y��L��qJ8=��������b�+/O$����LB��	�����i��r �2K5j@>���ɏ)���.>D7�e^����ȋG9�A�>�_���X.�5Ё'�Q����f y�}O�/	1;c��p��p(Zv�a;���Qй&'G��BL:�ou=k�Z;�_�[a*�?�(���20,^Ԕ����P�e���{J˥]����A`�����&��k�(?�#�ȣO}��,�}J�>FN��0�>�Q���NI�_2T���B`y<��/&�Cݨ�3��@�ӊS�o��Op� + e���G�� F�}���a�a����`�v�h��!*x'�~��'��9�c3�<n�y��ٲo���d;%���!H��>P99�T���+�����P� ���TQS�Ɯ�?0%I���t�}�xH߮��ց�rӔP���BG�*��y�(HhԳqڇ����]u~�r��HE|GE@h')Q5֝�(�o�8�GX�g�Fd<����g�Ι���RZn�-�@H/֏��LQ�O�&PL~ܠ�SN�=R��)p+\%2��a[h|��og�E��ߴxh����D)u���D,����FN�h@��>Zr�����]�O;�W3.H6B��BLx�t�䷠g*��P�ޜ�0�%0�W�*J�;0ER����M�)�P�����X�i2��s��b��U�.��K��1��AA��.V<��YM�l��e��[]y�����=c��>��u�xl���4��w��o����	B����T$7�aj���(8*ne�ːہ2��*��d}���阧n���ˑ������`}y_��-Zd*�Aṱ���X6@֖,�#s���ҤO$������;8D�#�B���]���rw#�/�q�h��-��^5��8&-cQ�J{�Ȓy��]*1���Փ1,2�Kj�̆_��-9nO���i%�Q�q��5�_��+��I�WAu
���]�cr�����ҏ'��=3�m�.z�8����\Y*�H%�<�(��c�\X�g������ �4�b���:�֊in�c{���>'��(�+��Y��X��ul�0<�!TGQ�ڄ��)��Au2@�&b;���|2_Y8�u~uQ <��+��h�~�,����[D��w�y���4YB���,���X�#�b�0ӭ�#��a�ET��rU4t�Z�'�S��ϲ���H�+7 ^T	�,�a�@�C��c�t^Q��9��3ѽ�"��`M�']�� �1c�1U��k���C �.w=��|:�������k�������Sb�x.�D�f��� :�gW\R畲(m͍!���e�Z���%�\{-�5 �ģ�x,���s?z���Hw���^Yۋ�ڪh����D����/���܇���XWL�t�t￯&�d���� 3���n����W̝��Z�rx��8�J���$f��x�T�{�Q3���k���g��?|���XM���K����OS�+�H�=Θ��,��V�\i�t��7����=���Z�W�O���}T7�����~Ee��$��F�����a��߬�:2�A�Ï�B��J��!E�7\
:c��0�
��r�	BHn��2�W�6�]3�Gq�ݡZ�b�Z;]�<�U��d��%{h�˅J�(�l�O�~1ѹg@}�4Ҝ���3_��J<9�l�� <�hA��S�=w:��p�j��G�8��jj�Wci��p_�&�E�8$�r}X-�qa�L�'�7A�����S�خ��1�].%CC�������6�����O�U��y�{�V6@���g�e�K�`���`��G�<��Wh�Y���`U.��+s0z+����~�����z5>��C���)��6��4[$Ħ-�t3W��ܻ:�v��Z����<�Ib��?�W*{�O����ݵ"ѵ�bTE�9�E>zR�D���N����j�ꘝڐl�[�Gs{��E�=>��f`X��`C�!!V�T���M�r��^p�S�����1:�?�/��^C���.;�nh����:{+�U�+��+x�[Tf2��3����`K�������[���u��&�J��:�r�@�f�ҙH6��0���8���ퟤ��V^s��3���rG����1q�<џB�d^��øQ<�9�в���f2E�X��fC�:m�=��� ����1vr�T7QJ����"�l��Q��s��C��g�×��hC�{#�i��=�����8'@DaP04Ǝ/�K�S_%�Ȟ = L�!�/����yO9��,.NNi�s�Zk,�%�ؼs��s��a�T�=;��}��&�mF�[�8�M&�Oo*�f'>���A 5�P�,��dSi�v�>��30��ތ���}�pr� �}�יm����T�`�dbG�kۃ���z��lD��32��v�G����<u��\�xeK~V��Y��d�1oJ]}&��*��!��*)z�uv�ъ.��:�=��M�����4�x�����1v���T^y����8��LV�mB���Z��RO4��i7��#��~�^�7�ۛ�V�Gm��!����o���K��3X��[��g;nM�r\@��U��e	�K�d�҅���9*4��7�RaY>�)�l�\a�f\�������-b�):�V|z��*��+�_�#	Q0,��^�E�*CF��#�����a+��/�'v�A���ob׉*���
��"	@�aVC�q>��G"4�~dm�Z"��jq9��>v��U�����}�R��H�V����,�Ġ\� �,o�C��%�P.e;��`����(�#�+�U�
`���������~Pc�,JK=�-�{p���x�X>�_3-k�`K�&��jj/M�d�s}�����,�8XI};�a8��?j��ނK0g��@��ޣ�'�B���>b5��:�Y_�#稓䲈5˻��E��u�:
�1&;�1)�廛9��ںr �n9)�Wa�bq���<CTN�wZy֍���9�>*?�D�A�q��3g�J���z�\��Q	� h�y�4t�s�%�@��Ko��D�F��y���s�=��N*,=�VHH�=�UiIEI7��#��2���$$�"%���	P���ܯ�ڡ����(�OEi�Sn��(;�Z�)'�.�{���_��xV�t>���>dx%����t����D ݊mb�Y�1a@Rl'GV��8a�tݫ��"�Z�m������ƪτW�LE���r����Qs��W�9�$4sȤ-i臛E4v���B��x:�P��1*^����#I���.��=�5�YR�0I�Ѣ��eα5�q`����\��LHĠ�
Z�c�m�]��������H�Qz��n��9�ͱ�Ep�Q��W�A�#��oA,�Y�c\P�&j�Է��co2���8��埦o�撫R�S��o�	h�7�]��j!M\�P�M���(�N�sƉ��Ќ�Nm.��垌���>&��2�nB��Ld��UP�EOD�I	��|����a��Pգ�����*�r��/�AO5x�;l'�mmZ�º��ˆf`�->j����6�M���-X�&�vq�_�ԏ'�4������&�O�q�[���X��{5�û�Y�N��cFU�Ǒ)n���ƍ��2WU{�͚~$�'������*om����2{��1ȇ�KO��&
S;�d@��{���6�֖q|B=y(� �g<�ι���c���Ũ#��	8�~@}�?�nie�wv��Ϊ����>y�dN:v�P���r���t%~�����^��p�����t�2�����4=@e��/�M���!�jZ��nZ����DU�V�8l"A<Xg��oTK��N_J����(�3;P���vG�8}F�6-E4�&�h��ұ4W�.��f������b" 4�r�JOH����YX(6�9�L蠊w=�}��bD��A��a�4F?�Q�b'�O���TåFU���5�
/Z9�	Z����W:	Vu��O,�Pp���a��Nw|�@��.p����Ļ� �~��]	�.�wF�$��Th���U�B�|�a-����4M�.� ��c1����R7l�	b�25�?���1]��ry��o,��ɟ�Ѐ+7"y�ʦ�V`�?�򵊽�i/��f1����r�w(��1䙤�Y6T���|��ű�
�5�9VUgk�;/�V������~f��"�Q��2��澺)(2���8�yfu@-�|�0|��L����үG&�9����\�����Q�ڿ����z[���e�v�{�;ä��oĸD�6J�!�0��BX>q�^O�M0�5r�@��{��WX��Zb��`�f+lx�Y�w�-!=Ő��Y�s�_Ž��4��GKB�MX|͆�\��ߗ�U�����z�`���ҳ�v�st�c�鍒��� zu�e����ߨ�Z���0%;�IN9�"Д-n]S�'5 yبj����T&&��n�ꨭ��&bT?��J�W�Q� �_U�o�&�)���t���Τ�U}�A��N~,�菞�,����ۘ.^�[f��{E�n۠��>f�k�B(P�;���t�RXP
��g����$���}�p��a1u6�ҽ3� ���I<Y����VS"��._r��)�������~�UPrǖ$�DS
���OWϜ:\30�t�1��~�ӷ��nEץ?©-`�8���}È��+�k��L0#�"�3`Ub��{��Ϫ��22_܋��xX��wV�C���EP���Q0F�Dh/H8O��#F�D�$Ŭ�aU���,6��d�3��ѕ�/�����v(����2��R�ф >��NӶ�q�
Uޘ��Ч�o~�Z$�9�q%��qnn���@�*yu@*;>Ɍ��#V�����EI��&VMͭ'���m��5���#2�{�ߒ�&���]���^���i��� h;æ���S���Jč��ڨ�<f@�?=�&8��QG=
7ў9Z�2�2-����x-�?m��i�v�\I��������U���@��������"56$0*�ĂG\��wu���U=�r��xW�1�f`�==;���^�$FO��P$�c�v�9Y&'Q��&�d4V�
ê��m������.�'.s��[:�s ���7Z~�eI:F�z�vML� DG�o
��j[L��2�׾C� ډ��b��ܔ@���Of�T�@6@��c�/k�nfu�|c$���������Q�ٞ���v<�=����7x�\�)-�G�Ķ�����x��|�nd�}E
�J=��I�ro:���Z�W_��m M#0M(�o}�n�$�0�q��g��R&Мn2��W9�n�!����n�(��e�����d��;�Ba ��a=̦~��4y_O�`���^`N� ܓ��i`�b�kM!���Օ�[�F����8w�H)��9�)u��:��Ւ�$�q�H��-�yGGԿc�Te��hٲʕ�/�*%^7���x�7�ց2���f�|�u~1z��d/�I��Q��f'���e\��F�s�=]!�:0��h�sP#��ʴ��3 c���|��2�C�E#�����>�8�L|U�ۦ��U�7+D��������h�w���|uUC��Z�CGl�H�ѫ
S�c�ȼ����5�hI(��)/ז3i碂\'���%��P��.�1���!�غ���z�O�y��n��+��lF0�wțABa��}'с{���E�E��rfE�Ug���pU���ܞ��h�A������f� a:='���G�n��o�p���@���U�����7�ztdk�nZ%��t�j˴��n8T�oeX�)��)���l.�iJSX�c��_�P^���K��zq5�^�bY���_VH`5��	�eis����VF��R-g�M��b�/��0󍃩�(�g�#g�U���G�^9�1�a/(�_�I_��#b֍.�V��G����B^��)��M!����&�~���D�=3��7���1�CU�o_��<La�Y
�'ӌ8�b^�@�C��<QK��vF��ű��L�����W����aI��2!y�{m�`�kx����QTJ��
�����TK�@��Q[|�ʟ�r1�Ĺ�3cg70�5��9�oЮ�n��,|��޼�=�e�χ��@��gh��(�XY�e-{�%h�p���حã.�P&E�l5'zI�:6�0�|.��g�z)�H^�D#$���b��x���uU����ZS�3���eu=ɍ+$bs�j�9�c\�����~��XljZ��@Yt�B'��� R'V"_8k��3�EK�d��9&B �%����&iú]ـ�GQ#��*۾��b�_���S�T�ں��~��šݗ�qxf���a�Xٓ>�a"еR��ڙ����x���uk�-W�"V, )$2k��_a���-ڍ�l��LsEЕ
E�� �U+�k[��t)�n�>W(^Vc���tPn{�\��d�7k�"x�'�2s:�W�LIvur��F�
��'�)��eHd�"��"����/� fN�m���!8����f��
"�Ի.�yZ�c~9|u����O�wrmtMY��Ge�r�]�I��.�L�N7�fS�ə��0{1E|%�%��'W"����t�*�ՠUH$���kb`��R����á�>������͉~���KQ5'�TL/�6��m���8��lH>q[�Qh�1�f��E�?�[����av�e��U']�^�r엋]�w<�iZ�=M.P�� [�Z�8E�z!5�7�^�>���u�;��z�⑸쟜������y5�Đ����	&dnҶ��`"`�E�Q�!HR�8�IYz;��?� bQ�9o�EG���6�+��be��IS/�iZX�J��UP�y7G��W���)8_�`~���y����Ov�.C8�l �������w>�������Q�b��)�Pp�Tm�5t�\h��դ��~�����v= ���v�̼�E�ikk��it�@mőP������Q�Zr/�εv�?�� =c�Og5 ��6�'a)����S�ڃi�yL0��l-&��y����gIh�Jip)f& �|c]�<�)�������q�������_X�9��90+�|�F��|�Az)�\/��ʹ�w��<�����׏�Ԕ���؜j���ā�k'���2v<��GT��g�}S���VF��^IK�yQ����(�i�	���;aG���ee�dJ���؀]hD�-6�#������ÜH���A��3�T�:U�-�i���W��9���[QA^�s?@���[%�s�|;��F�4:����~(�������tq ����H���_� ��i�/͙�$P��įX�d{���ˍ}��]�DKt��0�8��^��τ�Z�/�RG|�D�n�a��y;f&�@H��4=)��B�~�ȳ���
��]�>%By�L�דO�hx��g�:V��W��QVD4��`lw����(���o@*�c�T�����#���ZE��)�Q���nT&��f�����d7��4Up3�"k�r ��2����|m��,i�^ϱ����?�^	V�J��(ي ��~ږ��,���І���{�)��	�����N�n������A7U�-o�W(Z��Ϳ���๯S7OXF�u/'UC��,)~5܅
Z�76��:qa3���H�s��iEY�t��U��Ʃa6�͔_~i��h�# C�YV���r4�:���Q���b�}s�l��,,R@�%���NMnʉ�J/ny���	�v�b`���7:����<	@E��C�K��B�c�C+��	��sSO��E8��ebp��Ò��:�sO��@�@��I�`ӌ=m�O�Fh��p�f��{]W.g��,�`<�7Ī��ZN�k�����8tp)�|b&��{)� ���BK�@�3�VZ|�j��ܻ�(��FwF��M���,�-Qr�[Rl^Mt[!��127'r�9�J�&����/tD-X�{��R0�&�6�`�Rנ#QpƬ6@�G_��i:�(!��>Hp|����<Q`���4݈���=�o��Ů�����U]o^��.y+�O�Q����d��S��7' ~�~���~��Ĺ�MϞW.1V@��lRA{�P4D���GM!�Vq���n���Jc��X�"|D?��O�9��/	(��N�<o_��q���Pߋ3�\$[��>^�l���7�������P��w�Q�h�ݘ���)�w��i�E�)L4��B|�׶����W�6������-�Q��5�Z�����j@���N��vm�J����y�7>��h"s����o�!���,�o��7��H�j����gy��(>%��C�d�ƻ,)� ^���TN��#�8�ZǽԤY���n��Ǭ9��V����ȋ�M_7�I]�JI^�L�VEx��a5# �[���NPډ6����k����gsX6C��*k�U<�u��c����S�\�j���ӄ�6 _}1�����JW���a��I@��i��)s\�����ڪ�BM:(~:Ѩ��*��[��h���'3�z��3�\�ԻIxc���$�����Lǩ�^2����P�Z��Pr�	��N~�XEkӷ�<+��Ug�j}IO�r��9��{�	{~��G4j��u�p�̿0Ӈ��!��z�K���wķ��LA	��7�"�K�<�Js�� l����ۭx%4�V�HG�`��mu$�'H����5�͈�x��V�2��(���ü���sPP�a"ִ���*�Π�%�����%m�(YP���M���,�	?��_&�j�sᖞ�=���
E�&�������τ���v��|rK��1,�0�E���Ij�ub����X��L<�WTy�<�иd
( ��N�-:����L�p�yTnF�(��������:�ǋڷ��|X��ٺ�|*!���/m�#�"�A�k ]cw���F;P�\�r�跗'�`�_�w<��������&z��9��Qǅ���_��Z�%�V�A��G��Ϭ�G��XG׎9Y�l!������e/z���q5k����	)ᶁq�m�I��i^!������!�73����ά�-`c���z������4N!�N�A������-z�A٘���\c���*e�v.no����VF�-[݅`�6�Ù�S���p�uR��n�N��-��3K�"wQ����q~��d2mř�:W�L���Iݯ�k���������M�&����v[�\��΃߹�-�7u��)[�`9��[������^�e�3���N~q�:BJ�����Y:�w�ߊ�4�ڸ�*3=2���8�W��۝���3R%����q^�i���)	����/(/�/�qX��]�����z��1f��.K0sr85�'��q(W<����O\��p)(^v�� ��+#�� 1�-$a�v�Gur������e8�c�%e��Y����o��R	��6%qR�X�^�z�F�xv&)�|49�Ǹq�U�N��"�迹.�.�B)��ݸ�ZB;�B�Q�$f����06���D�@%�-l�5�m��H���9�'9�E��t?c����d�֍yVg$��ZnJ�����ի�!�����eW���c��ұ�Ul�D!�ҙ�ΡP�.����ݪ�'�
�.G�LL��V�"T�)��j�߲K�S��5�W���͗�z�{����v%�ѓ4:�2��؞�Ӹ�)	��z�t]|!�ߩ��h*����*iި��#|}:a�Sˡ�Ɛ�/۠��c��%ɉ��"
�c�aP�>	e�%%_B7�G�孞�\e0țS�QG�&�9l�A���9B�"!�rT'1�ڃsɆ�GK�g&g~P[ɈX���pC)͎,��X7@s�M~ª�� �!�dϔ�����8MН��D?�=�7�Y��jn��_�a������9���9�+;ϡV����>`�y&p=�>���w�Ұ�#!�0R�k+�M�XҲ���vB�)IyDhV��vt���g����\��^�� ���� �4$cb辽���~,��QЈf��wӉ=����&g9K+������$#-���I�do�=�A��.0���K�B`iϠwT���zD�{�wh�#�5�"ŧL�D����E��'vhK����IBN��KF�FhƁ�;u��b:�43;�:Mݎ)��b r�z��mWn��P�EM!�NdDV�{�C�	͆���S��|7�O����܆K�_o��7?�|7��L�'��Ug�É�-|��+B+��'G��������oo�����&k0 �a�~`s<�����S/�K�2B����(/@���E��f�>f�WL�*�}�:=}v���bK��#�R�G/�3r20�tE*0 ���Ř	Y�&I���:�ټ ��^n�_�,������o'��o�̩$rrJ�T��0����vr �ycA�dX|c;�	�jI�@�{A���po�Ɓ�^�\�09b�Q
3t�����E��� _ �U@�c�%�)�#r�m	��UE�AH��h"�8��7�&��T6V{�����vl^�a���s�^� .�m���[�G��~�K��8$���)���N�ȟ�h�!9b����1�(�,���a$����2�`�"�Rt2��Q9k�c4�W��ʝ�uD���w�/��g�#Ƥ�xu�Z_���MS�f�c�H�.��c؏�ְpc�
�Dz�����	��	ⵂla�[�|�ua��[�Z��!��*/�4S�D�F�ן�K��p*�08���4�� �/ք:����a�a�wZkٲ�5��MbT��n)�Ⱦ< �4��zEt��h�f��,t�b���Fy���,`a�@oɔ&E��Zt�|=>Y�)�Pgb��_��WdM�Ld�e�F���m�6"0q�Of��#�2�8�%[-�W��D��h���j7��ѻE���=���8"CF29~�X�T��.F��|�v�h�=S�y-��Ea=Q��*�������窠��Y���U��>aB@\�~,7<�����X��T�� ��H��S/������#�2��b���S/��zO?by����ߊ�2@�F�)n�f�	,j��b��y�����_A[��L�=����q+a>2��|��L�80<�Ԛ"�W���ya���������N3�Y]�+cO�WS������2�~�!;��7\��ן
��p��(_�Ç�!k�{�	ݷ��5����n��gd!����ΣHT��t">f�G�w��=�蕙�^������������:�/Bz�ߊ҃�/Ź�
��ow����d�qi;p7ޏ(�˱>��)qH��j�1g��AJH�8[ְ��P)0L�{�l���a;=#O���Y�R�XO@�I:�9f1�}���_��
�.Q���X�?��F�����:�ӘM~ҥ��P"q��`��`����y�2�]�m���Ć������/eX�)�邲޺h�C/�U���^��Ї_�q=R{N?݋�D���o 85����p��w�֝k�1:�3opF۲����F"n�Ӊ85�|��[j��X�~su��^���Ϙ���ts�T�f@�})�jDc�T>��ux���H��M��8�ڎyLHf�1k�8�Z�S���g�. �}r�U���j����iɽ,"�|�ض�EG����լ?��pȴG(��~yA�aMG٫��I�����?NV��Y$���o.��D���l�[����J|O��y�$�fu�܉j�����ET�
g����⎧�il�8��8X��-cz�ǹD�W�A�W%�s�ݥ�H�%�C$ԜXo�^5��&P���!Nu��m^��2�19U����n%�_L������OQ6�>x���~Q�cl��u2��n�f��;k/H����[�R�{���[��m�t����I���4�R�F��o��⺥(��b�y;P�G�v�\��"�=o��q^L٠i�r/OO௵�2�TnQ�uX��*R� [�O���NB�Y,t��D(k�{��<�$��贿B����9�-�2��J�%Ҿ�;a��rL}3���G\�p���*x�΂�J ;܅o���'���磜�����v�1y��u芹5Y�lu�mXqb~5~V���b��VG�F�
4�p�����{�$xo8�t�浤�|��*}��KDK�n1v.4c����NR�-��	'�dw��#�GNJ��VYq���_WO�)&*�t��3�0h<?쪭��~�펥
6,�N^v���rfI�UBF���Z�+�	��%QH�y�p����"��W����_�C��[�U ��j�w��:ʖ�L�W�RT��m�tj�Y�
�q�n
�E���[(/,���BP�H�1iN��:���In2tL�k˱wK^��C�A�8�i��D}�]�.����:IL�Pc�Ӕq8\u��l��_�C��v@�C���9�w�y���6fcL=X��ǉ{�4�0�^���('��U�kV�<�K�q�Kh�����c�\�r�{p��]���S�h}�?�Rhk;���o]D�N{��F��˫��	��u�4;߆���!�[�U��<;�(�Kp���Na���#t�gT�⪡����|�1�i��	2!q�Cy �:�q��U_&S1�O`��J�&)�S�ȯ*�����&�R$�|Rd���� oG�C��p;��,
����}��z��=�7��P�ضZ7������p�_�1��n�`0�"w0�a�{�)t(?�Z��������Sd��4d�k3-p���p#~*>W�s����,����R�� �¿��䣚H_��;jo���
���n�!"�_�I?��ͭ��qؕ�07��:F6�Ф�;`�LO
��}���ya��7ɼɲ��_�~�"6��*C$������L���RF��k9E�da�^�	�O�G���O_���
H�a�Ht���ze��^��~�o�	&=�������n�QS��줌�(�ݘ�rK�{��x(h�]�w�Ij|�j)���׵w���D��A��س;��b��Ǯ���(�p&�Ϭ����2���6��P"�P��Y�ДT�}X�ؠ(18Zy2���0*b�|ՇHD$<.l=�Ġ������#��I��'�'��\���L�,T��Q.�%�p��Ml�߮j;�����V�<s�nL���F���K��J� ��z�ߞ�%�3"rWƋcPu�O
������h|aS3;0���X����^��+�S��W�/���Gd`D�L%�vPL�Be�����t �D��%�G��_(�L��!B�P*c>�g1P{B���b,�n[��d��km���4�~���'���J!]zw�nbqu{.�XF)��tUÛ�w�,[g&�(4�q'	�;���9����=�Žf� ��~���5���J��h�F���q�Zź��NUȗ���|�"�u,�tP:s�f�hFm�Dw����1�#!��C�v�5ۭA�T�Y���&�H��g��rO�y��^M׺)ˋp��/�6[���⸘P�5����L-F��v`��y��$���;篱#啪X�I�0T���}�2YV��r�N���T\0�WGLl6���v��Z�u�T9�Ӕ�J��� mh7Xm;Ldwp��ǎ�Qӏ��QOu_�Q����^����|�f�@ �/��h3:��ۣ$'�c��[�r8�(��*k3�v"ɕ�}B�2��Z��u		f�8D��v]�k�ˑ�cy_����d{)���r�2H��+�ڌ�l>���p�TL�n>@��R$s�D5��K��lˉ�1��y�̪������q�k@A2#�F��t�0���>�7j2/S1��?Q�AK���t�.�=��f�&�U��?�yJ&�Q&����iք������*��_���(�
��Ծ���ܥ?z��i�1_:�qٮ���]��;��d(E�5d�����Q�b�ua������ j;>�0�{3E�^�&|�uI8OS`q�4[`%�L@X�9�C)��1���dZiu/�9�1�rA�J��j�*IK[i^�8�f�q�9���v�C@�	�o�#�D�!�5�����(o��~.Mj2پ �����o/*����U+q�͝�)h�6g� �O�*�^
8�~����L� <6�cي�y�NN|��H�ǆ�v��+�iG�\#ߟ�C��Z��%;�m=�K���D�bJ۟�tc`\�ߔB��	]���2;���m�֚���xE�N�T�����F�4
8�G՜ Ys�u-F�r��g���Q[H�	����(D���&��j�c@��s�ET�K�j揻}!�B>im���r>��櫶লZ{_���C�#=	:C%3���-�S����]�}��2�����(4����i��5�v�ȏpXU ����\�7:�N�9c�x���3�9�=�s����X{�����2��U�GT��z��5��f�(	������C����Og�_�h1�
,®b�rH�S�(�<�d~��8�M\ ���̴���1��W6�E�ā9�(�i���\O4|嗱��𢓴h�	�-Q;����h�f�z	M3WyK'��Y%�A�q�@�i]K����n�j%k
D�YH~(΁�\ZcvҰL��)u��]Og�g뷨1^^��cP�D3a�������a�_6j��I��t RT$t��b޹(Q`�E��|�,Sʓ�del��;A������&�����f�!k��H���Z�1j�B)�mĥ5
(���WT�t�%-�σ;��3�d���D���l��j�A���4�y�n����5V�dS�)-�~��~Ǻ�p�q��ǩaP~(1Q�"3|N#(�b8ph:K�`��<�<]�����2�-���W��0{�xJ�m<ݩ���e^D����D��?k=�7�oi�,4��VF�3ҼSu�o<���̀��茇&�x���;6BO_�k}���N����R���o*�瞏U�35x���X�5����O�$)�;hS��<>Y�)~..�޶��^��uyY���F[`�y߃k�]����(���A��3`;��%؄��y�8,~d��`���^�``�ɺ�M��mjD���*r�w�ui�ga)��l�4�ữ����v��hж]��o-`T���^P7�CŖ����q���T��D��������iq!����o�z�jM���	��?�w���_�C�c��"=�Q�5����+Q�0��FF���N�w��:��RO0�r���I�F&���*8��UC�r`�VU���HG����˅��&ƅ�U�֡(��
+��5獩��F�Jd�������h����(_o��%<=�Y�܄�6�1b'9��dk��w�]�����0�$�+�9��S�U��`�W}�ɖ>TH� ���_�t�D���Ȯ~$���N�@�	0�[����?(׶�y_x���ya$��tk'��ޱ�T
����2�E������rU� fM)E���.� �Z�%�w�m��AS���F..!��qC�<DBv&UF5#�ěs��y���q�e9?�2b�S��`�H��[N��SE�"��mR�QP��e'W.�2v�P�0p1��&o���s�8�����=9�Q��dS��N2�� X�lb'�Փ؎C�4���˿�+( ��1g��h�nՑ�|]�:�����9M)��`97O�i{A;�{�䜐�r���p��<�er';t]���vO�� 5p��s����*w���9���� �Jþ�m.h����ۛ�h�!����D�$����E����$�M�P�!�h���Goi~*{��ږK ku����� �����f������nf��,����^��S�����:�����L%G/鞥ɢqI;��{��*I--�`ͻ����~��(-�D�M���˻�9����?7zd��mk0�����UQ��:9Hm̑��JV[M����p���I��H��]j%=

��
����#�®�P~T�T5��>��8Y؃f�=⌥�(��?���0��r;����^N��Mg�n&c9/K��c؝�3�@n~m\�1�����(�P� P�`c�!��Xlu엗jf��<�L���:�WG�� b�׃ ̓ޟ�"�]�{����S
�qp�U���[r��;ԝ��OV�������``�~1�(�����i��^r��I�ɝ]�f[�?yD΀��ps���ԃ]��OH{�C�}}�>��,u�NP��ŃI�E/�Cm�0x��̵#'�S��-Ư�����z9W��sC�A"p�2qi��`�)������yz}��z�q��������+��#3�H��|�?��+�Dg<\�rh^1�rd��G�#Q��ּF��<��z��+T���+��GW�p��f�n�Tu�*�B���[DFx�̘�4+n� ���|��k�>[w��[N���v�ط�Z��aJ����S���u�>T�m�; ���5�E�S���7=[7$��ŉ�^��h�����=s�Wi�S��x[u�M��Қ�����@�_�`�����9���w�Y#��p�vh�������k1Eޏ�K�Z�,K�ݤ�H�r##A�!e���0e��i��f��9�`����]2�,ĉ$�ax�0ȯ?N�<4���{SA+`_�����	g3\����;��R��6�z�f�'t��G�%��0��c2�{�Ѷ����u�E�q% +!�f�z^p]��f0�#�d(r2�
+�ϑ\�
���ϻ�n<�3H_��:,ʎ����K�H�d��ĉ4�� [+�����J{�-4$sZ=@9w�Kk���w��
4�Z s����A�����}�b������S�b孛�is�5���6?���I��=�ӋN]�:"�e������)�Z�\r	�/��0���yTVk}'��ƎGlmYY�^�ju���A�v� ���4[����#>@�{�ع`r�����k��.t����R�ѸIė> )<��b���8}=��Q܈G���~���P��@�C�? [���tD�]L:���B�^+���
�Z[>��G���)�IjD�2_׏JC������V�QD����L�����ܨ��0B��+��� ���⁡���S�I ϲ��B��)�
Jl�a=K���x|�#�������8.�d,@W�}�e/,�h�ʂ78Lr�\�0	5�b��˼*8Ģ��@��7!c��-9Fޓd������_zS|�7�����23c^�9�4y?-A���rJw�ۈ����MI:DnAV�u��n�WI@d.�5�e�6�I'�T�F2��	��D���|<��@9��	soC3D`��Z��ڂ>�R��ym�2+��0�7��b!�Q���G�5�a>b��)E�ުGnk���ո�T�v^�P.�uo�n�<��R��@�:v?��>�庭r��8���4!H���X��ip��J��qU��ߤ�@��%K�
��h�+��H��^a������)cn��)M	A8�b3��;ʭ1�a�����"YJQG�<�s=��9�Gk|Cn[t�����`3B(���X9U��z�w8vgW�$��=�>�}�{��*h߀,f�Q�:���"(c���{�?�\7��F�ul�rK�R�������,I��{��8�a�R3A��]o��YbW�S��r؛>0��"�]��mS�0YDJ7�� cys�=��Õ��$d�x�߻XSmn�u�T��e�u�V�����"�y�Sv����`o��}�Ą�1�#QMఇ�����W���4�Y���R��������M|fY�h�ɻ�~{Җ���.\"�>�6�$τ�t���͗�B"s?�\t�D�&J�9~��AלFI ��a��2�8������(r�,%��j+�������/���FdX�e��ў�]�Jo'�fZ�@z1�k�c��M_�EN��� g�`��� ��၂|�`ʍ��Tg<%ȗ��,���"�B��ŏ����5�����ҵ$��e��l�K��#�]OH�E��f��M�/�Uڗ>ߓ�|`�<��U��0k�z��Y�5��B���x�K~u3����S�����?���S��^"���E'l�����dg`�e��E(�^�[ A� ߾����맆Gn�Ȝ�R��6�/�dS��Ew��amq�����T�: kFJ���h�T��%�y�Ư4n�v�05)�)Av��[�<��a���V󹳩4~:x�T�g������L�@ѣB�W
��@U�@�Qf#"���f��L����7=�'�0d�q1�2'~,�g��z��&_����5_�~g�R	x�q^�7%�4G�����>�rM ��.Ed"��&�iO�EqL23��ѓ�J�[T��&v�aą^��p�aEi0' �1t�#W���o�����4W�{�䱔���0_�2i�Q>ƛ��Qn��yUG�^#�ٕ0���2?�2Io^#���YH���GGW�e_�n���ʅ�M�"镳�w$�m���e#nhS����������buXs�Lp�Y�=�]а�����kl�Dߔ�wT�4�����QP=���?l�c��V�q��������Y�	$l<g�x�o6~��N�Γ�m��� �K�Cb�3�T~Nl��W�X���P�/EL�*�=2ZV$K����%+��jy�[~��RRI�F�f���s)+�}�G���]���VT��]d�d9��x�#�Dj����J
�|}c�Tɏ���lɵ_��t����vW�A�����Pl25d��)d���z{ȷ��8��҅�����=�\�~�9����:���o��-��ӀD7�ܘ��
�F �5
��X��{��:W:dUv��K�a2� ��vC?��\$�i�N�k!�޹�f@�L��-�RۡQ��{���W���˵��;�J��.η���Yя���L3��P��k�UY4E�m'����Զ�&�u�4wkR�UÁ���j�1ߜ�Ow���-��E�r޺�����q�P�z�n��XNy	�&��j&M�����­h=б��rڪ��h�yH�[	��/1s�'8F�3kh�� LmsN����{��i+������)BKs�fO薈W�uq�vv�`ad�:�su:�qpU�،H� J������W�*����ؿ. �Auba8��̸Ă�t~1�?&i�ؓ��F�+��륥}�;�a��٣���
���L.C�aВK����X�6���"Np}<5�`�5q���Ť�k�w�d���!��q�փ�� J!��9Uh�~�̍����E^Sd�`�O�FL7�d%�f�� `�ot�?-�Kn�K;n)�x�웹;[	���ia� ���3���CnL�)�a�>�2B�쐘ԋ�w�)_'�\T��զ��P���h\�|�*
bh%n�׷ߴ�A�L�3��0�+�/�m���η�]7��(�Kϯ���Y��:�6���L�y�2��t��X��_��8�3|U��N�\�"�';���E���t&��j��W#�ņE���i�S6����]()\Mx��ۉ���G�І�ۣW�����D�hê3_�8p�
xE���9R�2�ˎ�)}�+���Yu����@Vz	�ͻ���/�9�9�P�:�%d ����Q��o핧%:��R�s�
��v1`�A�ɚ$;�i���
�Ac�b�֨]���ڼ�&�&1���qH�LT�{]2�ߐlf|���^
T�u�u!�K��@�O71�}}��s� <x*Q�UP0*n"G���'����B����6	D�����(ͳ�#-ΚΥ�!l���7��<=u'\ߏ��lui�&� ���I�>y�e�����e�~�f�aQϪ��z�J�a���^��:C� l#�)P����T�#��S$|���~U=3R�^ �O쬇�G���X�h��<�`�=� ț�ug/5���z�́����F��p��"[5��fоT�-m~����S��R�sxd��Nq����p��n
��p�N���j�)M�/�p�%,(�ܑcI q�2�z�u�����!�ۆҒ�F3�a$�tK�h�'@��i�s�Z6�r"�3@��(�e�PG�y=�ƞ$�^��ή��a���pZ�Mk�;fꩪ����J,!���~�Ky�.DC2��~7���`Т�7�Lg[PH��F����!�)!�ĥ�9&�1�@b�=b�]zv�խ�ea~1��4�����ב_r��+�p��з ��k2�p>�"� l�а�x���y�o~|룯���jsL�<C�~&X۠�_�5�28�N+�1�<��QS���<��mI�z+`!�tN��#u�?��+��	��T�h9/�;����M`�<w�ωB��?��ba�d.h����W�_��rp�b�<-8�xP�2*ݤPl�R�[T5��=��5�Ӈj���2:M�s����)�~��Q��9κ�ԴSl;� H+���=��evm�
�=(��W�M;r��W]�8�����/p�<N�If������i��3���es6�z��f]p��L@�٠�}�B˷��O�K�x��ll�Yң}�v6��>_"���0��[���/��?�S�T��?x�������WlEӍd�"����sB*�ӷދT�}�v��=̦�� �;$*��۬(Y�boxy��]֘�j0���.�C~���6����]kPa�3�D���I���z�2�8{�q�����u0�˶[ޕ���8A9�J<�4Ú�o)4��l���c� G��v�uķ�"�7Dܑ�h�����ښg�SDo(�@cy��{�6l���h�!���{	},�E�{.�5�x�yWH���K<6�� j*����p_��j��&��01�U�R>�,��]|0�X����P�:0�??�݄��sM�;�o�s�6����� ��qi50-r���1G��{G�9^m*�!������甠hf��7y�01��yW̚t�"�ђ�<V�o���V"�x;���:H"��TW�����i*�z�������{Z���K�����w��D�V��#�IԖm:0�3�Ğ_�k�s�Hk��=�&�5�}�h�IWGVD� �W@���j��3�����n}�C3������\{�7B~R!�3@��	�ҁ9�	R6��E$t	�x�~S���	.�a~��ٿWK*�}L;���JV� �����h�CT���F8R���)d�6U}~L+��ۂsO˥��(�a;ft�>��q��VѮ�?Գ!�{�Q�CD��5r`�F�=�O���n6t����2�\V�U���$����l�3J�C��|/�&�!@DꌖQ�ۚ?�6穇&�C���Wk����U�%� Mq0Q��Rx�����-�DdT�A���R�3������ԚZ�2�$���K̙�~P�ǹ��U�ӈ_e+�k|"ٮ{�z��o�p]��@&ɴ!N3�J�1��_��L�OdM{�&�'o�cUNʨx�b>d$׀�-��v'���0k69!�[z�1��%i��9F�ہ�`��\�	����ӰF8gI$�]��}M{#�==p.O��-d�����=�J�0���=Y�{�����wb=�Sb�:�pʽ�$A3(���,N��>C@v��Ū�)�w���E�Q,�hK/g�L�+��O�I�J��h�G�T!����gL��0���t!�>,kϏK\�>yC�����{R{�U5��+�3�kq-_!�ܛ{@/w�'����ᓼ�,����gѫ�j��e�_��y٥O���9�;X�jbց��Qh����T�2� ��������ڈD@ΰ�`��?���2&}(����6�:����3˴�f)�+ڔ�$���H�9� /�����H�v�ޖr����=�p��l-��*�+?�������n��|� >�~)b�5�x�Sgz����sY���V��w�| 	<�<�p��t	�3>c�DH�������7Y��y�w�(_�Im��;52�#u�J�Ͼ�t�%_�� �������b7�^��k׉g�Ϸ��r(���6��Qsʹ����vM���.�S��ǲbċEa��ф����"�T�e%�.VSbKC°y���-�� %��j}�T3��U�1��ykqw�UǶͷl�j�4����cg}se��|k�e���qvf�T�������o��Jk�P���Hx�|�M��"���.�!%��0�����ݷ	w'*$5ę�Pd�b�H�PA8�1��u(�� �=�c�IQr�S�è�)���J�6Qxd�Pot׼&k����%�b��|Z�Y�����ˣ��z-d�P�\�kS�o��>U҂�S�#���oD�+9hd�Ee���?�U(\:�9@�-.-�"���,�Wz���k���|���V@2BuP$�/��c��9T=�Ǽ��J4z��e ��Ó��Җ�����@�c�&�6I
N�v�{�����r��?�� /Gr����ww�,6�i���>@�@�o-J��{��S��9�9���mϬ����mI�����1�����I������f(c1?�rK4��'~B� E{�%hWPƐ���ѝWV�1`���t#��<e��3�5�b�1���x���?#:딒��eum����*���ri��}��}��푏ޝV}�9�Qb6FohI8#� �䊲�	N�eG�X������;�'�i����iUs�6�R������̎����joWu5�0�q'��|P@{�)��qI�W�Q�"}�Y\s/c��d�6���(�b�� ��b���T����5I�)������<@���Qfb2 oPǞ�$F=��yO���&7����LpvN�G4�h��M��8�O+����O���)��r�ȣ�3H(� ��y��� M��Or:.Ҫ�֟�1P	qs\�p�����!�!���8`��OlM6w�!����������l��= "��n��%QOM���B
�4��t��;5giG�^�ɸu�.��W�8k�xi�>��b5���'�q�9���,���>c�v]�a7! �0��:��T�pP�%�����:�#��#����:�n����y\X�4#j��\R�~f����\j�IW"�d�&����N��
�b�Ց��e:^�(����Ji��H �-iѯ�o�̰�.�M:�# .�����V�-��d5�l�{ה�R}�8`��m��_gkcu�Ƌ��X��W�G���Á$-��6���<n�Tc�aO��q�7�]��˻ؖSV�ר��?TҊ}���ƅ^0q��arN{�f���Љj������p�x�m`��$�蘎�S��8��kۋ�<��զ�kM>���0DK��^��|. �^���'UsL���L-t�3��x�`��63v�l����ߕ>���n/f��v�SJ���2X�;�>��?��l�g�k4����L��h]�HK67��Z�hŗ���e?���)'���ZKbgX���֖V���K�=��c|��=Y.X�iJ�:��~(.c�R@�{Y�\��L��!����'�H|Q6�N`F=%@A�'�o%8�ȅ�ì* ���p�24��&=N�V�����Ұ�awD��4Sy���ot�Ȱ����I�
)l(�� �q�1/�=��m	�׊� }֤a�B�֑�{Uq}+��aH�u�/Y�4�)�~[����7Ja1��5q��9u�#�
"I�T��$�HR�#�\��(��ړʆ�A �P�
j�/"6$�O� ���.���P�P��{������:�2d�L㾷�_��J�����tCX{w�N��h��{6��]7�����R���_�������ZGu
�]O�x���
-;Y�b�7�O2���?֐h�E"ah<J�������荴�Ю>�x��`zQN�hغ��M��Y�A�� �оɄ%4�Xd���c{�I�L��g<�GZ����'��.�~����F˛e��8���Ul������jU��A�}�Z����>�t��|�*��(n7��~���1��g�^r�N�0,Z����+DS��,�p;I��BP������ɰx���(��L�(�\�}��mK��S�6>I������D$�ۅ-��� �v��>�ȳ��k�WH`95z���Ə�"��ǣ��`����̈́�Y�Y������y���t�`��]��#0u�ߊ�H���UvG��c̜Z6ΫhC���r�2V��
�Rd'�s�7�7&/@�C��,�u�Fh�X�-�
�'+�uې��C�v{�@]�,��tbD��)G�C�o&*JU�F��"R���ː����������-���F&�7��w;1���H��7�7ċyB6��/AB-@��R�y�H�S�Ps1Ly�$A;j
&�"T�̔Q���ҝ�m���+�Q��C�zM%d��2�H`4�wd���]lí`���ћ|Z���)SSl�����v�a�F7�Z=TED��7Ö���(d}��}��BG��~�(�r�f8��I�A�ňfV'/��\��^I�,��*o#�bc�̂��*�e�K�L-�5^��/O]�揵	�FU����<�f�� ��'[�_�Ͳ-��p7U���K�K /Yu��\5��=:4�����@c*���]5��v��!�O��DK��C��Xp\5򓋢���J�P�k��L���MN�z4�H�:�Yț�ȕz�����w��{٤�O!��S�7̶��4?��1.��J�ͫ�#��к�,=�����5ɵ-:[DG�!kxv�
�bn��[(�.�Τġ�F�E����$-���!�vZ5�`A����vȟ��A�L-�X�L���X�V�/��0)����?��A_=,��1�Ư8��}Y+h��2�N����)���4tɹ�S��[AN��"�Q �6�~鸑F܀7'������2��;���{x���=��3�!556����kZ���<�d|�2�	!$�����IR��ʆ��Q5�w%V��xRU|�ëQ%7��J�S�l��y����$�Y�2�n@�Mx�-{�_B+\�3�~�o��^E2Ym���gf����#�p ��8oV��0P�AP����{���+s���0��C����opjλ�6{�!��YY0���X��8�ߑ�дp&��2]R����&8f�*{7zI븯l�<�"h��{�vGn5z*%*��
��ZȭU����d�?��J]�XW�s<�otڐM�������Թ�B�)���i�p�l�wiﺯg�;O�� q��6�D���F�o���s�W9	�4��&����ZP��2c�hF����w���k��&�:s9�|qE�ܦc�eJK�y��| ����h�L◜��,�X�K:�5��F#-=4�_�FnV�%�^��R��E�[	T�z�R�S#Cj��d�N�J��������� �,V��s�ޑ�*,��2�q>�_,W��ay��W�^��V �´�c��B�M��H]e6����Ȓ������$!�L�KLO����YV��6�б�~�9����9Ν��i<��S�V���B:i�릘G��"\<-�������@r�p��	�kO�Al���Y��� Q9x�Es��Rr���I�#:3P
YNN�lJ�����*��6���09��d�^����sE�,���H�0��gس�*!��9�%�xL[c��!�����F�2�π�o�7�bSF�������vtj�*�'h���W��Ǜ0�ފ�.f��fa9���������$E͖��3�v�	�.�谟q{b��I�J=���Q��I�d�ze1p�M� �՗ɋ5�g���~m�
xd�Ź���, �x��\^��q/E����qo:J�{1��G�[�����B�t��ֽ������u�M�?@��"�����sR龌����o�[�\z�g9W��Fj\��Ť�v}��n��=�:=28��������]m�к�%��V���g�
�6hp(��"}R+`r��gG�2�Z�.w���)��ɳ~=$,�]?�Y��&Du;k���QZ������O�����'bV�Ѧ���g�����Z�q�J��A�%����9���Z��-ߘ}y0<	�].�0�%"@�%�5f�!P����g:˗�.85��}�b����NDsa�%@��B��,�ݢ	�㗍�4��]���^C�qaMA[�N��͖-SO��O��*�� R�F+��{ʓj�d�~Vځﾘ+t�یo=y��aq`������Yt�B��	x$�}�N��\����&�PuP��D>��ݝ��3��0eDAj����JN��S�^C?NГ�<:�c�6�T`�Y�zb~M-��7p�JՃR!rP���d��ش!u9�h����x�4�sY\i���S+Ό�Ls'Iu�(�������u�0���{c��8L%ALD�P��k#�6�S���R�=�0V��M&��F8���L��V�3Xb��̡�w$�={��T�d��D�����b	�e>3�e*����*P$I���s�D!�	x`@:��^�6�ꢻ0"돜b��$i�V�d�ח)釂%M��̕@$�� *�;����/t��J�z��95�����:��]���_w�d��>������"�b��҈�*�0�E|�׿�Z�m��	�G���yO�G��p���E�b� SsSe�h�W��D_��Q����7�{I�D b/#"�H�Fq���r�����3���.�Ք|w���[+�����3�,�U4��I�;>�����k�X\>tP�<,̌§ ��Q9����Ÿ�G��6�ڤv��a��[�t��hH���x#q���Z������!�eJ�!�i�Pd�5��Z�^�E1�q����سh�3�v�� ��6��#�~3ɖ��k�a���Psv��� ��+�/�l��$�&�jz?'0���X��Rz��D��>�'��<�}����Ê$�լ@Z�m������v�-ѣ�$X|�����unN�fb��R�!�Ņ1��yְ�n�!���'u߀�a7k_��IN8�Ài4��U�d�줹i�
r楯���Xf�#�ߤ�fu�A�E��׶{�ˈ|>��Vh��m��+�O��	R�ފ�O��w �2�~���a�)c�|<�45oF��\�@��,�����Q��^?x��:�H�}�bp����/�z7��#�ࠌ8��a�����]���gd�� �yo.��)�(Ӊ�
q��DTq�p���x�y���4T�Ռҭ�(��@{Ӄ��>�N�#���:�S � Y��y�ߠw�|� T{?�K�	sp�]+� ���-)�B��%��$��.ٜL�N��s�=0�\9��?z�6[��=d^�V�^ۋ�{װ���4�<���N&l�+8�\�v�R�
ɐ-�Z�AEVj%5��D���M <�1�<uY����r���2��-|�󵭢��S���?�)1\�������Ei0�E����۫�Bm�_ţҕ�zqY�F�\�����?q�HW�8�%I�R�w�<ޘ�Η���Ot��M=��T�w;�6e�K��@�g����S��Q��B�=�o\�e�T����2΋¸����X%�P5+�v�钥4/�E�u��z����rԮ��§�*Q[�5��?4.���'^�e�O>P_�����WZ���FF� �	o��
����w�y=f6��������H�����%�|���Ն� �����\�kqA�kꗽ�3B����`�����*"!�dTC��Gy�y���	}9�'<�=̞]np���p�� �5l~;}���5I��ڟo�aDwx��j&�����F( �t��uLa�r�'F����#u�NPgn�X�= �z��/�(U�p�3��LV�Xl>�D��Eo�eW�c�� l(�('`���A�����%7�Ĺ �y�&�H�g_*w����u��4���X�IDe�pz�<F,����I�73�ރ$��p_�R����?���ۏ#�ܒb����Mu���Q��ѺZN=0����'���pL�xP%���Xy��Z�!\Shݍ�-��R��#2��+��.�D��G�_ꙻ��{\f��c&���C�!�|4`��Q��}�#3���j�ʙ?,Yɺ�dh����x�ТN�������}a4̳3��p�E����9.u�\Ha�	9��]�V���Xkv���+�ki��{�x�+������|�l�|���5� #��bw��tZ��%������吏#���~�����x�쫍���V�F�%���q��z�6�������~��w�ɱ,V����b�)JunM���QN�L^����X��� ����<hDV�]4CRS;C6v\,Ny�E��S��o%>���5}~�?&s?h�~��U�5)�@��8�G���u?t��,��F��& ���'I{Tf�L��Y�U�~*���Y�7�?��+~@t���U�����6;C�Q� *0���&
�h�:ݫ
e)}Q�۹��������T�g2hx��g[x�$�0jRť8�-���*-�[ZѸ�_�:MҟT���|�r�:��4QF<f�),�y7 �Jy}}>A��6��JA�oK��%�B<aG=!��%���-��R�`��F��B����xԹ����f��?����n�~H��	�\a>{���	 ʙ�>S��X�|q��c��2�9���L�㐞~����Tں%��' �����.v,4���9��2\�l�F�
����M�� ��m$X�vBK��(��!�\[�!ʗ����#��2D�JGA��c�� ��Þ˅���8�`9��uof�:���JI܌��ƹ</1B�NuӚ_{��q���Z���t銄�T��d�{WY�l��ee��5m`��;��Ѕ�� ,���j�{��	ʛCx��6b��v{��	�>X:��1R�6"�u�oA���+��6d�%1v�| �m�����t�DK&�i�O�	���B�G鯜r��;K<�(�,n��ӊ��h_E�@F-2:MQ�F��CA�3�D{�N��U��K٭y��2��$����0>Y�~鲢�e�q��.G�[O��@�4�Ҍc�%i+�:�dp]|^:���z�C�\UF���##��/�y�!²'F��fe,����h�O�V�-��4|.`K�=1���M>!����)�_�H]jZ��d����kI�v���뵕��π��\�Z�
�j��p��ՆȰ���|�R�:��^�}�*�|1�/ nx����K��i,`w5���<@�d"�t�E/�O�<����ޘ��NG,�H�D3`WG�v�Y�m./<v�RIW�f�(₤:���V0��Fw�����t���.�x�T��k�6�g�]؂v�EqQ�ˑ��N�qG�Xl����{[]���u�g�% ��U9��ز���L�\�8��\�9�e��vk�(\6�G��nW-�RFK�W;=���B����`���m�?ú~�B`����fɨ�F�(������Kn��z����!15){I����%�4���O!���ĖX�^o(��ô���}�,���V�ga��7�QQ�*,�J���`�j�BM8����o[Jd5
�bwkN&�&|{����MUwK$yCpB��xB�Ȕ�g�-�����}y��уТ����!*�m�����=3�# Ĭ.?"v�'>����[& �)+�o����i��(�^�y60�8W��C?1昡Ng�/u\�����,ݯ�T^����_�V|�?<X��}W�����_�D{<���ɰv}hH9�#����E��O�X�Qzŷ�&�Y�����.x����D�sL�ꗘH�7���V�B���B.C|����?��ƭ'�����Ҧd `<�ޞ��u:
+�w�O@,\���W��V��ai�p���E;��ҲR���w9"��
�{�Wv��0���������nOԝl�oG�4�H]�a x�-��f��|�
�L�5L�̧r������N�����(���76��?J8���⯪&G�k�����茡��ȋ���(�a��,�cT ��;g�j�����Xtjj������m!�G�g7r]U�����+�>�+Ϻd����R	��+��蓰t��tk{7��h���[p���|���3��t��Yɦ���[�g�`ǝr��.�+�^�A�M��C���JAJ�qء��rx��5�М��tgm�cL����xFd�D�9$5�ӫn�V�_1�`ۣ�P�ėA��� F�grGp0@��0>ؙr��h;J�����@�����(~p�@�{krLe����O�=;|h�p
��Җ�5SRm̑Ǒ���h$*f&m�g�-�˲�-�1�*�܏3�	ut�o�Aҡ%��w�#�v̀�'0@����i����Ӛ�����dIu�HIG6�������Z5�� �5<À�r=TR��Y[�k��W%��t��:�$�$����2�G��Ϸ�<� ���?`��V��1�2�pg���L��4#�e���U�Rѱ�����x�fS��gTU�Vu��r��.T�U������GJ�[����+Cg��->��*��b�h�y�ܳݕ{���<���ش9�1���9��"&�64��U��l)^��-�
�1���.�1�:�C�9��d���/����Rћ�浒&�<bZrhP���soҊa<��Ҋ����Q%5d��� `���٪*
]��.g��o�7��rz�jqF�{$�>��h��
�{�8^�:qk�
7��ƶ�l�˽�ϳ���ZX�E�V.���v2"��
,�z��\����k2l�X^��%PLn!SE�;����ϵ�k���P������흳QUS��+H�x�&�	x�������[栉�-(�V#d�4	��RH�d'0;(��:$堼l緣�t�o:!�0�oy=�1�8t�$������\�>��3p]|������dǢ�Mv��$�4'��I�2X12kN�5 
�ͺ�R�@����R�$~�{1c�6fR�Q�,�֧Y����MUps𵅡D���&���Xt��Į��5����u��@�%��*�k� sˬ	��������`�L*�n\�]�a��L�ʂ�:(ohwbM���q6>Ŗ@�L�E_os��2S��Q̕E$�1�����wĵ�|l7���I���2�.8b
�3����s;�T�:�
�꭬P�v&�t���L� ���E�#�!iL�l�$�%���I�O\�u��Ǣ��c�>a��A��j�|í��f���Ch�=��\U��{�ŀ܂p�� T.�`?���P<����NQ&n�(�a�_	]��J�N�Ԍ&����o �Е�c��;�6��sˈ+��ai5�A]�s�؞�;�\	w$���� �R[�KR˾!���ٷ9���CW��My�������X'�D*�[����QCv������$�2�|�5����(�Ek����Y��� �ơyujc�V�ĎM1M	�C�M@����U%=0yq�v"� �Ip�ݗ��嶭rs�'�*�U�2�@�	|��X��ǧ�]�0��t����R���Y�j��.����_[&�8���7��\dAD�&;2]:�ZE�ac�䬛|~0z�Eq�i=@@Pp��OSJ`�<�a'>�P�Gȑ�@��o]�~�+���g��򁌢�0u�<ɦ<�k�æ��GQF�X�7S@^�I��+)���k�z'_�P����*�R��l��B`yKhFP۵$N���\��
�mT{cO�b��Gu^w�ʢ��G����A�Δ�	�ſ鏯�c�;Ƨ`�:&�c!�s�n��i������zP^��TBëd���yݑ�K��/3���ᆓ?$���1����ù-��I��G�9^�bU�u,N�����J���C�WB߆0��u�S�0x`r���!�*dESxϮ�>xZ�s<^�~m������q� ߺ����˖�h"�9MRD��5����?lH���noR#�	G���WȰ?���E���\�NL{�����b��H����B���.�:Hw%Y�����2��}CӮ�0��Fk���w�����U0���~��E��֚�Ɣ�*�6TN �F�o���6��?F2����_=Q�j¹w��$}k���fF|&���o����'k���?-�T�с�ʹ� ��c��UE��*���'H��|�th궚�Il�0C�����)��hi����9W�&�S0��tN���S�W���-�D���p��{�q��v�쒔�k��*��w/�S�;ʁ�1�z�����CQ~~���X���dY��*��;�٫�P��_�E���6[��Eі����͵&6��֮��1�H�:3��Nv0~Y����Dq�$�U�4ȷ�}˯���O!b �K��aH�I=QE����Z�
\�>���}��1���*����c{���Y#���Jj�~`�#�$ޥ�����n��*�^146��������í֮��E�S�T64���UQ�W���3!�V�o���$�.���4�]��V9FM�Ҥ�~��˨i���d��O!�*�nJ��8k���(���C�~IY�J�6#鬵�iM�lc7���ܪ�ު����F|�ܛ��D���K��;k�[π(	� �d��M�+����u��za�!#y�#�!�۔>|e� {���D
��fેe'\޸Db[9!B���j�y߮N�׍o�BZNFڠm|�'V�(�0���m߂��'�m��0@3"�r�Ly�|qpok�_�/Ƕ���HI��1��-: [�Tڨ�׾�)Q�.�.%$��C:�up	K�_�5��`�ǉw� EEN��Ub~��!Cc��ܡ�}�̹&��A�u<P2����o-2����[��R'��G���7J핞a�"lmǯv���ߡ�U�&t��8�n_m��g�W7�����i~�S��&��:̠�JQ#D���^�J��G�2�mr� �`/��\����j5h�����ڧ)Ð��H2Ȓ[X=� ��&0g�?�g�]�.-c:W��g�4�z�;��7���Ĕ�*�N��u����������T�)��KFN���l.�ڐ��/!�6���k#���>���u��G�++(|O��@�B��C�A���.`�e��b3���@��OH:��nw��H�E*)��*5j2]�O0h��J����i�C̸�w��cN��G�3�!��<�����v��$�E"$�)FN�jk6�3д����܎*�JiΒ_�xjI�
u�5؎`ڀ)֢_ R��R޸7kYul'��7�o�q�m6a���0xM���lDcjы�/(�DB�Ҍ�2ŕH�Ƚ��/���KKAtMl�*s�����{���ŭ�E������7�J�l��%���~���[L@����/�c~�m0	l`���i�W����
�5s`|&� �kcX��o�>b7�h&��&$T��F~#dA@#���k/Lq�<��:�i k��g~��8[�>����E]��SM�����aMQ������� Zזb��Q�k���r}��tR֎/���d�&C�����	U�+�T%5I��}�]�(	2@�%-QC
gX�i�8�w��\��5���zJ�j�j��}���H��;wWf#��y+�yF~�W�(D;�Z�4қ(���V3�3���C�������db��]���L�N�&��uH;�%3jq�m�m1M���v�y��jU�|�
�$��!�P|� df�<���R�"d��Ͽ��ԍ��'|&��C������[$�r�]C`l`]T�N�a\$Kvų�p�d�3��p8�̱GQ�x�e{Ҁ���ܿ)b<pzT�#��Jc�3Y��&{nr-#wT�LE�K��w�}��|(@��t[7鳬\Bղ�����97�_-���!��#C��Ю����	��=5:�����&�3�	���i)��˃L0C~�ܠ�!Y��a�U>��2V "<c���,䤠��D渲;��,�1p��+�4R���3��--�i�ƨ�p&ѶА)���R�.��;�},�����j�枣��lE�ֵ`�e0�����F�'�����ħ��=�'��G��Ŝ�ӛ��"% �d��3�g!hq�U�1\ㅿ��>�f�9�w�e���K -k�8�2���"�:����]LH[&���HL��ȶ".,}�u�~���O�L����$�w=
r��_���:$�"w?�����h�ů���;M��)���d��)h��q��/���vq �4�(ۥ8p=�sU��:��2󹣸@���!�a�X�b�)Cvg�F����>*��8��h����B�-��i�f������5X-[���FR�e��ǈv �mʗ+�>����5A�՝���+9����ux-��.���C2HSZ���,S�d���&�8dl��	/m�Q�a�-�����rg��,��O������"�����TT�|�����/Q`��.p�Pm�U�����<x��"�4p���]�.]��ֶ" "�,�P��Z�d 3Z�F���:wP�n��\��-#��<UO�Fn����x4Y���H��d�.��^�TH�MN$�<9�Wa�wq�_9�ָ0c�����u3��iR�O�~��ҕ���n	&'NQ���Ya���Δ'(�jkE�E1�T1̒b��ǜ��׳
����%t�?Ẅ́5�2��g^kT��[��h�%g6�t�7j,�I+~H���jэz���~����,��BȠϏ��-��ˡm�o�\�w�IutNfԴ�{��ijȇ����ԏ�L����^�DzEw����8b�C��m>�ЖAH �l:�kG���)��"0p�џ���a����.z�i�{�zP�|�:�Y~���r~��H�r9&F>�=dj!�U���P��zcf��
׀^�Gw-2F�Y�I�?~`2<���Iiɳ�k$���T��jo�	Xux{�TQ�W�
�<34���3I��=�.���o������������|��c�ԡ�Ev�X�ʿ�����cz���u�r��b����(��e3��	n��ƞ�YJ��J0n�B�s᮵��Il��eu٠��6ƀO.@
d�
�B��iR���ӯ��Sj��&t"�}i�l�F}P2�[SQ@��/�a�c&���d�[(	3�=�&ym��n�u�Nȡ| 6yhғeDAe�҆"B����M7�&A�m�\I��ǒ+4�wל�e�I�>\��Fg��v�:�s-�0z�tG\�r�]؞G����Z��p"(֖�����s��SqrP�U˩�_��5��br�,��dbu��ٍ��6y��QG�Q�N���ICW�O�OF��z����O1<�S���=�V]4���2�@&e`�R�?4�r� ��*Y!jeϒV%Yf"@�5�t�����T�R<�Æ�"���"�0�I��iκǳ#s[���nr/��V����"�ko3�)�.N韂��9{쵍/a��P=�@5���6K+wx��x��w�`'�rA��V�K��n��ۚ=Z�ʹ�Êښ�Z;�������`H~��+
6�`�*�(�;U��臘.�᳢`�cD,V�*�P��]|BH�C�T�b�L��O�ޣ���2/qM'4u�ɏ[S&�~�����xm\��D�Xr
�Z(�V�9<��8ap�s|�ێ���W��tVXB1��x>������N�{ǣ��]��/>��e"d~K�q��q���b�&��sE��|������"x.�K �zGX����k���K3p�ڍ�tŞP��.�[D/m�5!\t�����u���Y�'�c�{������4��!���'%,�5j�z�
t����j�Q�T�%����#!��Su
��z7´��b�h��}g�v�2�uF���V��2��UKc����.pgm푦4*�����:��s˿��PCz+��~���<~��tdaʗ��d��ɭ����vo�PB�����*# �*�1\����
h��j�+��&_��X�u�;�W]�F�'H�\��0�W�\��K�i�Pv"AYp6�*c:us�o׻�Y]��ڏ����z��Z�cf%�"�߈��󥨁�t9 f��cJ�У��&x�w@�������ׯ���Gf_N�Y��a~#,����2��1�8&��ȹ3x=y'}?�w��⵬mW�͍k�Ω��͟{!¶]}���!E�]�Ռ����
|޴Gc�i��ñ>�g4W6ӥ(p���Sޫ�Y_z���*kNg���Ǖ-���?��Bv����tP	���6_�����G5������!��;̿���%��F`���c�O��J� �����c3v�ˁ�M
�A'�--d�0��p��4e Gr�Bq�h���O��8��]�dJlؼ�F��>�&�]Ώ1����!������*���l]��D?*k�tb�����Ua[�&]�]a#V;��b9eӵe��D��e\�-M��df,1�W�B��F��1QWZ(_c�5w6MR�XXdIF-P�rF�(����9�UIc:R���fV�?9���h*QvU��|�K>�3	貆�3O}V�q����a�#���|�6%S�'Q,!���������tN���bb���8�~o�Vj���z�[9I�`�@.栠+f���V���}*��n��P��3�1��`K`�}�/�m;Pg}��.���gc�g|�h���Ԉ%��X�	����u�y�����oz�%��|�,�9���E2~2���o"��(F%U�L�=-C��Z� |0�q���p��*q�|{�#`���wމ��,_��`q�R�̇�+fӶ��a��'G=��-h>WhEXn���۱w����_���J��Dmd'd��L��6���y������۰���s-�S�'��/��D��MW(2�E���:��c�2��r���ɐ���,ANN�m8�2Ε���.��/��¼ٷW��Q����{d�r�Iq$��j�O��xC�=-�1�LIm�[���Zգ��������b�YI�u��+	྿�ٙp@�~��E0�?P�5|��V]t�c�Y�G,[9�Y�Mi���=���2H����g��W�'�+;O�?��c���8�C�Ԩ����]n-#�4r8?Wp:�4�����s���9 �A6����@:�i��m��?T�N���k���q��o��s�ā��k�����g`1�4��9�g��t}�L�^MI<�{18��R�xZ5�[���!�@`5xP�Q����G����ġL]*l���B&��C�`fD���zT���&���x�'BA��eFdU�q�ݮ��3ß
K�F%�^[?@?8I��Ѥy��,o_[�VlW����� ��s��,�)�[{|�o˜�T�ao��5�V�`�;����\��_��}.�FC��K��o��T�]s]q��ӑ_�16j���kW ;Dtd�����D.$����f��j�a�?�X���0M�-Cr~���h! TG�<kv�L�%iXk&'r���ou�����K	(����P�&l��,k�����gV���=�pᩬ���g@�bܕ����xh������l�����V�c)Z2�%��q���cz7�h�x!��9�(����=PYwx$o̈���t��3��a�S]�@w����L$YUrGLyAe���n�������P�$(�zu��(_g�'q�Ů��^3�?+�=��u�'҅r̦}����"���>)�On�����/���\REKi��㥅O�&~�<`5�n�ʃZ�s���G���?@�Hy# n���?����t�&�S������E�r9�ߪ68̜qM�V��R1����R5\?,�\��Y�t���w��7 m��^�'��"L�[}��'��,��[�rb�`#���4]H�n\J����s����s��W�}�Ϫ��%�<cS�*��^)Ѯ7D�C�ͣ<�
�b�'���&uI. ;�9,¥z��R��'�>�Ik��!B����:[P�˱ ��2�K�~�!j�݇�G���+و���CL���D�5m��3V�v���o%������������<�xp���c�-�)ƒ���$VOm#_ �R�Y;�9ݟ��\��P�{�#ng�t(���ӵ�6SV��KTg�̇Tx�|�:P0d�����_���&DC��#s`j�&��|O�ta����*Ofο��K*�/<1T��!Vq�()�(��9B�B��Y8�u�q*ߗ/�f�IK�2_��ݯ��/�;��nJ�x}Z�2al���s�$��q�3��1�d>sX�,@00q=.P�qB-9����s�N�O|l	���o�}fD���\�Ԧ�<�L%X�^ߝ֐`�� ÷$�zS5J>3j��������QG��Jś�rg<)s�2΃�=��ox��*���K���He_AO�������z�q�Z��m #rг��Ҩ�gS�W.(K���Qd�`��p�?�F��!�Vw���'A?��d|�DuxmF�N��c�"^��u��^v�y�%��T0��\��İJ4�6�90>X�<xk��UW�X�z�%.�ҡ���m♌#[�T�hT༮�)[Wk&�g�_�9�d�l���6`�����R�1�czеH�d�8#WLݹ�k<��������Fh��oX� ��+yH>��@H�i�2Q��%�6���)�?6�PSb��N+=׬D)�.����	W�[�ծD.�V�k�V�}�/�&�nyJ�@���8��Ĝ�HG���_���_��y�,1c��8�-�n_��d�7Ll2p�jƱ��͟|��:ܔ����g6r|Ι0l���h�|�S��1��,9n`��Xz�,�A7�7����|�����8'=����6��,�@���C��R����߹o�"���䝽���	J5�Y�;h�m,y
>�^r�Z�a������m\n_���A��k�D#��tյ?�����1�c5T���1N�΍�x�SZ���3������c�岦�˯���=bĒ�VhGih���3i$h������6lက�������c����i��߃�֒1ܭ6k��H�/���f�M!எ�I���?\>9����Ļ��y�u���x�Sg��'�rɩ�����8X�s�A��Y��ؑ���ӧ1��j�d���qGDo�-L%;�ͯq�2E9�C���e � ��2j�V�S�Ew_�7vۿ2��D�}��7�?�6���%ȝ�nx�3��S��_Ͻ�������ɬ�}j���
6�����ю�f�'�`	���w�Y4�����m��K�gD%�a��O�10B���"3Cإ��=��kEc6HF��B0`�C��l����LE������4r��jP�Qv�_O�3�%ó���!y��<��ج�rPa7�[�9;��r;�kN8r����Y�=c6�{����6TN\i.��Z�S��tF��R��IM0�OkICV��U��USl�Ʀ�b��)�?��t��ZbZ��!�4�vf� ��zc�LDg|��ekި|�'?���p�h����!P�lQa0?*��� ��Y��f���fI�a��}ؠNX:K�QS$��4�O�چ�|�c>Eu�6���LR��$o�V�-'����qy��*�j�T;i�r�j�	>�h#�wm�Z��f��K��ܮ�%�g��k�qC]%�>h���쌍�ɸ 5m��)z�hȴ�参�����M��z4 ��eo�޽=8�kѨY�.��m��A�)����bVjH@�8�d��Cd�t�4������ ��qR阣��/�=��_a=�g���f�%1�/��n�+2��moUl�\�|"z����Kr�U9��YR�(
f�[����\���u�e��? �>��<I,w8ڸ�Y��8T��v���6���2�����/��0�T�u) �%]�Qz�%ߖؒx���T���5�@��EiZ5�&@��3#��'oGcg��+����mt�6H��Ec�}��E��i�%��ES�T��q��"�Li7 H�uYEgs|�rG:��)=�@Do
7ܢ�=7��AP�Q$�����l��C
�!J��~r��.g�p2�OO���=��,���w�%�t�C�rR�F��\�Z�Xv��l�qn��{?
���)#W4v��^�\'j�'PU�a��5���*��=��3@���S�JK��.��#-�;am7��ҟ�R��jw7�֓�Do��oB6�$[n�5Du2�n�ؽn`'z�xÕ���(��
���tqq� (�ԡ��m�	U�, �۵��ZMd�mPQ^�H��L��.I0��Ǒ��dgEQ�e)M�bh� �+��Q�ӌE$���B'��6$)���Q	_ѩ(�p�cn��0 mB{�N*'�w�� Y0�A\��K�톧8%!C�p�e���d_�U����}F؍q'{��\N���?�
 ���H([]�*\�:$�<�B����*�,�b_te�]8A>�4�8Sڹ�
*��}�?(��%=���ck���C���>�5�`��_��=�Ҭ�I���p�S�.�ar,��	D�l!W��h��^"�n����/l�T-�RR���*����OD�6!1h����9�ay�*[�5�z�h�).�w�767��*�Ӽl�Q9�U#�n�Ԗ�|��uSH=��ͅ4e�^���'�t�v�`�3�C���B�NF�m���/�נ���~λj���J@�H"s����Q@�[���ꑯ���.���3o`�T�Gʣ�z�����,]q���8��)�ƻ�
�S4z�u�8 6�W[����7�����k�e*E�:>�*׿o)���؍t3/~��v�ҩ�
Y��-��}��HP,��jl�B;�Q
$�X�
V]T�-N�VKz�V<k����]'�1Ꮳ}�q�~D�[br��H~Ykx��.O�s�����I���ӟ�
/|���~�M�+%G�M9�����I��֒�D���,`9(�)g�\(�/�!̦Y5A:����xH��#,w9n�i�eF>��YW&V�t�[�E�	�24E��g.��s��+�쪐ٔ|s܇�HqK���7IM��R�/�Z*˷�\�r�v[��\{cJy��OՐp3	��Y���*õuB��؞��d5�>���7�]�X<�kz�w�Ɨ�d�ɥ�Q��VsJ���A��L�WP�
���6O%&��mS(L�W���x�K��N'���p�a�8�_�����S�`����DR/�C �/h�:]�s��[��U*�r�<��T,��N��̝�[��a�0M�W���ƕ���H/o�μ:�<đ}`��m~Kú&vZ9�"����!0������rC	J�B�.��k9BTU��Ƚ�X.�з�����%?������Zz���IqO�=��{j��* 3���=��QH���%�^YGn���l�a!� �U8E�m�d`�;�@s�9bMBş�L��Wb@;N�+&�S�h&&�5�b����5$��S�[1P�/"��2��g|������,���ҍUn��8!��+[�a�Ⱥ�A�JP�����Ý���<^��p��R�����?wu��?E���ٸ���Jr9X�4y�v���7�
�oVQS5����i������Sߩ��14�˰'!f��晆՝L��*T7]�b���M�D�pF�/2F'��b�lB��7�㻥�'�%��ӫ ��,#_u���=%.�\1F��X�D���GD���䜦_0;[/!�Z����gw�k�ĽsT�P(!���H稐54x��/����/d6��Zi4X��t"cς�GWٹ����b������,+im�&TZ8Ѻ�g�ЪdT�D�)J�u���4�m��BN�Xqaz��-�"5{�	�_�wʙ��!��FY�$��[wX�)v��Yy笌�`Q�9����ԿW�=$�_�q\֭�8؇mO8]������$�,��a�gPw���1j/WZ�S��OJ&�h.@Z=�rS[���ǭ���_�1�(��3���J;|p�\*\�FO)a�l`�[sk�����E^��Q\�յ����Ȝ��*�3"�pO����e.!�"J��WV5)N7��u}h�|qR*�5��(��NǝshL�����,�J�Wl���@jˁ��F�n�_�v��j���>ɒ?�&�~zh�k������3[��>w�"����[����~�Jխ���W���Ʋ���;�Q��\�A�_�|��[1
��< 'Л=��VYA�pUKor=�7$L"n�]���fƣ5.ӊ
J��@���.D�}�/�4����)k�9�]�"S�+�+?`/��՚6��"b��!�֠"���x��j��m�C�lGvW�N�<�\�GEO�Q�8"> �AW�V�>�JH+���L��{ޙ�I��!Ȍ]���7U�(���p�|��uׯ7���OPۤ�Ӑe�,&��^ĉ��V��`&E	�^{��r���9�ɜv��Μ`�@�'֮�s��U�6eo� ���������J!�q�E�]i;���Y��F@�e7l��������,�L�3[�a(�\뻝F!!/I��V�28A���
���WT2�J3HS*�Bl��YW:���,
`w�/О6T5�X����8�O�}�chJ��L��7����k�W:6�dh�x�"W�$*Ǥ��dp�����n��{0�Aa|3V{\c*[���\Җ�S#wQ|�Ĕǲ�du=e̎����O����&������E,Ң̪���@�����ȵ�@"�h�
B�^@. ��m�ѭs�
�����֔�wm���B��`���kRo��.��(	r��8-���p�Q�vl�!�ź�[_�J�w#۝i���)������Bs���`y3�S ˙2�gp*�=�1��k���zC���O�kS%� ?0U걊��@��Cơ�2�ӓ��h��:�1CP��~���?P0����T��P^PRU�����SN�^�Mw�9̌��Yl��J�)N4�TxM[g�p>X5�J*�Z��|Ob�]��)�tT�c�:��ً���"��Ug"N�Q&dFn�7 ��7�w�$=�  \m!�:�	��O���Y�������=�w��m��c�D���X5�e�7l�;���Kرהw㼀f""��l�(���`��E[5�dJ�~m�r�sC�������
Z$��674)nY�&�$%Czn΄�����4:�J�/����9J�K��O���ga �� �0�#siz��HĺF������5@x<�$D��K�>׷b��]�ʞ��j⼋�ine'�&ּ��<�Q:����P��c���Xx�L��T�.��5��]\�1��a�75tTQ���r��RPwLf��O�R�`�D��b|�М <J����7���t�a�-��J�HΟ���-��\|�m�ݯ �>���*�S`��	ݒR1s�
�)�I@^تAG�䆶Q�#��脧Z���E�|U�������g�u�-��:�b$w����VX����q��T�?ۛ���������X9<F�-0�7ab��(K���� ��
����cRl���T4	�tr��kxcVO��x�E�2������B�� ������H{8X�+~���ڪ�P"�E?�!�m�|8X�>����qkf�k��Vg��~CNO���ؼ�1p��@�)��Gg6�E�l�TA�y��J��D2�`��H_m�h�œ�A�WZ�Ӿ���6�FC��K2��Ƞ����cO7����~yJڇ��o��`M�;!�TZw+�x�~�q�f<A��OE�:1�F�:u�8���O��-[�G�GM�~7��b�wV�	�
��W�+�o�\�j��P,Te�v�-��{-M?[G��r�T����ج����x�b�ګ�Ɣ`�`�(�)]Գ���E~{t��̧Ά��:J,	����V� ����ZT8�.��#������v:��I�Dd��*�7���ȖZ���Ŭ��9�^����@yՏ��|.�7Xq,e�sml�����6]Œ�}�U�(ƿ��ӿ1~�u�P�y�б#�x[V���"b�Z�2��Sٸ^��g��.
j������0��l�w�X2�#���W�(a�r�Y�7�c��h�%9�+ⳙ�Kh��~4G��ܨ�X;$�4�7l���r|(h�	�}L��ݨk=F���_u��a���o5������OOS�n���S�(�i��[�n�,ڳ3{&�{d�=D����4µ�*��^<T��ץ��	�"��GX��qw]=1�+��h�)���ˋ%R���D�$�´�Mx��3*s2�Mc���´�u1i;�A5ߗՁ��F���Ā��0/����u��Ũ�B�i��i�=��Ԛ�v���C�
$�e4�݄g����N����epF��d^Y�=g��&�S���r-Fv��Uܬ#8T��1�ի}����_�!b&�#�����m�.�_���Щ��HA�]K{1#���MIM��[y"�Z���|�Y#B�-��N[�A���?I!+��ר�B��}�2�<TD���\��j�ӵ�����5�\�ql~���X�����moN���E��7ם�?�&���v�A�Ԋo{�|ڷ���|mz�@ ]'���d��؏�f�J�h�S���]hx*V�l&8�_&�૓��>�*�Gdlx972����1���9��CU��ǟ�kte믚o9��� �:
"�%o�-ς��	m���-*��^Tބ��`v����}]ߦ����Ώ]�9�s�7V�W�ԓ1�\s�wڶ��6��"��V�9�W��)�_�
N�zK�<_5���ت��ŵ�YF%�!�G39GpbT>E�zx)�LWs1gU�xŌz����HA@UK�/&^�׍��I��j3c\ۯ��$��������5uU:@��7:o�h�i���
O��E "�~��S�_@����~0ܱ�*!��熰��:5�I8!9z0<�4}��W�Na���
�~k3�B�S�ţ����sX!�We�*M ���-�P�Чr���+z�����G�W�"<���$��OϷ�o$��}�r�����
19xg�)�����%�K�[��y��5r���������!Wb�/���S��;���B��ߛD}CɊ��i�e�m�{Ԕ4�e̤rѕ�Z���9W�B��aL_�=���{����[��*>744?�N�-��HV��^��a�=�ff5��Z�sT�_������}�j�N3�W��^��ȡa�L�2����;�s�@]s��bZ���K���5)B�?���
4��0�4y�آ�M�3M�p#�l;��#�S����E�����)s����^޻�2%��O��<��>y=���)A�6:zU_[ �Zf�Wn�B7]����>���N�Ͱ5�G��e�?��є�����yG�B-0,U��wrJ�+PPQߒ=c�p��)ط%��8Ю�	Hn^q���ph3{�,���t	Qۍ-��oK�S�2Z�����^-�/@An=|F,<' �9�֗�CFl�|��G�I�� *!f���~�wC{�_O�X��v���`њB��tp@TJ<>��I��RX��< ,�Q���fS���;ٿØ�H�����*2�� ��h���/�-��$kU"R�Hi	xCv���C�
�]ȡ;w��ߍ p��������־��$�D���R��d��bl}���Gve�>�=�x�U�L��\�Ru�	���I���H���<��s��3j�$�PV'54�yS�(*Oذ��%D�m#�T6x��Y�i�v>:��WK��8�l�j����s��(��AgjvNA�au��´K�Kyc�{��L8
�	�kP� $�ʰ)��`�Y6�BH���*�Wt�]o;��|��+��0�,�ּ|[�9�x��ϼ�>7֫��i�#PO d��V�c���zу�x{_����ǭ�g��a�\H�6ǃ�����2�q@0����pl-k$p�7u���(���œo�$h���2�5��4�VG�7���ej>�o�V2�^����!T�e� ��\QRa�d+�2F���!���CD�#��>;ܟ}����X2ck�����Z�k"و>�L;~���s�D[Լ)�w78q+�D)�قL�*�!&�?�$Y �BЮ��.u��ɣ�ڊE*S��b�R�N%��R�J��S��'���r��>s�a�ʈJ��F������-�7}A��*'+�ǩ��7����WЩZⱺ;���F+�k��ěLLح 8c��gƤ-���V�M��ϝ���.]:]0Aw��v R{��4<���4L�b+I��>3�T	�V1#������(�O��n$���"Ύ1���ZE>ꔃ�~��XW��V4+l#�)8D��6$/��a����Ih�XQp�<�3���߾Y2Y��ʢ|�?P-ko���wl!~���93R/3�ae��$�E�A��_!�� �"��T�8)��{��8�?	�*������!��'�_��,�!SL�(�Q��0�(�NKA�z,,|��������-U�n��\q��$�`]�sa�K�/O Rޒ��e�Z� g^�@�Pn=��4~��s�l��r咻K�D8	��{q�H����Z*��<QӪ:�e���$t���l4��/$Mot��f F_R��w�W"i�����u�Q|��	I��˔���X�zpgq]���̷j�^�Ko#�2H��$�D�)
�Z�a�����6��QUa�RàҎ��4p�$憁p$͐ �1�~��'����=[yX�I�g���+��������*�����4�ŨѲ�J���B ���FͿ�?����k�PM�C�ul�7�B�ZPH+���R���ᕫ�RUX��ީk���K�w����uтf��wc�uݖj���/TN�}~�t3.�n�<��݆GX�xCz'�1d�6C8�/0		�Ǽ�ݽ�(�vP�5ᘒp�y�ƥ"L������W@�`�2��>M�����g���JB�ɘ_3����EN���kc��JM����-2*��yh{{�z���,~y��M=��@7�E����>	��y�;?�%(f6�k�߼ U�L�ͩ ���p����]Z:����N��N	{��Hݍ���[��d�e�^w��ݣ_�jaM��,Xɲ6٪x�ot�R=�����C�rf궪���Ȁ����JL¬�,�	���� z׹vl��3J���bvgZ$��*��fN���}�ѼɔE�4,G��c7}�^�)�j��!:>���J� E�� <�*�-��iU0�� V����>28�����W�?!��'B~�tt�㼑�˚����j7~k�%k�P���1O���E�1<�N����!i�g;�NǸg�k�P�㨿){ �j�UMB�����D�V"�OL�x��*���3�$��8؟�=YN�Xxޛ���!�a�偔�uO�I�qsiO�f�\��m���J-��5t���mS�V���D�AU��M��vө�ОCj���N�8��S��vcK&']L�?�����Ao}��ך�B�>�U�~�:Go��3a�w]�+�h5��hǾh�HD���JvjG�<W|`zT �@=%+�]��c?�%�|�y��P �m�Є|� �(�߂&_���be��l��s�\L/��ݖ�:`��"��׆B�{��<,-�g3D��Ɖ�3ht��<�P���Yz?��m�VU�

,�z���=�h
��\'��r�A���j��m���&g�d� yɣ�Q��֤$<W��`)�̮F=��Ԗt�����~w�9e�̧�4�Q���4����^���~۸:��">�֝��
���L/��ͩ^�M���>�=L����K�m�2�W�ƈ�z0���=m��H�j6�[��`v�v)�_iU�au�W�l�X�qVIoI %*3������/��	o����Fɢ���Љ�O^�#	WV�S���Yͻ�T5}6G� ��N����0��.���"�F"�����M�NS|�Y�<�.�^��P������ߋw�d�w׳=KB�M��x;����0��򑢡t6L��p��^')��Z0:�"�V�@��{ � ��Z�M?Ǭ�l��1}�GҤ�B��~I "��w�}6�@��R���[��B8�8�4��Ϙa��� Fo�w��ؗ/��}-N��E�YuO��}o�[?�s]��Vs!�������t,Y��~��cr˵2o+V1����(�u+��6f�YI�:�]t D\��Q�\�O�޲L�'M&t���{��&>>��nBq�) RU_e�Jf��-�,}~h>;�@4�f�>�|\�:-���*�:7oP�9���١��$"R�6�����@F��h�:������	R�b-�g�FM$g��y;m<D6x�4��9k�M	��C������j�Q���=ӌE`=�k���U))<{m(�
Z.�I�Ň� ����E̮)�SU���4X��]��) 39�"��(d{�7��d��Y���M�@���Yk��$�D6��+�0=�͗�FI�p��n@Ϯ/iW>��\#�Z���ďIȫ/�m;e�T�I!B�L����D�.q��YBRc�ٌ.�RC���.���-[[��V��-!>�P�
_�7����(�~\�	zΑ������C�c.��VgO�����o$�S@��j��Q�T�A������ǫ#Hvy�k%�Xy}�%I�j�q����U���P�����\�(�4 \�@�Z��_#�g����Z��GM�F�<ᣂ��� �R�ޞt�Dc���.>�kX���k^�=a�JHn��Ɏ"�7=V4���a«9�♵0�
�
|��O�)�Da�C��C�D��֩�����f��A�k��f�����rA崸�!�o��8d"-���+�d�#"+��B�㌴�� �=�X�)_\t��̐a,e$?��i����d4��[#!8��(Ԭ�)Ԙȼ���,X�/����V]�Cdl�3I�č=�ϡ��_?���c��VXo/�Q|��9c=�C���q�[����S����KI<��T�5CȦ�$�d/�4>�����F1�ee[u�D �8K_����������p¾��*�ǽkͯc(��)�H���(F�F✶<*!0U�f|Z�{N��]�i�U�e�#*� ���2)v�w�-�;�O�X��KH���e�ө	���UI��d/g�w��l�[KR�o�h~�P�:V���P�L���$@�9�Y?���u�l��x^KF�w ���I'��Zn�pʈ��p�%����Q�D��F>�8�rhI֦�E0�"?��\��]*�XS�rL@��/�{B��T����6~�ف�������U}ȄY�M*�f7DNHĕqw6O���a{~��'~?��6(��.c��B���F:�Q^	�L99��!牁Gs����I���T�}�ŋ���r8F�_��8�uq!�4Bj�A7�T��������<P�[�)�o�����ո{���G5�j�FJe��tr�e�W�
M!��F�l ��l�y)�E�@p'���j<�kѦ�Z�����������]�X��h#!�$1ot>tw�W2����yba�Wx)
j����$�ǅb�K)9;�����+$�OK���{�<n5�9X{�TQ+�x'sn]��"}�V�IO63�R�{:_�g���/5�Β�cł�r=SYGa��4�<����h�x�<}�`O��:�m�.��b�1�z�E�\�i����#pT�*�,��2�[�$$AaV`�W!���B�=����������r0MR���jN�wĞ��}s�܆��P��E��ɗ��i@�W�!��^h���V}�U��#DC*I@q��b��'����[fI���qCZ�fUϛH��d��@�4�p ak�6��_L��o�r᳠�U������e���IO)%!5�^/����XH�|97�����P{�� ���pw0}Q!���Kd(w�-~\t�[A�E3n��d>�~���Y��T��R��G�Yp�ţz�]j�$�p��4}�$.GK�{���2z]��;��-��v�Ls��� JK�N�N���ӟ�5N�W�Ԧ�w�g�~ �%I���5����q��ZC��G�G!_�kn�J�Ye�=��+����F�gh!������T��H�N6�+�;�'�E��@��
A�͝5k���:�� ?Q_4ֵ�+�'`�� Xzŀ�^?J����1�\��\|_�K� ������/��1pwmt��X>�Z��H7��)���& 0�]ݥi��w��S��0 �.|�׊��^�aN%���(�5��8���bt��~=Ho�̪�	n���BfT��C�WK�*�M<զ�p0��/8{�掻�d�-#�#��a������ ��&�#�@`RoO@�}�-��G�l�]�r��1�(D�������-��f�05Ē�H��|mW�6{�^�p`�LK�`8�p&Qf2���B�Jj�E��13=��)�POi>2/�ï_�CUk��'=�e�Ĵ�ĸf�i�	�I�� �]�� ���zI�y����VA�(m���ï�x�Q��O��s�}��8Ͳ��A�@DVJpܵ��56�Jl9�%R�X������c�}�C5���ʹ�<O%eC��z�!VG��+\B>4��¨���a�=��qo�����Έ%�O5vH<{�?��H9��k����?M1�8y �q ����u�'�߽P��n���}IЈ��Ù�Yn�Ș2��Kf�Ai��=�D�8Q&ߒ$�������7��bw�ڒy/T�dz
�B���-�'�l:���B-�E�ʵvOo�	sȫϡ�]���W��|�g�Sb�r ��߯�c�V�גɄ�@�b�%�>�X�`H��\B��TF�jt)��ـ8��t?:�3���Uˆcm3Y�������6� ���E��2���ґ�8����D�]�no�k���=�AJu��a�l��{¡�4����@��E2�
5SS�;�D��g+П<'�Z�@Po��i�ޝ��Zg-C��!���|nҁP�G�ZT��BK��ȃ��@Yj�B��M��享���9�+��PA
�QT��9:=��c�#3��W��vyN���XQl��K���A��ZǺ8�`'���njbG�����g���h3�N`����+�::�ܰ"���	V���n��F����8�#-�����0�f��6Rt�[\}����{�gQY�Y�Dj�I6몁�C[CD��罡֠�#��0T�W��J;H(�O�]b
z��F����`��T����=�mn���J,X�N�l���Z��ΐxXt�MV��E��p�!^1�{��<��M���F�K��L�AkT�� F� v�����#0���}&��E9���?�4l��P=E4{���]V���]پ�J�-��.&!���x��/p��	� ,63Hs��<cQg�9���Z0

��?����|A V+�j��;�/ يx.Qqˠ���e�+�p_��h0�+2k>�������1��~�9X�rkpT_q[Yɖ�585���zZu�aPw�q��R߻`����
q��v�x��2���x�i�'x�!z�w����i��Crk�OrK.m�G��jCN$����}�����0��I�N�̈����"��O����̧3�/�V^	��aw�N�&����%�[���m�7҂攬���f^��za������˷P��[#��~ ����\Ʌe�	y�8����t�p�W��9>\E�:⤒��C�B�*>H�ݛ"z���j�G�\ۖb��Ny���";Ja;C,�:"�ĕed.��S-�xm�d�/��E��T�x��&�u�[�0��g2��j�FI����P����Ӄ��B��W�8���ǪG�4p�SJ&F���&?V�X�3:��Z�S��H7B2���#�%n+DhwOI0d0Y<f��i�
������-��ߝ��oQӓFԀ�|�����mb�3��>s�"�3�{����%l��E��D�+��ߩ���Z25>���b�L� �p�m�j�=B��ȪL1:(]s�`~����Ύd�����k�5�|F@�0fM-�Q�Ne"h��lV\��m���Q�u7C��"
4��q�1�����^�Ÿ/O�M���G�-��3X]3Ž����$�J�Kk��~�ߧ� 7Ia���M��,�'��h�㼅�P7��@}P�������`�I���ѼϤ�x=�&�*6��ŵ;)Z�^J��)n='��Rg�
�����y,Ԙ�T���
�UͶT��r���>z�gl�~�Gq䭐O'P� �-�޼����]�	]�;���r��πŝ��_����-�b��,t�aK¥���n� -��Оb�w���� ?�`��a/�F&�����k�*�iO(�	@ᬪ��h����S�趋b(c�=M��U�����sN>�U/R8�|ܠtBs����<T͋PJ����#}�?�k�qy\-7}������g�F�����|珸�Ii��%u����� 8����A�53�@�<�b��0��O�W��l*�f��{o"���S�z|�Y<C~><�=L��9�B)��n.�l]���.t�zOR;��
�T�����˪���v�������~�t�`fM�{N
�L|<-�Y�x3�_��H���ޅ�ni�XMi���40z������̽��5�>��d��V�I߲�73x�O�]�j?��wd��P��{���E�:�S_�m�#BH2Ҏ<4P�]���5�Pb͟_X-��#85<����b��'�pd̪�Fp�T6z�z�Cpd�cw�CV���Ѱ�s�qO�)�m۝�/���o�ڷ�zƇu����Π���{W�T�����|��'ɲ�\ILƣ�f��ǁC�^�)��X��p�u��G�m�q�)�7B5cF���I�w��]�ς�Y?ŧ��ŵi��A�Pd�X��L�O��:��j��"�f�8.׸3���yc��D�U ���^>���h��y(L��Ǐ��܌DAȝ+����@��RT/_Q.<<�R�1��B��3ͫA}ȱ/��!:��hg��vW�ڼ+	����ԐRDjl��d>�*������
؋��~v����V,�&�2�E	�*�':z(��Bg)��{���,�X�e�Q3���X� sey�*�"$\��M��U��c�e$-��]��Y����^&�R��j(U`N��9���߷�ig�zetHӏ��F���|���H-o��T�5�4�I�oU�W��;#BH�����j�J�ؼ�L����ӯS�U���7��\<k��
1�m' (0�Y��͚�=��"�D�f��7�߈�?�i�dS�.�7h�o�alu]|��κ���#�1>����h&V�woQ;��rU��� ���괥 q�لl{*�/P��;ַ���ױ�x�9T�N�ΎOH]w~��q(��L�AP���~�A���}Pz��UBޅ\���3���V,�Tz̈O���ce��߽L���k):�-a�e��#6¦���>�Uߛj�������݃.�xFn�̫�l=jD��vSE<�c�jA�oْ�<����&�ME{�b������oOk^$��:� ����'ˡ��Q�W|�Dx��9��m��5��+���ټ�t-���r�n.�-v����0f��"�׊�*^���^�r4V8�G]<ɧ��X$�+��UCBzV�r
'ןr�]��C�:lܷ��􌹎�'%j�,Z����m���[V]�(٫7���y�FdI6�v��}
Ȍ�b�p���G��p5�45�-��e6�zCNR�����k��-��v|���Ѽ�D����1�r���Z���pI�Y��TO��թ���M��%�1��H��\�qSVH�#��#k��k��,ָ�Y�]}iE'd�
�
Ǟ/�2ڀLc��K6�P��%�M&�?jI���
Ų:A.�����=��>J�c�Jk�WWW��f�����AS`T��`��b*�>������]L�����̧\E����8�5�*�.#"���g�	�����e��$A��Υ� ��f@��"Q��aZ^�;��,���i���ݡA�!'oVk{l�؁����4�d"��6�%��	$�m��pTu��.!��t���b��+�^�'[�4�g�P����B\ZٴMj�29�OS���	�l��(pTۢz�'�S��_S�ݠ�)2B�Z��u�f�>��.iͬ&���fC3��uz���� g[E�n1Uk{��B^�q�`-��;�c��{ �ֶ�i�Q�:-P9M�4_;A�i��4�b�u���:H�AHͱ��1��i3�ac3>ɗq<}KJQ�}#� �'l)ė���4T������k��<A��&��÷��bU�����Q)�ɝ�T�?��!ߍ8Xݎ��ex�� �I��#��e��߻��ƗW��]�9�$UF�e�it���͊Q��8���=5p�9N�(�&�� ���Ci��ub��/Cֱ�|������~���E�
]m�������m�Cc���Z�������ΗKaqi��������B�Q~s�%�+�8YQ�#�F�x`���ň�j.nw ���� ��_K���_�h�+�� �.���(��j.�m��Yz*�x3��:�l��$�J��_�ݺ<$w��$��w��Ƥ���tz�qO��[�^�M�T��rɐ����l�JE�X�r���!F��ΐť����T�= �0o�"T@�5:�٭��0���@N��`�-�y�ɛc;�
t�:�LVC�y ���R8t`��`�O7�� �'��0�1�EAz�q'��砠���R������1���V�G���[T�TKK�Ϝ3I�A2n�Е�#�uSgo��b��y6kSBuB���3�ũ�%���<m>?���{4�}��G��C|B���P����@;$J8<)�>(����`�l�r'x�:Z6�]����8lc�ڞ�V��C���Q]�hL��d�د��`��H\�;����i�o�>�v��Q�n���7�����~nQ�5���_�_:u;(��O��+�r����߅���(�H'V�#;?�נ��e;���)ۿĝ�gp�"!��'���i�[Z�Hb��Z��g�{��k8b�V nd:�dT�3F߈���\oI��p��D�����,ik�A�Y��Á�m�	�;�����r����%W����*#��1n������m��^��������<����J�Erc7��E�-��Gv~q������&.we�DE�$�
� m�O;1�E��v,�d�S-+��݊]�]T�S/K�\wGM��U��V��>jɨn�ڟ��������u)����N�=��tR��R:����#�)�W���?y�)-��K�T?������Θ5#J$��UA%�3��8�{dZՙ.�T�!`i�"�1z����z>��}�5��	S/e����OsWPt����08
 �M�䚤�C�v�z�L�Z#�T�s#���h��Ji"$X���/�JxW�ן�]Bq�p��p9�fҩ�L�����T,���W۾��o{1~�\�ɓt�:���0��@ta�^esaO�R�T�Tn�Î�S԰��x��z��b�U�iee��Y]���R���H�P*2~�=䒖ʸ�շ�D��U��%HS�ՈH���h��e�Q�W��-UnGa	qG�9�ҕ��a����W���#im�QfY�5}���J��������og*XfZJА�+�Z��ٲM����a��S^�C�͢�{�l�֡���=���>�)��s�1��Z�jF�K�vW���`��x'-�{��T�G6u�c���g�)�C��C5Ts�g�"�
�c`�u`�H�*��` AX�\�^˽ �&:�Ѿ_d���0Z���z���������Ӣ�آ iZ����}r�"Q7+a�	��
�)���$��%	iK;�펭$m��q%��K��
�M�q{?x(<oDD0N|+������wS��"d�ku�ь��Y��T��%W;��h��X�R%j�EL�Cry�̓���Gy�G^�k��T'��s4}�gG+O
��lK]��ҋ	0���ͷ-��д��.��������m+Zl>ՉpѠ�S0̜�ؐ��������G<e�q!��%��kSe,�s�ԓ�Pj�F=;9��H���P�
���C�jUR��[Ǘ lm �~d���XoX�!A9	8�p��eQ/=3k��UgIU�M�U��M���F�j ��\��Vbq��,~�*� ~��<t�>���w�����.��+l&,)�m��'��S~�C
�r��� 9O��6I� ��7�M#�C���Z�2�g�.+R1in�X��#���z["��'w���;����&=WF�>�����ca)�˻d�q2��V
w�e:Þċy�rrH��T��+��/%�NrOD &�"��n�
�Z�H#�1�D2�P.*8Z�I"�~�6���Ⱥ#a��&|y����L�ڣ�`�TC&;�6I� �;Aꐼ́����_�m]����=g��UN{|PH�A�90�No���V��\���z.����|���'{e�q�n��l�r@��W��� K��j�z�B��^���;E �����<W�a�_3����������vX.tq+�7�I[�r�j�Dє���ex��Ŭ�'�bB��#)��>w��}����e&���ۘ�f��������X�Z�����yh�N��(�2�=�[�
�a��+�`,[\��˟�q�@u���%�j�[j�F5��*�.��'�V?���X��/rc\�$�|��6�腳���<E�&"wԣWw0��Mvl�L!�����<�	���X��;�+NT:f�7��Qr���FK�*����+e�ڟ���N�5	Ti�aB�$��|��OJ����&�ۋ8����o�BA�z�p�%�1��T���uW�$�z�x'ݚO*�Ъ}k[�v��5����{S�2m�ӵN|�G���=R	8=�*�.��wB��J��c6���t���9-.ts�{#۬�(R+1�TR[&+�b��_@T)�K���'i|T��.���L�T�`o���g�;�;5�͕�/�1ԣ_mMo�v69��*iw+|��$���<=H��a\��}�K`smK��s��F�d_�B!�Ԧi�u��d�mہ�"+p4�^E��G8i���$�������[� D��o���\�`mЗ��WЍG `��k Z�7���*Xm�:jkٵ�uZ�"�_<� s5������bzl`c"�*�V�/�dˮ"�߱ۿ�Ɩ����V���yQ�o�&ã�	��ߚZ�7d6@7ĲLж��H�HvN�M@w�r�K�;��}�>N-X�F�Ò'vh=!���P
�#{�q�B�pp���7�ç�U�n��i��L�xަ-�O��Y�Y}�$�F�pᗯ?N}�ȉ�E	�<���8���Xyl��C�c��1�h�з���g�x�L�]G���@G��o�u���pLm��"#��\MU��E���8%A@z:���
�/yL�{���7)�I120Ci=*6w�t"a�rs3�~,�+��F��%�%f>�!�jP���v(8�R_Ņ85�%�)g���E �F2C��<,�A=-Cj�s�Ȑ!������&�8���k_7�TW
��-d{����2�̍�f��Y�W8��1�\
�0�|cw�O0�X�[�ܢ�&�.YC��<�aH�w��j�[)I?����ԐR��[?�=�d �!��Zw�J���gyk�ɩ�qq�[�l��L�zH�;�Ħ�����W��['�q��=���&��+���+�s1iศ6�|(�6�Tȍ`	�;�L+���L��Q:�AL��ʠgge׎��]5������_�>5V`�]��6K��H�7�6kBN	�*xe{��Jw�vz�ƴJ))(�i/N���ۢ�`Ό� DJ�{u	��&�G��n�e��=*ý��j{�Io>u��DG��>`_Xć�9Y. ���i�]���z�[��٣��4[�"�����₆:/IpО�>r�K�P�9)@���Ñ�pX���5� ��	���9 �\@뱪�l-�FZ��yHD~���<=N�4��Nh���&u��\�"�����ϸ�k2�̍�f������]<P/FH_���0 ��+���C��u^
���\x<�2Α9��\.���S$����!�N����_ �둰E�a#h��m�]*���H
T�:Q�D���d�WּE�s�+`�ilr�ѝ��������H%rľW
>T���$��f�����~��d#�d.ˈ��_�	厙�9�kc=�.Gݽr�O$\��Jk��rz�D�E� �Lz�4�z�¿����iCAs��ArA�/���P���o�$�,���FiEk��?��YS��@�źc"!dY4cة6�T��V�Ty��l�ڑ�Bx�tYi�M8^C�X�cK�^�9���@��ݻ��sN��{�G�ڍ�	$�|1g>IcY&l��,U
����(CK/}z��!���O�G��s
)Ђ���+�UWP��_cؠ3�W�}��v��kU�����M��>!�����ͭ���$"�����-�l~�<���f�"�j����
��To~�X8��@��6�i^k�O�L�iݷ/[�z�#v��Z���I���o�M@!�|!�1=ջ7�{!{�K7�
�����/Wd/#��>(N���4���I�(�y^�S	����I����`J4[�{��d���G�P��\�U�$W�]� �PҠ����8f����GsjGLih��KČ�+����R��:�\��K���Ci�<�5I�B���١h�rA����q�jCV�e�z�1�u��\��;-A;���Xp*���^��W�mb0Y)�B{&r@�6��wo�4�X�9i������n��vw����D\o�-'�T\↬��"�X�;j�&��9�� �Қ�l�_H=L�ih��t/����_�6��wo�;�
8���N��.ܯ�to'5�>�l{8L�4��u��ϯ�/^��IӺ�mN=շ�����E��h�b(^�p�;���&���1D������Y�z��6_V/�'�Q��M;8P�ʇ�]3��Կ5��q�>�.�������aI�3}��V��$��t$>H�R���Bk��yk�xì���{ɪ�4��Wwh��Fl$ԫ��2���[�q�2rTcdB���"k�� �&ӎE��\��ܪ/�ܼ߭M|���RP�)�@Y������҂An�L,o���t����aI�a���mbFH:^��h�MQ�z#Gů��o�;m�PI?)<�1����#�|-8Pd�=�ሣ���-�e�ʔ9������J�R�8#|�NY�Q���@���P~���b��u�:�-���n�G�A�����e	�y��t�|�l��*�w1����_��I:�]¸����&���N�`�/�`c�=ݓL���>��
 �j��R���u �%���m�#�+�B��B4�	��3˂�c�n���[��;� ��mM��8�)LC��Y�tg�A���Pa�=;��G����𞞹D �kXt1������6����{��І
vx����1�˿u\/'�f\ODU7(Z*�B_E���fj�[v<�Uf]F���+#ST N���r���H��xr�����>�WH޻nr��]xD�W~ԑ:V��8T�Ko�C��!e�]!�Kq���z��.����^<}�	�FflR�n�58�n�
�(^S�y�Ue�|�"m�<�N0�o|��v�29��c�45NܾF�)M��	���c�T�s��Z���+���W:���P�U�P�$�]0����X��ʸeŞ9�_��E`Y����J9^��=�u�� .��,��_�Rʎ;�
����Sk��ǔ�>v�{v���`�5��q���c7��`v9ǯ<\Qv�*�;�n��!����J���s�L���}Ĺ��
�t��3�Q�I�����V`��-�%�|���]\�BW.�<x�:��cs��a2)7Q<����Cn��$#@RU�A8��%1�[a1$�0��y����u/���x-r��I
ЂȘ#o��1��-kF������m�P���m�RK�A��hX�0����w;PDED�}�X��̛��O����QՁ�'6O�HؕBd�H��x5'���_ O*�U��/d��!-��R�g`�HP�`��u=��F>�ώ2��»��5���C�- �J��ň�������9e�2����u|%,\I�]P��l�?��ԗŬA,���2덅{
�g{殖���� }n*���Ԡ\m{[�w=��!�3�����(�<{̹z�}J��y���_���"�>��?�ʵ��cm��P\6���u��5P6�3��]�1g�~��:��,�E��=|T3�W������tw�\hy<+d�.&!f��a�r��|$��¯��7�%�;���%C�y����o�U�G�����D�r���DF�l�;���	LF�M�坟Xα�_���E޴p�|
����� ��rT} �m;/F�1���@ P`���{Sw��e^������*"UY"ܽ��RR�UN\�WvQ���	�iL�aR�?yA)Åi�&��!��)��I]�w5�.�6��R�V�?��H���	�	c%ܒڟ��2lv�:)�U�{�ڎ�A�ſ3��������y�c���]f���6d.,�*���sz>��Q��i��1C��eGF�)��9J0*m�w�l�Or�L_6	b^x(��,���0)�>VoȤ	ĥ9��¿)IW�|'���=���0
c:>��1�=��qKk�	
��L\�@��⎷�����N�Jz�25	:G�M�Ku�@��K�Ճ��]���*%˟κ�Jƙ��/�V!�L�Abu,�Dye)��r�-��fߑ�Ɩ����0�v��&��h�M�"=w0J93�
���vf	��8z�o��M�&���Z5袍2]��D[.���vچX���t�$�e�E�R�[��X���ɧ��o�CD�D��	�=�=6��jr���)��K=��������Z���>���1c�t>"^T�����r?�	�E�!)�X}G�)���2�ax����W�Mn�?o�N\W8��(%<x�9�d5/��aH�d�1�,e��gE~�q�%2�ٵg,B��x��~�0�Љ�i����z�������r2Q�=#�E ���J`,F��3��B�����{K�q
���;`��u{d||Z��j�9Y��߼GFp�sI��v�1��#���%��0Y�{C���S�G[��k�?�Go� >��Ղ�yu�磼2��W�j���`�7�K�<;�oj}:��b]������|,�/M�@ Ƀ��lX����c�0��>n��H)S�|���U��M�����V�H��aO���g�<9�Vߥ%�Kҹ�!p1����|�^���IIbGG6�T�N�dr%=���A��n�=|���Ҋ�m�o9�h'�1���3� �`��Y�HI���g�ao��,?gG��yc9�e�a���
�bZ��**�;�  `$:���[٭�Cx��6�'i�gH���5$l1	U�o��]8�r���_�m�r�\\W�1ئ���x��vԗ�u�����)Q��t���1�{������v�L�H�N1�,�����D�f��HLd��G¿�<�������t[��G�r4�H���W��#�	 ��5p��jmy�3^!J;[;�d��X	wv-I��n�H������S��>����|��3}_�ʉ�ou:�Z���dU;���,����魸8KT�)���b(���4���ܴ=�d���W���G��Y�n4��
��M�=A}�7M��<�L�ֵ}��+#U��J���qTm�����qk�w���M�Ľ��Y��o�Ӌs]_�B,ap�u�py��l</����+�ӭ���v��I3�2���U>s���+�A��Z����nzC��>c>��B���^c�����S�������B�n��^�}�B���Əf��'�R��ߟ�q
����/߇f�x�<�>�X�R��8��GZ��-� ��`zQ��ܠ����We� +>Sl�sG,$'~��!.����R��9��с��{���z�Xb	�Nx�QţJ��(��ESc3B_��Jbo=���^���6�����+����"B�r�������ᦰ{�&ɗ�?K��
t�'!�	�/݁ZS0c`p8he�^��є�U�[���fT�P5�/�h��@��P��6�����#��8��2�L��U��@�To��b�&p��8���DYK���k�%��e��A���o�K2-h�}���ӁfJ���t�T�͙�,XI\�½�}��4��H�]�A�E�l�.[r��7��͈��?��l����WHn<x�9)��:PH��\�^"i՟�������� Q���l(�q/�X�t��iΌ^ .u��hPf�-�^�����U�Q}�y7�Z���Ϫ�<��љ���,�&i�������gM��C��v)�0�����;�h|��-	 �}s�T�j���o��\g�U�J�����3��~�]�ˢӗ���ͱ��Q���S�y�'�w|���}H������<��W(��^A3Q��kn��W
�;�r�	}�|"�Uǎ$�Nm�Ϻ6�HUUTd��M<��A.q�E9fB&���@��w�,��G}�:fM�2��~��>h�aM'ļ�:.�"�=�54��ʱ���8e���~�����\�\�M�� �]4�$�V9/���XN�mQ�k,;	�$}�
��Yp��O�E��ќ 9���,y�g����SD+�
�}V	��ܠ4Z�$+����a������\y�:�eo�/�0��s�c�u��ӊ)̊H�>h��׏��j{Zb�Ny�c0���~G�]���l��Ě�?��	\����)f��A,�[nJ�e�?4A9N�AQ��p���B��%��+���HKKf|
�&t۟�G�j�V�(OZ�*���o���B���x��R*�@N��ky�/=�\������Z&^�FNG��'X��։e�q�<2�pz4�7���觩E˪=x�%��S]�Ig��R�PSpJ�J� 5����g=��� q�� c��ï����+)�����4��7f��S�M;1���ޓ�٣c�:7�b����n1��(C燣�cOB��93vP���R}k�?P����;N� �ѽ��>�bm"���q �ϣq>!w9�͡g�������P%V�j6(���.�b��C,�Hvz"�ߩ4,�ceV[mʭfFVt']�JF7�c��m\�Le䀄-���6��|T���t����q��t]b�7a�Q!+fu�bh��թ]�����U�iY($�Dᐽi�e�2���N�?�_h$���)�nW��"��S�3�=�הj�����? ВjH�9ү��ɻB2� ܰ��;fT)�������*�NQHIcx;��&�ykPƆ��nrk���Y0��<&���d	�+��U����F���=2sRg�3^��Fd���;�K�5h�FB��p\b���-�����0�"�r�s_�����{��f�86m����|$����6B�L&��������Da.<d����qhG��� }c�| �PJƘP	�OK��,�y��0��^�_[N@n��_Q�0k'A&R/��x'n��P�t�����Zҟ�!<�k����ֿLs�H'&�[��"�@A�ү�˂�k�r�1ͼ��hYpִE JjJ���".�s� ػ5��)H��m�fALD&k�\57Tp��駝?6/�IPQ~t�k(� �N<�R7'�@�]���(�6�ƬkC|�ˀ���Dؽ��G��_D�Of V�"e�R*� �>D⿑�d�1A�q�mV�n��j���}'b[9O��і�py�u�Y�X��	�����vǟ� M�⯑#���!At��-�#�=�M� E�S��E�H���|�SR%�ᅼx&�$��'m%6v,�	��m/f�j?r���+�B���e��b��>T��=3��Fj`C���)piT&<
��dE��_!�a���E]�%��c����N���&�3H�s�f9Xe��m����}���MN����}�<��V�Ac�^E��?�W�!�h��0;y%��9\�]�#tQ�?6!<��������J��ufN� ��:��'�.m�7�^yr���֚���*3P=(*�;�3�M)�6��j
}Ë
��.�T�̤b\-2 �Ne�l0C	�g��P���2�� �3�u�����'@�Y�z�X'^S&Le&�eTw�BY�̲��~b��	4�ޒ��7�y��E�Lx۴���ߑ>�0[D�SF��pwƚ6��S�5P�ͫ�f&�b�j3@�_�`h�bŹL!���>�5���J��L��젽���R�yoNs��>��$W�Ĥ�:�K0�]J<1"T��G�6�Κ��A��8k&�5�.�����M��>��X@������	��9*��D����jw�~\��#gᘡ�l0������:�m�M���vY�R�>�{^.I�|����B�Tu��	��j�+�7�R��J��BՍ�3{i�-b�oV�n�W�&�7����#�p�8���>W8�f���ȸ3D�]�KX �G A�%h����O>��\�'7*�D���KN�D����n�m�",Ύc��ֲCBc�p���8ߦ���o� ��G`��m�H���&CA&��l*~n;��[_��в��:��</���9W�v��~W���f���1�q�z�F[�U�ZȺdŚ��Ȭ�z?�)�Mib��3B��ޭ���b�Ώ��'��a��'���	k�A���\o��,�[Hf�}�x�2+��e��X/ ���2��\�wE��o9DwH$���/A��V��i�k����2���l-��?/�N��+e�,�H�����xɤ�Qx�ժ惥�;-`�gU��z� 	�K��9�yi��8����K��9��p�4�.��"R���St0E�>��%͔��x���V������
?�d)NZ�gi4n�D�8�d�jg3����jcy�k�L��!�����.��H�|��Zc�J����*;���(�;���ZK;/sp�c��^&
k���U�;���z�@��FC㝀Q'�@g��`�p�kH8}����萈�4
�f�n�"7M՛:A��IWD,��Ɂ���|s���y+~o�,h���W8��.��]��]o�O>�R\jN�/ƀ����Ď�mhV�M��B!�A�s�@GA7��.�V�ܖ ���'��s�0��R[���8Bc��Z¶8�?���D9k2�+�)�Ճ���,_S���M���6��14N�P�h+d5�Z�kz����3���>U�������]�_�6�<UzaF�%�y���'�?:�������T ���b��V��|�B>��R��c��$[�Uc#�q9�T�Q���4 >�p�g�w��v����ԁE5����	95P�ˮ0�x!�TI��; ���]�Oا�	�HlC�Iޥ�W
�Zr���@\��J��	6��.�C�d�f�YM=�6Y�ӑ�� ���Qߧ-Қ�=��q�ʤm"��H�p�V�I����[���z�P:*��l�F�{�7� ��mM�;7[�!n�����9?w��2w�<�G��рF�'��{gT���F�t�G����g�b�c&��r�L�\`Q�����w�v��bFF <�H	��d�F�����9c�{$��I� =����Lr�$�+\�]8Ճ.�(���i��E=<�Yi�� f��6�9��:�{�\mP/�
OY[�#����$��@���$�Y�7�[�=�1S�W|��WZa�����T.s�㙙��I ��W��;�?Lzm"��̝����q���T��*�MɬD%t�!�ޱqyr�P\��x|])o�l	����(r�����iHt���p��2�'ѥM��%P��H�c�z�ם����A��k�F.9;f�B�̉�3)bdr�@��\c�3�Ch[���^�����΢������D�)>&��ƛEJ�.�Q��3v�l�R5�w�E��%W��i����A��-?f�/11�_D|oL�����V����t�	^F�xg!o�A���DM�v�6��wܲs\a3�}�p�r�<q��0=������M�	v��S��xQ�Џ�����vGM���~�v7�tM�v�b�c�vkr�dGո��[�4M�5���'I��c����iw��;����ҠC�mӖ�&fj$l�ݦ$u�@�F�U4sB�V't��Q��[X~l� �E�Y��b|���ѩ���7�8��J"��yA.�X5c���`�:�%�� ^W{X�7#��\u��s���=��8�I)�, ��ʈ�f�Hͨ,��5���c��`�$� �`��TN8��zh��}V�m���)�@fV�S�J�u� ���X5 �1��#���p�ԑ��]*���-����x_
J�48�Z�"����C�~��ã:l�����D�ӎ�|��Wjg;df��9a�񱃝5���s1'����� I�9Kk�fn�!_��ؽ��f*��Pmj�`Y��(��V��'c�n����J'}�H��c6Y�wr�1\>�<��C���elg�Y�����~B�湻��>�a�T��W�e�0qO$G%�
SJ6��C���sHYĀ��TM��x���tNXQ^s\M�����mj���+�lO@�*�\�,W%�r�hċ��ά�9(��1|�M�J�����j𹫬CQ#�~��qS@��T,�'D�V,��QV�!n����ѿ�Y�1�8�%�w�:0������}��B[��G����b��3r�`c�&I��Z��Ta1��Q��f�&�;;Z�}C ��v��%/
����.-&F���o{'EC���٣�7?�*k���#\�sa1���<𯵭؈oe팩F3D9��������6Rq-Yv���SE�LD$>Y�+H*%��EZ�X�n�F�G�p����G��B���)�TP�Eiʱ	5U:��~!ԣ��VP阪�h�����84e����|Vr��+*Bb��`پ�̝���);�6�.'M�fϤ���u������gI�Ts�p*;�Α�������Y��Q������.b��Cns��e�X��u�����>����� n;�� ���?���lE�k��ΰ3A��J�t���-Cg�δ�1Hŏ�,�Nv�����{����>���z���zW��5�N۴͌�᪄S$I��-��q����|�	a���1r^�X����y�ft|yxU�%D41ܖƂ:�[��Z���Q�+�J��@��:�\��.��5]ה���#��� ��乹��p0*�_�����3��-��>�$9�i�PS&|�Zo�w׍�������*8���D'//c��(L 5Zx���}a5gc��AD�����CZ���RB�+�Qz��n�j��1�`� �C��Ɗ!�-��(p+���!���G����a:ʑc�|����[�"�¼��RJzʩe\���T����<�$=
���YI�>r��/t�����]z.�+�&<'���l��w:��6������־����S�w��	]a�T��m�c�v����d=w���ڥޮhF���{���t+M8px t"M
s�"Ж�%z@���Q�i�ϊ]�r
��ަ[\h��^C�#
��x1���4P�b�R[�޳R4\:���7�S�kef����w�E�� ߰��Kт��:�������ȺsT����ƍ7�kp�;��u�8��A����M�� YF��_Dt�خu����`F�;g��I�;�_�b�P
U|*I��k7��r+�o8�S�V�]��-��#�9�#��ɑ�6|K"Mx����P�.$G�Np?,�]9��R��bm���o�KJH0�"��q��1j�09P�iNښ�cYh��gR^�����FO� C���p�A�G\b �����)��M�I������?(���[��dE`rnteщ��C�Lܢ`��y��;&H��$;F�#���<(��U��qd�kk�aά��;����!�G�m#+�ܗ"�VM�n�*[���2�pb�����2)�g]�YJ��β��'�O�$%�l5z�pv�l�
�)<9(�1�J?��2cn<��JG���q�z�k�Q �a�F.b�����#��@���#}��T]�7�i;.`ϭ��:%��m�g5�|mP�-��$H�f0�J"Q&5ɏ�� �P�r�)ܛY��E��	[����pP%|��VT�u}��s��7�p�RR���$� �z'�[Z��_�g�b���'Czy�p��(W}�B�Y���3�O$��NVS���krQdk�D���ٷ���j��ލI���Kń�����+>�_'�*K��#������P{�
}Os��r*2� �y�0׍GH��|�4������[{xh\�˿�&�z���H��pQK:μ<ƛ�'�)�	N� M�4X8�FΈi��ν�&(ۢ�._����Z/{�u|����t'�������i[���o]����aNo'��/h�,�����d��zz���;6o��b��I�:�wH03�4�����GI˃�=Ѓ��)�W��(�}�	���p�%�9�sL{=�y����Ŏ"��{t�Z�H���ev��N)���OxqW� ��z ���c�=�}�����mDύ����Cb��C~���>���¶�Jr>�,�g/￮�P��&_��dwx{�o���������>o#梮�-���(gޕ��oM��z�å�i�nh��ǧ��_f:@�m�D�[;��	�E0j`3v����c�J�mo߄�s�z�[qi	��N���?�V�c�OZ��ap	L3�-f�3ȴE:>�X��:��.E�(a^军�҃_��+#��\"}� _�CH�u�� ��7�i�ǽ0n�Qh�wt{�ϩ���0cr�e��M��~�/�П׹�p�-��b@^��< ��i.�֐@�v��;��~�.Р� ����=��c_���L]�Y�����lZ�����J��A�J���&�Gj1����Nr���8�1��{�KIdi!�4��E�����{��:p��d5�rJW٠�z�.{V�����^`$)�Z�m^����-H�ڟ4��i�1��%\����<��6��\��ITSq2��,}�&���)#J
��$n;[��Y�ғ�ʃ^U�qHm� �
���B��r*h����Q�7C�JN�;���
�z�)�6:x������eg��iMv/ /]�c �ޕ�y����yA����B/|������%{Z��+�wܒ���髊�9��[ڠ%\K�9�;��B4��1���o��ص���Mr��ڲ�]�჋[�����fH��z�@R4	�4�lrcn�h��"z��_�]�rqo��I�W<5��$[bp��I���.VN��X����C�IV�V����<�^��hdt5�A�l� ��f)���q�"{�v�����'�=��F_��:�cn�Gw����<
������9e'p(׶a����A������K��V8��a�P�pԎ��꾕e��>�1�n�a:l/�f"}��2g17O��e[s��klD�ҤL����K_(���m�J��bЮb�pϋ�R�:�B�)lΌ���	&!;wJ�����=%��]�K!����('��L���J_4*���L����f��>�y�ʈ��(�1���Dt�{b����f���s"2	��:�J^ص�Ҩ;�Fb�t�~΃���&qh��"T7��\�Љ��}՝y'韁m�tFz���}��0eavjS��K�t/�2mRR�=���ޢ̺~�A4�os�I�%����¹w5G��R��6���z~
�P�q��tJ/�������@Wv��x7�1m��x�+��uj(y��-�q��ױ3%B:�zP
|΋��A�z�ݬ6�	��a��B��i���Qo6Z�πQ���(EOT��̺3*��+�#z��i�n��� '�@G��t�X��8!�[G�+�y��]7VN�S�i���sDcm��dg�H�[�B�×� �Dyw+ � ��ޤ�I�1�IkA.��g�y��x���^���h�*�$�j
�}-)����$B�j�����҂f���=ïK.��B�"�Gl�Zz���.I)�^�Od�qrD.�cG�m��"� ��y�'E+dM��$j&+p\�9���c�U):�4*!J)'o�[�k�XR4�u���� ���s��^�w"~�bd�n����K��k����g��}6C��e�ί�:r�c�d:�f'\����5�:� G�r=�R��*����.���7�i$����Qa۷�f��=(��j����͗{�����W�!S)��2"�o�苸@��P��� egf��G���?�sR2}�F7)�>�Ų �W�Q�j���O5����+O��/���S�,Jzc��<��yV�˪�ֹ|F1��9.:+�f�A  ��t%@��,U��:#ijd��,��UL5��Y�~L�L�-�*ٸF�a�'d���X�H��w��.[�嵻JH-.�9O!��xVj�+�QZ�U}�, ��,���9��/'�Mk��@�;��@���Y_a��PgP)��$��n=$��1� �e��B����v\�����~�Ǹ��F;��N��@3�s	D� "X ��A'��5#�(�Fǫ���V��+��:~̀ 딧��z>��-V|��3�.|6��s/� �pQ�2�Ȣ�tU�?s��_!։_}f"��w�ڈ�B���	���ˑg_��q?z�lQ�i�~F��ǆ�!��KtU.���$�a|ی;%��	��2ۋy�=���i��� �7�\����b�����'�J�<�=��O���`de��� ��-�y��ɝ*�������G�|x�J���H���.<u���ٔ��`�2��F���	ǵP�5�/���B��b�zB*����+�G4(E^j��*��D�2�Ř�)��PQ&V0{�~��hLj�֡�$I4�y�>�p��Ԩ����jy1����[L+�nd@��Ѷ��Pe�T�(���VtD��|H$�dI��):Sz&�!����K0n?��"�!�ifݎ����|o���i��A�g��z�jA��Y������s4酫90�7��H�(J �Z��hF��(*�W-F�h�%&-�,DI�|Y�,y
��f7mKP0�/N�1y��'�n.�62LZ+u2�泴g^	[���FK�5vht�סG������j'^�T�����>��{X3�}�rI�f�K� �ɗ*fu�9x����E��&��f�g�����B��*�3D=.ZO@���=�گZ�*���"�5̽*otׄ\������9��\�����*�(��#ow�2�����t��3o;l0[�=XX�ɿ`v�R�"��=�i�y�QJ�@����VR�>s��})s6�1�lC@U��	�3��lm�u�Z�]L�+�qƷ32��wѓ�!�)��u��XR�	����n�o	��k.ã�W�
��ۚ�Dn�^ó����}�U�����i��r )�bV�_�]�
�u;��Pb�}��,`�"f)�睱G����_��G���q$#4YxS8��:����)ܧ�d|���Ɨf��|�"��}�(z�rѰ�������aa~�5A� �Iu�CM]�~T^�L�Ӹ���Bn]�/�9뽉ٱor��3�F����On+o��4���:�v�\�6�N��FС��j�8��=��rW!�EE���Ut,�������Y���j{n���V��Q�m{ƨh�# ����g���+{�
g$���L5=�0�E�E�S�U�-n���o"Y�-̧ġ�k�Ҷh�	=��+շ�����%� ��'�K>��?��;|�ҟ.�Ս��/�<4�#�o¸�����[���"?����5�&S%��~Od/�������J\����.�/g�v�+����8+��-�����F�1���;PP�_l$�󧪠[�g M���U����B�V��B"q�k�I�j! ��zp"6&��F���t���8�p(�E5�g8��U�$�d���%�r����8�J��=��ꍁ�%�	�Z�i��{ ��"��zIq3ϸ-:�8�d2�@�ԫ~# 'zb�ܨ�qK0r��JѨ��X�D���D�wɂ���Y(ܺ�����}8S�"�������HPc7ep���ʸ��6��6�ׄ(�i����H`-{`�(���swA�֔�8Dz�@ N��(j �������~#�x�}�I���%��q�nrP��9��iv�ch�WR��y�q�@����*����~�yOݺYfˇ�b�eQ��
Q:ޘh��5�߼��aq��yc���}Y���/)c������h-���ӢAu�k�e��\�M�?�FR|�5ϣ��C���?�d��\h/~��BpsY�J/�T,�4�py�t�@�-ؚ�qWǾD��^�@�/Q:�)GX�ڟ�L�����g]J�cϤ+z�6��;bRJ֒��7�vI,9��"
)���'L��ӠYB哧��)a��re�Zt�(�����s��3�������#󏛄B]�%���"ݫj�k�q�
�w��oF���<A�T��l$֬/��N��J�F��}�H���~�� a��(A;u�*Lr3A�HF&���.�9��SH=���X�$d��B�E�Ple�=faB��a~��hI�������,�?0��-�,iWv�U�$3
��}��V���\����Xկ/��i����i�v'k�U��+i�AB'!��E�cF�Ftai7�j"y�L}B�m��Ӈ 0�|��o����ī<n���b%�ӄ���x��	�����~P�:ҼXz�$��Nϟ޴֎��5���m}�✖z`��x��t-Vl��B�\��Є�s8�f'2�g$���~U�ͽ86b.���X��DJO:���ZzgK�Y(`�gNl"��2��1I؆ٷ�s�˞�L�)�S�
W{ߍ�C��9U5�w�}T0����2<&V2���At�,	P5"���|A�[%�k�]��փ%��N���E/#�����ը�0��a� _����۞��.��u�����XZ)��������=yA�&�m	TБ�1��m�י��.�m���:�ǫ�yk�FT�6�����+O����Vᏽ)M��	Ʀ��iu,y��E��N-��^�*��
[rD�~�Y*c[0$�9$�NQT�x��P�����w��t����/� m����u�ƅ���'I9�[T���M6e�����U���56��N��4�������,�r�oSJㆍzΝ����ew.L�%�g�r<b![��ʘ@����L=v��z�顳�i�0��3���Yp�;� �rA�tp��Q�#��'��/@⚄���&��a��M���E�4}@��E�t�(%�w�W��p��$`X��w%�8��L4RG'��6,u�5nU�(N"lQV�ʦF.Y�Pπ��Q��p����L��w;�a�ϩb�XM��I,Λ���7+�T��/�ׁٻ �v��2�2��x���s���A��A���vh
��7{�I�gj��Կk�gޞ�&?:�G��Jc�D�o=��k}���AF)F��r3%�u��y�91��㷝�dZ��D��@i~o;ۭ=G��.O����Y�c;~Ֆm	��O1���S}@R2g�{gq��p�Nc��5n��f.KQl�< ��a:���w�$��	A�9Lo���]�Cݑ�v`i�Y�KD��ZSGt��I���Or\чXC��\��tn�ޞ�:#(T��~[�Gu���q� Y.����=S*����f�Y.:����&=5��
g�h��qzv��Sh�K���茗�{ӈT@��j�	RzwuM���z�?4lQL�έ)�{aҏZ���Ut�/s����$���*� �c���e��cZ�lx�2*4��g(*���l?�c�e�C9>��fC4��yzC!��N�{o��=m���Ә � �n�4P�ƃ&+م����JLn{lJ����ф&��h�q��u�$
� �v�Z�230�w1i�(u�KUm����6l����e]h�� ��wh�9��'�F�wi'�q��e�4^�Ig��Sƛ����4����fe� ��-4�Z���R�.�G��S��6��҆Z`��y��]F�s u'�ɕa����)��Gq��ȱEs��[�r|,�O�91��Gg6Pڽ�����6P��6EJ�Z����?���|�(��V��#�� ���ч9#:�<8Z�$�nv��D�8)��I�]ׯ�LB}uC��Pw��̐^�Ck�n�ӎ�mx�||ߺ0����U���tĆ��9-�I�%^i�v�\�b��p��>��o����"L�
 ,oƿ��`�eG��Hc>��QN�2��V\���~4�+]����8��,������ٗ�'�2q`�{2mw��9�غ�6�^د���DI�W���C��5)�󂧄�>\��,G�yN#<��V�=�A`�V��
iPt���PY�e�H+^޹�B��C� Lq�������gՕwdL�<��;��T�T����z�n.�!�Hԕ��ڨJv�ǻ!�
ƺ�$�A���&k��/>�19�i� r�ݿ�-��q/]�y38�='4�=�0P�r9��Q��;��K��7vRe_U�������&�7���<���鴝�E1nzJI���W��+V��]P��[0��F%����8���2Dh��p�W�BԸ#�|2�Ɲ�ʎ��V��&�~�q��5,�2�om��[���C�ո�PH�{�N�yX�)�p�ᘳ���5@�� ���,��ǉ�
��XG�����>�j�J�ˁi��gN�F$�}�,{�Z���h:��T�����l�8u�i�Q(=~��zk�X\�����H��T_�kj��`���>v}7�r4�2w�]'�pj!��Y������;�R���Um*��=����v3|:�Y�eAi)b��c�pr�}��&͋�і ��[��]Pw�����qϨ��Bdif�p��n5<����Xߞ�0�ЋU�;�4q�.~�#҈Z�U�ׄ�|�l�v�fkn�VI>x��0�%O��
ʋ��Ms"9��>9��� c�G��Qa�B��Y
�E�4��v|���k�^��{�'~tG�
+N�C�@�
�/�z�	�+�`��88��]h���.8
ǯ[�$��Z>���D��t�|�����i�����y4�(�[(v��<����p�t1�o�,߅v���@��+s��a@ M�O���%s�J�}'�g��(�ͦ��q����o$�_�����"�V�s�or`�-����KX��`$D���J��x�!��!���)�6ߵ%�ݳt<)�4�V�zAj�BEF��B<wb$^n��7'Q�G�6�I\�Q�2�Gw��m0��SgТe{Q��N�epv�lTت{ؠ'-���	EJ��剥�k������H�/wɚ���U�=�)Pz��e�u�*�r�Q���ᰈ]FpA�q��\���������>ᔎVn�	ܡ�>Ƚ9��J{�ڦ�q�r�m��H���j���W@@��I�K�#
g���c���j�����옜}xvN��L_T"=B����U֍��hH�a eA]
ծC�P7�X�W�]x�4��[၉*$�>�Y��rs�\�I AϹ����}u"�^~�B�Y���i@|<t���(J�pN��| >��#D�_��Rp<�}YI^�W���ܥx�	���{ՀLg�B�pW R|����3��B�A~��%g`v����080tP �F��2ڕ�#���.Iqh�ܦ<U��W�+�]����I��A�/ŝ h�y�� ���gr�;��W�K�{קY`'�6�m0h����?��DbQ�lUZC�25B~�fn�l����=�]@m�]����e��^ż'�?.4gL��]Fm�]�5M"���Ur�y/�����܋�)�s�,:���1��TU6F]��Yt�/x�����y��Q�d��|���g�J��;xwf��*�s�n\��S0����kyЙ�H+�mg��� �R����2J�c���k�.t��gz§ 3^���K�R�"zD's��j��7
�7�8��.����o'ܩ�9�P���#7%9$�v���'�<��N��l�ȏ�����R���f����98���jPb����j�Y_1��kmNVY�w���>�lf0�a����ۏ��dk�(�!ܼ"N����/�=%,����,Z���|����0E��E�d���?�� }j��Nt	w�F���Q�V�S�_Ԉ�K��f��-�]�IjA<)���x�*��иb����Y	�5�Z+#F�xC��Rp�~Z`t��qZ��r��Ω�C�bܟ/&�g�,,N�!S��v��0]7)me�=l񁵼�d#��/�S3$�m德:�o��<T���s
�W�U�'���2&p�P	�k���r�FMcYӥ�p�1x���ޏ��2E�pJ��)���;(byS��e��Ц�l]$ٙn���7vf�ꥹv/��t':�e�:�(��$Ֆ�'Ƴs��1�3�A�7-�ײ�,q'T!� ,T?�i���s�Ҭ�P]|�d�����|Ƌ^=}��чH�'�uH�&�}��1���ƥ�b�`:�``7@�)�TE�U1�� ��<�l�:M,�� �覣m�1���A)������O�.�����7�WL	G&�tS6�vN��Hש�"!6g8�k�*���Y���1��ʥDbz8x����m���'��DB�[�i�-���tU���6�l�`�~��h���[�75HN2��O*���U�6�[���6�c~m=X�o�׍N�.F�"�����EY���9��iаY��z��$
����dG�����q7u��{k�Ԍ��/�Gb
�ev9NY������ٕ��5r_r�P���k�B냯ɶl�۲2>-:��L�~�����}|Q�x|�]�X^���PY� o��Ƞ���BV��2m����,����{��
k�ӵN���1ܞ�푚/���e�]kf��i)w���'x2h����pT
�Nq�c� aR������}Nڽ{�m�ߒNb����1�]OGcw[ѫ������2g� ����uK�-#rZ��3�"g͎�.��;��ͰI����c��x�AGc�����G��W������*��^�elL�^o�򰅨Ac�T[G�[I�l���N57�-E�[�:7�o��\dp�wy��UQvv3��q�"��h�F]�v�R�h�%�>�����6��/�<��ƹ�-�nS�c:)�~w�$����`���8�9-��ˤHm7���SNAy����_:��x{�0�;o-${2��o�I��k�đ1��r�D�;�1�+���qN�|������&şG/ȌBv���w���sft\D�h��/8���t'�[i#����Hj�������7D��Q�E��]q/+>��7ߑC^�=ۆ��#�bS�ηI�(�[|����R���/溸'��%{W�� P�ӌ�2�b{��m��s���;L�Pl���%�=��F�Mi*u+�IV�5��iB*?�5��KE&5. ��!Z��k��~���H�o��;��L�F�S��R���g!��0�[�KJ�0��Pڐ�Gm[��)M�
3��l8Xa�6��Cð'�4^�r���<�8+_(�e��4�R��Њ	�m('��q˹��a����넼�L��[ I����M
1�R�F,9F؝�m=�y�ƚC~�_Wf���Y����y)�����ժۚR�1�A�ng%��,��n���|j���*��Ч}|b`dR{.�t�+l���1��	����>��bJ��I����4�� ����O�6+�����q[ɱ��G��T�Yˍ(�g��b��?v�c~DO�;��5m�ɴb�)<"U{b����z�v�bǒ,�XK��i�G��q#��Ú�n���d6ac��ڛN�B��:?�[� �yGj�d/�%X�u�3��l$����of�D�7|�B����?�$�׶�-�z蜦�Dؘ�@�ɂ���|�-�>�B��\���z�臝%?Ͷ�Ղ�9��0���>ñ��-4�G�|�KiW����$%=�����[�~˜��[�H����X�Ȕ� �[��cE��8�!�G(��ߠz����bQ@դclOem��USr��5|b�ɋ��Yf�A6�ؼ�^X��Z)�9`��\��y3�n�+����$��L��	�)p$�D�f����ف0d���NЪ�>��_�+
2��r��ֹ���>����V�1N��n9o�Zk��s��$I�聗�-.,��C��q�'���?/\4k��U�P�N�C޸H���qc�ܙ}�4%��Z�������7��!ª�r�,bq��k�زב|�䅽��-&�� 4�����~G�������[ɰٺ�I��,�Iu)?id֪�n~��c'5��S���x=Ywt�`�v�$�T���V��l��۰ ��i�d*��~l�W�3�V�q��`�\�}/1��$�D�%��rv�Yޞ��*A�i��Z���5�����U �V��8�bȇ�xZ2Ib~��jz�Wt9��Uezr>�e?��1�LE�=��>��T �H��lA���/�B�]�9���������]����1���-��������>���H˞q�:r��!�V���ǰB*�W�tT,��/��\Eɢ����"��LW����9�3M|d�Mx
Ĵ����?�?��1�f݁�*aS0e�d��׎�;�܈�62�AJ���ΨO�e.I��=�=��̉�y�/��w�-�f�X=��=��jΚ
 �"xJ��'#Q/��4�ԉG�`��T��*^�X2��K���/ �0o��O+��M$a���$&ו�^5g.�ON����VO�j�-�o�w�}��/���a��$q�~�A�\����=;�sǳjD���6pˈ���5�۞��Z�K�b��b�(��Χ� ɕ�coI�G;��[`�&���1Mϔ�W�?4*���"?�H��{巋;�&%�(���L�thځ#<�"u��l~��V���S?	��Ĺ�~�5��ZB�A���k�lr������cҿ�����A+��L�<r'�A!�.�Θt�,�l7�}��/0�,�:l��Fwz�Q���lR13eШ��nn8�hb{��4���[&�� J��*|�@P�5�_L�,m�	e�����SUl&Dnx�Mĸh�`"5�����S/4V䋖��n���nW?e[��FK�7�il��T��_��D}J0�++��8ъ��Ԡ��_�ZWqۖC(p�bd������u,���X^A[�yd����3��/��y˸�S:O�f9�20_�u{�;ё`"��&犊��0��4�~���m�8B�Z���eٷ��r�;���Σ=b��*�۾���0#P�|
С��K20���B?�r�&�'�T�c��}QDy�R=��W�d7KE�k1���ܒXiyQz��{�I��Y�>����
�� �<��Q%���׈����������](�r�q��d/B�k��)'��(BY���4"�n�a���ρ���O{.U��yH�yF�t�;"�`���eL>*�����p�%����M�Lj�p>��˝�U|��
�����/�-�������#җ�û���i?�����9��%�F�)�����oa�T�d�ĝ`}����ip{<"q��(�V���V��T��l�o�A�?��S�l9s�EY����%���k��i�Ұ%�C�}�3�4-�y:M�4� 1T�㘅�n�в��9�Q�laUe�ɪX^��m�����@d��P�x��W��(��?a�ül��ԋ��M7��4�����I��~�r��T��Wk��PS�8�/�,��uz�7��,ֿ�ƻw�������׶`f�{���s�Pܔ��sj�8��?|��<��l;��g�����0�+�_�W�Lb�� ƕg�
� g�/H������x@�7&��'�t��{Re9�F������YS[��]�K\A���	�x
�p�U�u�C<`��%��bN��'#u��\dӟ��J)T0��˽a�ᒆ2ߴ��#��#�`��U���&�pkV���7�\fNɮ�]�Q�x�����=H~�O>g�j����-�ҘFT�ˠ��^��2�j�bas�_?�`�u�� C*���8l�1zҟ	R��������P���M�x(�}�'�ES�|�?�#�l�C���2Fy�	q_Pp�~�4�6Ix�]���8���rL�=��E>n�(��:<�RaC�\n�<��}� <���,NR����VZ?|��&sY����Ff��R�v�i-�V	����k5���a%�x)eF���+��ku;NK;,_�
���tsg��M	�[����B��R�:�!kǋk^a.s���MWU#t�a	g�R�HYؖ�UUΓ�s^%A�8�IwF�� }_����LQ�'bj� ;+t"��V>5IF�|���:S���v9ZNʹ�'������/]�5�=Iʺ�����]zG:��A�&��)��v��i+�D���  ���y�l1�߄�����4N�,�B�s;l@�Q���J)	{�?�b����?|�i��h1~Zʎ4Q�%�L�c�_%..fpgP���>j�
��.� ���>�l�`�F���4tg�v5�E�pQ�Jx��w&M<�Z|�v��G"l%o0��`�=o"N_u&��p��+�]&�+�͑ZOA���D��Ĥ6��8�UH{p��\�Ņ�]`4��̃�-��Gjb��ˉ��X�f��tS�J�����s']H�bhͽ���N��Uza̹�	
v;�\8����{��-OXMq}�طÅ���w$�n�U��-"����Y ;�}d���;Cfran)�)7A�mI�>U�If~,'�e��auޜ���IȅՂ�PO�A H���sYD!e��j>��S0�����wr�`k�F���A[�J��������ߑ��E�Ŏ�f�bWR�1|p粻 0^���L�L�Y���A���B�7�I�}k~�_H�ʁ�9���,k$6��%�O��I%ݷ:	H~6�٤v�˫�I�l�i���h3/�ߡ_.�d�9�0��p���L`aD|y��h|0�R%A��e$N{g7;I��*I�=w�]�~��ߥ��1�Pg�)c8����(-��m�����4A �N�ȐO�߮�!�C*������{x0|�Pa�]�����EH�W*�{�Z�����̭#1���
�l$d��i�v؆�?eHF�Z��Tv^����ދ��b�l�!���s\6�cHeJU����dY�H%��2���Ǝ`x]K�:fm= S���`_3�bsHY�bn㠒�2s\�r���
=�K���]&?�pO��G����;��k�l8�EG`� I�,π��@�E8������U��A�<�~;��B-�"xR��K�*Qi��q�(8�{�{=�r�` rU�N�c���=���N�<ݔ4x~>wH쒹k�;
i&��"l��*�u�I�L�e�<Iw�b��r��u�p ��0'��;F/�V�T\&8UȰ}�ɮR!YbU��B�K���کM�>�� ,p�(]"4���СK>	����`���Fn<�/	V���.]bq����)`}�p�Gŭ+�g��
�{��މ��w��G�~�Pk�О:�7Oź�m,��iծ��Ya�.���5���
Y�	y���C\3]��j�'��4&00�QJ�gr���	�_��h�@��6�e����i��_�9æ9��U����c���]��_�_!������Ȋ�K���f{+���s��x��V��t�����+����0���c1x��@�-ȝ�[:���bo�V�A$�D�;�e.���̬�菱��&�'�8hl����#���פ$�gp��ً�J�_^��0*h -��|q���������~V��	�����,�7����y�r	�5,wEp�ș�/���Ʃ����3'oΥ����|8�7"r6��x�rT5��T!0���<�(o�_��;2��L�zz��
��_CY�wN9o�D����^@�3��y�W�qt�Ϻɝ_�o��K8ŗ����/�b&m��D)��
8�� ZZb~i�4��*[k>)\�\_�r5Z�tW�c���68�d���>�߭U����w�|�=z�-=Ԑ魻��b��	lt���6�	����F��yU<�F���}��R�'����qWVyqQ�SJ���5���'�k�&�ְ��Z����0�ǵ��O<��W<S��ƹX���pR��K�9�k�-�.B�x��f�lu��G.��Ol��܅���U1�鳚Q{~��H;DSi;SK�ya��q�6�����f��O��q����ID�C�]8�0�>М޽d5�	�u���	0�5j���i<���j�	W��F��b�j��?{xa��r_��H��T�@�:h=�0Kl:��^H���}�!�45x	�G2{��qt���'�:##�Ġ\#��B=�#dDD��ECԃZ�>�#��4�Ê��bGv��&H*�!8��%����\Ͳ�l���!��W��kX���M?��r�+ԞR��O���`y+s��0�ʒ�e��i���c9�ܽ*N�x�zvF��aa!�^��4:�Y
���V�:����җ-��{o��sA/��慀5�}Uvr�f�u��OP����>t�h_*�QY�O` ��T^���;>qfi >S�p��{S��P?�.nf%���!�^���� ^Y�c��Df?���U��M���t��u��Z����h����?��L)@��\C���� ���Ԓ��PU����;��F5��og��k��oZ.o�A��5��^�^,T���;�ܳ�*�`�'م����Ҟ�6~��� Ӭ��Mix�p�!;��,��I��XŁ=p��j6:&��l�b�]��>r�<>A�y�w*:�]���H�S]���u;eG��� �Fl�֡��Ó���=�君7@�f����zs%�X��J(��}�e��m�"��7�M����c�nܻ9r�]L�� ��0��g-ҡ�HI\���D��"�o4��$:��c;&.UJ��	P��6����c���$06<Ȼ�?��Cv�r�� �_9��"���+eWA��c��3�,�P��x��g��+�T�䊉�
�Ft*����Y$?fp(�RiFT`��ZMT�T�ʭ�U�Ѕ�uN^�U��_��I�iWZE��s���x�Pp>;mc���()���:B�z�c&"������x�=�`ěF�7'.�x҈�C�J������H�ՀlR[4ׁ�u�DM�X�՝%���t`��
K��Tg@�s��yO�S�\ޙ���#���f|1���gE��cv~!��^�U`3S��"�@��8A;|d��*ջD����_�ސ얚K�4�w�!����j���hISǛ3� T֗��s�,�=uW@���)�HĞ�ض���Q��r�G5�C=�+�Yt�zў�;ŨMϺ�к����b�A:�����#�+�y�c�N��ut�P5�1�E[�>X$�Zw0�`y$��P�A����1�/Զ��X�@8�閦�<ŗ{/d����S�Xt�~��)$"=1�|m��r�k�G���1�UAsō�*%����yU����]Ʊ)ڽ������v��*_���c?Ce0��m��H��L)F����+��{���?̽u|�EE�Y2�����ݩ�E2�f{�޽�CW��Iݘv<;�5DH�u�5��TI���kWL���1[4gHK�SrKsj�Cf�i�#֊~�m�D�l4����`T�x��u�8,�RBe���7.��Q�g�t̓��k�Q�c����K����_���bbSY��a<8✧V_<x��F���~M�ʛ���cVX�!h�5ل�c��D����F_�R��I�q^���_�BaR~�O�M��{~�`Z�����!��5g��Q��hFB�R������ڼW}^�Os�s���C�y/L��cA��dR�N>��Yv�t�?']�;8O�:�<j#S���]���V+.[]�!��Ϟ��;�k매2W�.�u/d� ~�yܰp�-F�"]�^�mK�G�FN��MI�3KcƼev�
��!)�����7$#>)�<ׂ�*R��e���YL7X�^K`&?�v�[����v����0�#�����U�	���(6Z�V{Ѷ��_���s��]�jo�К��`��L�Y=�	���5�GO8�(��e���}�:�H:��h´�+�(9*�ѯdbX��; 빎�D�B��� ���7��֧����<}��!g*��DW�.�.G}��!K��M�97�!�������_B:0G�>Ӂ�����1�0�ғd�|2iSe��÷��et�&.Ɵ�}o#J�}?s�ͥ��[��ӟ��E������nA�M`�����+}��!:��3PO��p�2a/FPWR� �:��_iq�j.ml|`�����J� �y���ƏO!�	^;��f��3�'��O��6�=�8*��(<kf�2ȱyhd�U ��C�w�*����A�1��麼
_4����= �����S�5��fy�,�BD-
L�/J�Ɨq	�;�ǭ̱��D�ڜD�m#0�!��P�8b]k��R��7^��0l����m-#�_��;f��	�w+���b݄Ĩ�rtt��X���T��9�K��]��ݯ�sD)b$>Pf���о�I��s�[xUl;�����A�����m^n���d�2�����(JoM���Ma���R��l0B�;�9�8ʀp�C�KWO8�gU��w�pDT��L�φjr�z�Io���=�M�o�,���\ot�|�~"=�Ш@Þ,�C���
IS��l���c�1u?��|̕�+it�,42H�W��XfXY2�d~��8�J b35;_os=�� �N�kf��A�׳@����M;�Gܭ�'t�-��͆q�̗	�&QR<(et������{�O$��K#-�V �����BaI��!��2 �>Z;&�� -C�*�-��.�9l�!��+*�EE�ըpnӃ��K�5%Mq/��0*�J�m
���0K׶Mhfq�����A����JbO�oE���ۿV�o��(KׯJv')���%E���[j�_Mc���k�;���I���M��\��Ҭ{(��Wh��_Ubܬ�J)�S��ɽ0YwЖ {Yȧ�J�
��}�!�pͳ�rO�/�K('���g��{��V8AfG��KS�d�������e�rR�mӺ!mO���x�ci��jޣ��-��A�iF�)7Ռ"&r��X,6*#�I���IkxI�o+9Y	!q�94P�6+9X��e,X�V��Rgt)E/�<s`)Ȓ������S9t
�|�:�j���&�N���J;�F?QY�W�\���/�rj]c�N�,��*<
�[���(1�X:�6�z��+���*��#�:N�N@�"�y�u� �^��.$G��!T�+�5��x�����Q���J1_��<^I+�wE�ʳ���Q�d�L<[g����]{ר��u��^V���c	0�V˓��	�Mh�gu�1��������I��]6�j�
�C[�����j=���o$U��XJ�A�W� ���)w��^F@Wܒ��m��w<usw��]�-�/I�+�	E#�/��y�j(j��9�,5���Ϊ�տ+�)[eu��E�	�h��,�F^���n�"��+�4���D3���9����a�Ɩ��$E�Z�!<�H^�Nt�Z�����E��<�pg3�J�4���A��2,��
1{֌`�����}�CA���8�'ͪI/���d�ύ
}��%Ҧ�Ld�9�H��4|�����	��C��뛸�iv�E���fV�VF�0��ڽYFS�HC�9g���� �[��@�8�>�So̸�a��,�?C���F6Z��M��nM�^a�y'/��3S�N#,�Cd������X�o(z�GH�]�����#Y���(�l��p��Zj�诔�� �����N��l���E�v�0q�jf�<�@��We?�	���.�+��s^5Dv��2-�yb��r�y�m:eJ�H=�Vi�ә����~�yG�CvCأL2[����͗�K֐I#J�Fara4I�<�zo�VG�kxƃ��fde�P��;M�#+v�է��6ڤ�&�cO������A�%�<��b��w��_�AX�w�P�� �~�&`ˢ�����g��s8���?868����|w��)�]>@VBYhV>1.w��]krSK$<z-?���a�
`刈5Ij�"��Wk8O��ڦA��a�*L��3t��"/�ǖ�r.����F�G�9�s�	`6)_w�'攦��ۡL�v�L�ǜK�3��2ϩr��e �Ru�u�� ���k[��:*��5�EX�;\�cz5
L��;Q�!�Lxޝa��O���P�|�n���%֥6.�����s�⫟r�-�h���*�&�k+���s�������3�Rj��E/�?�ڼu���Li��`�N��i�}��@����H����"��q��!a(�0�X���&��>�����}��A	S?�y�3<yH	!7�@l��#|��J�����o�Xl�8p1�歫���6��ˬ߭0w鴭yA�;Z�G�,����["�U���ث��V�������0I��yp�����Y=�8���f�q���ܤc�� Ec�`0���J�h����G���;�^�R���Fu7����$�G��k-�5N�|�)�Q;ЗRش����X����/R�Zj��ǣN2�^e.����V�{���'�)���a�A`��p@u���8ӏ��b�SaQ�iYy�`���R��T֤���k�;�n>��0A��c�P��/���S%�ӡ����8��*�HEr#����ת,ɸ�
=2D��<��*����dv�T7� NAd��T��P������@�S��G��X���&�h2?z��i҄$����M���9̮�s�3l�S;�>o��)�L��Ffq�[��e��B���I]¡+e�p�n��8e_��4#ҧSX���'%\��g�A��f�v�Y��zC�$��6O(/��_M�,�/�ia%�/��u��!�Ce�D�|����{�c�6xUO����'O�g����4_���EI8|�:S�2�ES���j^>
@cK��x���)���D�;���A0�.�B����m�諭�䜚b��>27�ZC�@>�d�Κ� �Fm���J�
�
b���;�����B	T>��ͨ?�+}BX6���M2�O�P[p�c�$�%|A?*�	
ܗ!�rj�,�y��������'�!�/���,s���ŀ�4��F]j��j�v�R3NU^i�Ӟz�FLh���w}�-�&�x�{8 ���,��Vo���m:�K��I&!���%ݥ�x�������������B�^@����L����K���SJ���"�[�Ov�NW\���)>�]x�FM�b賤��=^q��xDĘ�a/>f���1����i&u�`����5�z�%�f��y�$rΨ��6N����vK���-��5y }���D�2k's	���y���]��_	���w:{e����yY�/�MN�@��S�nO% ��&j|����XH�;��0w�A�Κ����5RDBqq�Ņ�.�[�e�[�����0�:ۦ�����`Df�Ǘ尿�~a�����~�P�,��-���-$� h7)	�2F�(�X��߿�{iVHV��$|ل�UkC3�� ���HР�Ǖ����t�6׎N	"���:��?iI+�hǷ{��j
5��Z���|u�����P�W�284/|&_#��)D	�;�1��n-ý���X �p#�c��G���-��7Kԭ��_1N	aX�W����=LY��ctɦ��Y�#��IJ�7)�j��:c��q�W~,�ьު~�o����e���,�@���X�m��]B�pPi0��G���ƅ.�ɘ��vW������柰66v&��$)uY��a��ƉKf�6§��ع9Ky�Y����v'C�ޑY{a8k+��"~�+�t����fu:���jz4%�����;������5�k���������c/�p�gk�Ud���^�\�=�v<w��[9�2/���-QGG�f6Z(��`�
ǀ����@5~�P;ݍŐ�ki׭��i��+���]4A�Uұd`��U}>�Kw�$�#���r�6�8 �X�4_������e`����U�B`��� �ڑ:Bj{`�S�_�^�3D��Ѣ4$���I�OhZ������֘ɟ�Δr��PƐ��i~{X��|��&�F-�/A:|XWW�T�L��q��)C��'�#h��������11���*u>_�rJb+&��i�R`�Z>��Gp�y��Չ�j F�|t;&��0�N��kXG�%��z����®�}�t4~�Pj$A$c ŭ0�)�{+g�p���9 �cUp�2��>s�"hc?�65=�?�qK9�C�]m`���᧺���X���&�&����x�CC�}�Y��Ǌڌ��.�p!H���!�</�1���1���9^���E|#{sV�RM��v9��Jt3dBJ�K 2�7�S�ýX�7�0[��r�^�gFu�Z�(j?��_�.�_�%�I�E�;7&�=��r�	�z��H���C�+�g��h>l?��G��ʞ��!�O4���7<��^���h��6ye;r^ý���_i�Q���EŇp�>I���3B�>I̤䵒��
?��{c:�T&vy�	�o�IE��C-� �=X� (���T�0���`U�d�"9��H���	���o���閱�ߠBMߘ�L��Eϻ�na�i�y�n]���G|5�/�n:=�����[�]��Z~Tv3y���3�������wOM�
�-;��Dk�tݽ��W�YY�8�M�;J�֕ѹ���Hx��ȕ��sp���[my�+_��?<$��b
��΃j����e&:�}�x>��}�BC���Ԓ'4!������s�ڝ�(f��g_��m2�Q;��i�|7f�Ύ:SK��n0"$ ��`i��
�F� G5B>n��'�}��	d���|������p�>�OK��Ax�9ʭ�-�"զ҇O�F���?�q����a�~���e��A�����cA�M�G*�g"l���	�AN�G�]�A��{��$3�TD�c��ܚd����_S������q#b��|߿sv5����6����m8$�.홂/&wu�k��hV.g��6�������^�)[_�nYL5׶!�����m�E@�좖��AU���s���\+ok�q��EY�m�^���NⰌ�m,6�b�Cȅ�4��U[�.���{\�>�`]��[s��%�h��]ņ��M�ۺf_���:�U���1<�X�cj�ZJE�x1���R�&������0iV�s4�=S:�FQ}b����\hu��H�g�1���fx��)|��p��HL�)�SoYK�'� "5�;�W�<uv.�g���������O�=ϝl�����c�O6��cUz&3���%����K�	�!�߸an��Ӝk�]��j�I��4(A�\I`�4���Q¬Ş����Z��eP�9�1ැL���V
������i��@��t��l�#r �u#+�����X�2m&�
�7�qZ�w���ΆB�_�%�w*		#pA��e� �g�E��F��}�M�|!�9�7��`ϋ��&����QV�&��S���� ��1��r�J"	ݫG�j�?�Z��]��O��﻾�u6{�)u*��O�!����1����Ws�����m'Y��\�ޣ���o��w�C�_�畹�v�N^��DSa�?V��,dC��<��35I��X�^q�P	7d�?��6��PϽ�'�(�ˑ��9-*ϭ�(�fo��4�1��e{$������6�L���2�̠�����F"Y.�Gx�k ��x�6t���	W�F4��h3s����+--���&��7��G����Ŵ�ӭ�%L ����^UĒ������Tj�3s���H�����tU�7�To�E��G�.�j6��o�o�k�E�s���?�B���X	�W^���o�h�e��xa�L���P������CLe��	��߶}�'�(w��U8ԓ�1������ �[�zZ��s�3�"��*R�̈́��G�a�.Xq���R���+�u�Πwݶl���g�o��������jKk��5�aw��OK�ؗf�� �fwm����)cS��NM5�������(�e
��Bg&��c�?Rg�Q)�a�U>��mo%�C�~+���mk���/��HjȲ����6IZ�V��sr�
�Ӽ4������~�o���}�Y��v��s��~� j�j��·;~�o�˖ �@�C�$�0�a ��~9;b �,��;׶/D�.xj��ٕBZ7Pܝ�*��.J��77��f�5�v���ee�Ycu�X��1�(��?��4��2�@ܯ�C�<�*�/���gr�^L�.��8�+/̺f؝Wq�Q�-x��0�$QTʻ���C�V5�Q9�	���	����u����o���/��������0Y��~�b9��-��=�u�2�W�������j>�.�D����#�s`��-����mi4��||������8c���7�b�*yj����t-����;^�P��y��^�u�N�bp��:Ɵ2��ǒ3�5�L/�7`�����D!.j��`��~V���!#���υ�g�5�^�N_�Ok��z�f��MQ<ęã�����@�hh/�zn�D��ܛ}���(�脁>�o�Eע�N�����[�p<2�������P(GC�+�Nѝ�1��8��U���z=�-/dtF�#��J��VSV��3��٣/�1�7���N.CJD=TNc�]yW&Fҥb^3dқR�JA�2L������׌T�Ȋ�+.l��b��Gw�X�}�&fB��lE1y���t�V"�.P�Q��m:�PG6�g���zw�&*`�,7� ���<8��$����r�zqlO�gE�^��VS�n��ɼ�)0@9�$�|'�iM�H���Su`p��s_>{t]��)U7�����ܺ=	���yo�F��u?�2�1�,EE�ʶ��Z�ƚǥ�7��Q4*%lB�`&;q+�/}Ds���Dk*m�����k� ;oQ8
R�9�Y[��y��op�3e�yo���0S���s��y�ųez�C� 洍��`����Ӵ��b�,���u|Gg���J=X��y���hE�#�6H��ft�|��b���¶���g;�7̏���]���ܤ���C���zvI���u��x������S�V�EI�/:9N�PAH���H���P־�vx5��}@��7iw�B��y��ې��pQ�T�F�<n��`o<*��������	��N����Z�������r%J+�փ#d�m��7>`R�����&am���״�1���T���b�f���F�[�_Am��f�o��I�U��e���k�-]�;��]^;� ����{@��j)�d�GcW�i7"���k�d˶�V��릱]�Ĕ'niU}�j�s�t��kş"˟�Iѧ����dtxg����(�v�~�3j~Ni�RE_�_�U��/8��#��E��p#�O+Ҡ���1#��*0{(_D*����b��9��>1:�Z� ���5Q����A�u���V���ӗ�,r[M��}'=8�U�"�O'>!�r�ˌ������}C3��ހ/|~%`�̖w�w�zn�C+�I=����
����F�L�3������#�.y�,:$���/s�V�ueȑ�?)�
H���C�!�v}���`����|.G���9��W%�j����%UtA�@����q����t���ǅ��R/����^���h�aa�S��eWU㝏�v�klg���HM����, ��Ӫ  T½���vJ������o�
m #���.N@l� 1��STM��%@X�N�s�e%ɀ1��9��9���J�GG?���p�o��[6$�&�9�,磗2����]���VH�,�K��/���'�2��4*Zs1�09V]�@I0�'X�q�\�t*�@��h0��gP�Z����P���]x�T0��oO$v��� Gَ�g1�B���p�}�f�P���F��G�0�#�̥�Ǆޘ|��j+Tꣵ�z%%�w/��8��M�6^�}����T'�P�����%�����5l�ؒ3��ÇZ`��[����b�R�u���t����vY��_����ú}�I����I�9f`�>��kD�6��A�P�#c��Y��T)`l˿L�r_�r>-�w�$�&~?9�f�C:#�>�o����GC��r`;�i���U�hD�8�i|UCfsQ���"�\E`)�j�luA#w��3��&@U��i���Ao�p���E�J���{�M��\�#�M�E�T�Ӛ�t��K�0�
u~)8��j���R�G�����W�
o�g���]LD�Zu��帜)���w����"S�44���WzF
��౩�D.5߼���� ��Ӎ=T;��x/�7�2��/CL"�̋)�x���6#�PH	��<�ԗ:����D�.)(K�~_r��ڔ��ݕ��)��)�������)�e���,~��K�TJ�
	$3����M^W9�nr�=T��5�w�!���58y�����i9�$E�λ�W���=���8ܯ�p��'�v���Q�F[^;�]E+5�#��X�����X��u_��ڐ�>=H;Wȴ��59ĢqK��'p��J!����fZ>c��N9�R�>���F ��g�[�A�F��:���|���+�t���$#��	��5���[�Am�p�e;�L��I�����^�������@�I�~�X�@�����r���H�n��m�Ti�\a���!��q��5���=��m��Y��Lˮ]� 4�N,��&ND��hP{��7љ�b@0�y�C]&pX��8S�QA��fî�:Oyi�I���6c�H�:���*��@8;������e.W�4�L_G�4���zR���V8E�.s�m<Y�� �gh�*�Y}����F��{l�	���Z��V��!
� >��_��+P��f#f�u�<
Щ�*�0�µLi�M'�>��x�*0�;q�1�{�������
��~9����1
�:���"�J��|Ơ��if�xNO[��n�R�Ũ@(ـ��5c)p�	OoȲjf��}G4cb
�%ʘ cS���FIDm#+��w1ڎ�����W�RA��H�Z�2��"���l�F�$�e<:c���d�Q �r ��ɟ䞑�Y�b�~fJ{�����}Zrh(V��Ƌ���L�p����R��$x��cR ; ��'��#Ícx�-��6;%O����],CvW�z/d<��mذ%G�u9�La޼l9
�k�����3�<��Y�~���E��K��9'f���#J��/��"/%�*:�^C�#Z��ǼG�x�� �C�STˁ�!�o%zʁ�@����5v�i=��c�l}p�Y�=�o�\�i�n�V_��M5�>��o�SZ��IH����+��T�ޟh���OO_`�Od���dI;�ћO�;�?d�H����@qۋSr���8��NBjK�3�f,G&��9�Cjw�qҴ�xz������-z�fs��H�doeՊE���؞ #��GXҀ��g��������Z����2J0Ⱦ���c49z��Rݓ(�����������#��t3��- :���)��|��?�,��{y�O*&	�D�/�X#�|Y�?��x�{M��ԇ%�es�l�����Յs$	"?�=��3t��U��t:�V$������t��_�l���o/E�����
J��z�Ӏ�Ӡ�[2�=zj3��xnS�c��V�\ג���,rd�y �U���tZ�׏lY���2�k���Yw	����z�1"�pD�?L#7�e4���G}b�6X0����Gb%�k��a�@�,�?�g��h�u�^+y~�2d>�������1��Ye[&���]�	WAs4�O��1[��J�l,��u�_z�~�����Ui�8��7��0/��u+L�@A��vG�͂2Y��T5��?����yfZS��܂,���ׁz�9�1�\w�3����`?�τ0y=�m���-{d����΃mZM���+9su��=����&��6*a���۫/�GhG�ً7������C���|7K!�T���&��b�b�\Ϳ�Gp_.��C�lC�Y�w���ݣN���	�别�d�>�wE[�8��5%섐5�i�|��KB���iĢd^��4钃TM� �)�S�r�R"��oU�^8<s��Fr�qoX�e�Y<4�!��s9G��B<�1���kl�3��I���eK�p�W�����[��=��4`��L�9ؒϒ(�c�(�wԳ1�3�Ƞ?C@�4���Dg{����z�f�3;�0��p����b�����1�lxH02�>|}��i�9���MAcK�ٓ�o��4Jr�7KT�%�~�;-oL�̂�Y��E��Y7�~|�a�]��x�z�ߦ�yy������n�M�PemD��9$��,�Š ?��\!g�#�X�y���|f7���b��N�G �	Y�}m�f���������J��$��l��^:W���5��xC��w���+��5+�!&��|�**Eۭ$A���IA����޲A��s��-n%�(�c�m̑:�"k�,n�ΏyH��7gx.�-���ܝ�����}/R����"T8D�B0^���B�5����K�lψG����Ɖ�������yX��Lw.D���*�|@�k
��8���ݎ�ZI���y��p8Q�ŵ]&�Q�
�u���I2wJ�2���W�1���E'�M�N��.:�H��DE9�Pl��z��HAJ��L� 5~�۱K�������lcF�o��j�P��vkEϫ��BT�ty�(�N[9;M�"���<Lm� ��B%�_��.[6�E/��m�R�m2-�s��`�D5��̆��Z#_�L��t�(�c;����_Q�  ~3�ث\zI,:���T�jA@5PO������#����,�ȑ�&����_��L>K��6�0�� ��+ר$�fFOK����0����7���_�+V�OC�[�T�v�d����<�;���4]dF���~��_����x��$�>i}��	���ͷ��7��r1�g��eT��p-]�y}��)m��S�(q�Q1�يF1���.�S�:d�&P[�z��+eW��@�#җ"���Z�*�u�v�Gz�ȑ������W
��C��P@�T��.򫗻S��߸	��9����������F�k�
�B��;'����rz�R(��Neo���+B�8V?}�U�ffE�h��S �x�v�����@�D8�##�
Cj6<���#^4�&]t�/z�V�a)k����[��*i�hB����KG���'��@�/YmkAX�4��&�N�Nŷ��'���'~��L�cq��Q��1�`M�t}���븯Z�H�lhA�A�o�k2��|o^u�s��	��Ui��A�(e�pg��}���T���6jkoy,��}BnV��3��_�2��?f{l[���]�Ƙ��M�A�ȱ:�4��E���(J�TR��-�4�`�pe�~�҇�V�$�0fJ[�� �3?��fѫ���{�"�A��&����-:H������!qXm��"��1C%���E�_)F���2X*A�����<f������α��v:��x������\V���č\�Z�&gvgE�:������K�vh%�Ź��H?ȧ�4�RPx<��|�Ŕ���g>p�S��{W"�zH�^�5�Öho縀s��ot����xӬ)~N�"�wJ��2I{z��y���M�E��k,�AQ�ڶ�����)��*���4�nUo��U����џOr�O�~���#��{hza�r�&Z��^������?� t��_�?=������_�8���ö�i�_��k�tU�m�|�󘐤���+p����+et1E���E��1<�����Y�03�)6DM���;��Bo?��q�x�1I��k�*��1g0VEoH��:�	�w�"�ա���s�W�S�?𛏰�� e��U���w��[���Uq5�z���.�r��Ww)Y%x�K����Vjl�ɽ��XBH;���$�$�
��+�����C��M"
�5���=�>BN��RrDL]5%&rxn|"�}�|͉☯RS��%��"��� B�ؼ��j�*V�h�&R��V��.f�E��˼��;�Pt&>���ꞩ�=8K�j-E֪�h�
��p(��P�_�juY#��o[Z��zi�J�	��i7H7bt ���u�L��O��g�}��~�0zn-'~my��[��5:������FI��7*+��໾'ʼoU�X�"![��?�@�Di�V>��A���Z0��y7
��Z+�J^�ɣ���B���� F71�	Ӝi������?C��Kd�b���L�d�x��#\iH��!M��0����+�L�Mc��i�Cկ�)A� ��;�oƪ�đ?{���[��%*����k�R����w�yAK�̕-�2�P�I�ߩ.����Oݕ9�KbM����3� ~��O�^@�<��x�^�xi%}
閉�s<�sT3_������>��uL�bF)���tO�P���P<�n�C�Z�t�3+�j?�#���0Zm��r�(�$=�䞆[��q��1DU�h+c�p�����?G���`եU��`��Y-=
�p��)�+҅��P�R����$miR���W�+x`�$F�f�i�O܁�r���KSV=x؜񦴾2+�^m�;�IofחK`� �D2>���q$nO����)Y�_�{;2���)&�cS�ݤ�~��)k��j!�U[�9�X�I�����^���EI@�����+����XiqH[���}��v�V4d���m��/"!Z����p=��f��*	q3A�*|fa�9��G�D+ߢ��O���j��9�5�c��D�[�%��U�p�<k��J���H
�rڟ�w4�
������A���[8����b-H�����l�l� 
3w~�����τ_'�����_����.^��.\������k����.U�z-'�9��������c���GCQ��)q���̒�<[^kG��~GIM14�1��]/�'t�������qg�x��&�F�Ȕj��<��5Kđ���o�K?Y���T��c�oj��w�2����>�	aK{�3�$�A����d?����r҉�b����DEƍ:�.�Q�R��h����x`s�=$�������D��L�������k����V��(*��r�B�m�;��Ҫ0K-F)������3h+�t��B�\�SAaݽ�r�Ј~�HK�XmR��.���0�����E�8f�.�%�-�!&�l?�'� ���w!��a��k�D���8VC'_��������t�f���)%bD�&�C���$�T�q����$���v۝���=)��C�E���r�qpw&�tͮ�T|Z,��I��=�eoN翈�lspaK�l��O�ſ���N�.�cM��}
ZN��]�c�dvE��ŋ[��+���-/��B��%��� %������]�e�eٛZ��(B���
.��<� �"�PK��K%�ٸ��0#2b��h*;���x����.�z�q����kR�~Os�e��b�����j��E�3pӁ%�d&<m�9���Ս�В�;}t�r�}�|��kV~�w;~a�>C��zM�:{pB�g\}�{� ��a����_�Ǜ�%������z)]���L�8ɐ��?�kG�����\�����M�̲ƞG��c>S�2�E�1��^�+��
{�,�(�mR8lW�����F��4��b�d��a�J���:��⟁��\�^��7%Q�4��0�v����g�"�\7@9��0�ڀ�Ec0[�Zw��E �x���!��D�r�F�*`�'@�I�6��|3Ӥ�����b�g����2�I�*�������zfG��S�y�qfI�i$��^�.�~��Q8�r�l��DU{v׀��z���z~�8E�Q�k�gV�d s� �T���{]m�8�@I�r�)g�SAq_Q��*G3Jun��P������L
�Sb@�����_ �}�Kj�]�,Hm�I�kU��׻�3�r	LKܥ9:���j�i����ݘ�D�&)($K��lW�������H����]P|�s��/��}�*҃k��bM�� J��8�轫A(����M�3�|�j؂{�5�м:�I8'F�x��"��}��s#�[��z��(P#�Ÿŗ�(ps��e���6y��E#y�p����$4�xƸU�@�a�C,�(�ѨF�1rLr���1� ��F=�ԍ���^�_�gd���S�|t��I�tr8���e������]ȅR���H�����ИK2�R�5�lm�j�����Oap�G�	�}>��p�:_Muͱm��t�,xVN�D��U��M�Lf�$B�Q�ssX���[\i
�=�wqژ��d�DX����0n�v�`ܴr3u�xs*Q�ї�5-t-�b��EN%C;WH�4�S�`��ms�8]�^i���4�OG��J�o⮹߃tF���XBݨ(zjp�Z* ,!��5�xq]V3�����d�๚��[�ZY}�Nv��M8 ���j��cMIʓ�?Y2�o�T�y���]R�=��g�,#b୞h��X�4�9Kc�Ek
΍�ꡃvC�)*ڊ��H/�S�g���~s�Ǆp�) i��r��������%ymQR��(I�nk���[�Wݥ�MJ�����ov��������1�y��Y�<t|��X�J#i8��SU��U�����O�%7�k�JHUX�JԤ���B=�!,�nY���`���c+�\������T{E�)<�}�$C��?��k�O$X#�=���B�EG˕̠��:;O!w��)wa����
�腋���?���8�;,(Y�J���S7�Ιa�p? _��"���˖+p�w���ZjW'�$	������@�Q͏���V������J]!Hg�p�w��k���~sߜŉ��u%mD���^����*�Ůɡc���K�[j�uKP6P�9e���0���v�]��( �1\۹��� ���㲒l����@q]�1!��l�ޘ]�9�m�~3�3UOz��8d1
�Z��fP���ju~
����zr�-]O��=�C���ƹ�ķ6�٤g�Ti�"I�y$t��?�����A}^�!�Xҥy�����7!m�{�T*br�����JE�M����'VZ �J����;�q�ޠ��|3tI�Ȣ����z�
����r�n�	���`M�t
�.d����;d�_l`���`�j�$�qa�<�$`s޹v��/�PF{��4�����6����õL`�^�/���L�� d �,"OCD���[OS���_fC�d�l��ܯ��c�9bR`ջ`���x;��<	��^�  -K&�y�5Y��bZ;t��0��6��Y"FbO&g�$&ʂ��-u*��<'�����;Ր{P�0A�}_�}�C��H���H��7z�("���s\e�3ρ�F�92�AO�or�S��#ZY�58Й ��ov�ܺ�
��߂z�Q	X��)��A���\Ca�����L���II��~��R�6ϗF=r%�#�N�s��1 HN�棚�A�XH���!41��3�jx��>��٣U��@�lj������м������"����k>Ť�b�	���}qu���t��ץ\���,��iZ2r�X��QV�1l���!Lw��%��!?٠�ЊM�����j6�`��j$B>�l$�w�D��s�[u�(w�oj����<���#aws�9�]5�gq�w�S,T"���b���1�i�݅L6�JuWMJ�`H�����e�3WA�.�d��4�h{����T��8]�\��LUqslXX��me�g�Uc�a��7�*�K������%s*]D�-[���ipe��ߜB���ފ����.όUM�W��U��Ԅ	�{�Jg��]�'����z��~��c�M��Qɰ�D9ҧ���v򮦡;hm(�ソˇx*� Og�1ȭ��z�h)~`KE�  R�[<ݞ֨�N���;vE�Ȟ��<຅��$C�;���m7�ţ�=Thy�@�Zj��S{�]�/�O8=!�s�Ti���	��N: YG�y�к�<�BP���H��S�\��z�K���#���%���<եb���x��1�\�D���[��)R�{gAv[qqK���D�����䒙M��m�M�v%�pȚ�C�=O��Ǧ^_�������d-�Cy�r�H���;�:�q����X��o��F��!�E�f,.f�������}Fm���Q�
n>�`�W�T�s�pQ+k�1я�����!A�xf-� �N����]���f�ّ5ƻK�������T�/7H	�	�;ci���)�j��Ƥ0���ʒe�a�]p���)h@8.2L�w�D�j�Sj#>lzl�#��r�l���0�573�q-\p���M�D:�꒿�l���p�x�������<�0<�Py��`ZM~���r'Ǜ:����;���$(�:"h��LQ��v������ݨ"��F���Vؤ�l����4�\ӥE��d'�+ד�U�q�*^�w%��})��p(�[��tX�flp�l�_�����U�+�C�=��e"�x��x�h����	������.$�ې|��َaL}���L� ��5ޢ�k q'Vp��X��-1`{6-i��+z��<�%ʡD��ƾ6�J:�0���Cl�E*�y��(7�RM�l�.ެR�!Dc��_"�%y̎�C
���XE<��:��{�t��qA�F��.�U;�W{��Ĵ3͞(�hb������H#�c.�!���fzb��9��zn��s��N��A�ʃՏ�}��%�+���y������` �1v����eL#��6+��'��K��.���8}i��nVu_�B�غ�@:�l:Ü�l%j��z��\n�G�X���D紪���'�*�Q�^�W���A|Ea�AUa��L@gBeӔG)7tm�|O�z�L�	*��K�t�~��s�
��/0HMn���^���BHb�v�(}!{��Q���&,��A���$�S�3@ %����z~X�˰���5r��S�ڊ��CQ�9�$���/�eoRU���s��;]���_>�@�]c��h�L������K݅jq��˚}���;iێ�B��Y������q��z���-6�4>����`�Υo�Fٻ��7FDBN��i�	��9M4�,	$��1�!� C�G��n`tl {����oF������i�m��@<��¢^��{��8N=0�F��|���l�~
���,Y�Y �%&u}�֖��ʢ��B��g�����b�p(��I�Wִ$:n30֝}�\���i)�O�����|�l��f���!�i�,�E�}$sz,��c�mw5^凪�}�8/Np��L��Ym���c��R�����q�FN���o4ܾ-�����6�,齵u3��%o��ĩ��5s?�+)՟�R�`�Nc��F�'~ucʋ�s9B�D[��a�B5 �U�
88q'lØ�s�<�w�L����I�}?��ʕA�+aފ5ݑ�D��R::�I��TG��3044�]wzc⇘lІ2)�҄���㽟hѲgP.�G�p�z�(�ol4��9���_FH�M�7�4���o]��4߬�GL�}ė��<
9�qb��5yկ�5��v;�5�8 t]�o83��f!4��G��&J�b�C�(�R|]�5��B�b�-��k��V|-�\��������PY���L�@���_0	&�-�]�p� a<�:�e�p�:KNf��+�uWCoL[�?@t�r(�X�k��(Z���`P%�}�SE�FB���t`�����
즥<c�/��8/|��D�9eL���m�� �K|�ʒ�ꁗ�~`%uZ0ɫ���Ef��q �}f�)����&�;oL��D�{n��rn������҆��<���A��O�t��,}��qd4�v��߉�$���gfW�Uk)��M�*c�yZ/��K�@I�#��4޾�{��Ƣ�-~�J>FPH�KGXd.�����4��ʙ��}�K��mxQ$S?"$P�$�;uN��,6�jў�F��Y|��0��5M�>J�2O��3���4|�bDt����]��WI���I�z��z��v=��r�9.O��y��#���3g�r�K�[�+rh���qX�;�ZE�`�Q5�u~K�A"%3K(L�p�)J����T�]���f`����egSdZ�r�v�%)���'/���<>svU��p�BXf�Ϭ�[���T���/�y)����|l����-�e`�i��5#8��>��UVP|J��+,���G��2gЀ�eO�F��Ym�;�mꁄ�Nq�'�XU҃��G�6?�a-��dl�g[# �agF��6cRc����0ಟ�
u�mC��d��$�J�� �?��<p&+�3��SԞ��G�e���;9�'[Q�.��K�����4���U/�7�����=�,��V�#ҟ$�%jC|`^*�斥I;���7�}�z?-�
йu��r!FӀ�7l��$g~`���ȃ/�;-(1L�Pٸsv����d��t=�x~#���s��\��9�ڱqa�9�h2P�`�J���r�ΤJt�\#	Ҩ6e5��Mr��i�/B<1G�?���K_����V���3s�o��?&��ob�* ϖ��x�{ I�����,����	�|aZ�L�J�0��lg@�K�qLO��g4ppF��.�j���U;�3?E�C����'���	�6)�[h?�M?���b5ꗛ!�z�f�v���'	�<}'�
�T��K�E�c^��Xy5�8N~ȱ!"l <,я�Y�k(WY	m���å�<�R��ğM9��D����\��\��+%�O9\�}jw#kJ���rsחi3��D�f�e�`�+���[�(_�a'�r�'��Lǎ�'��c 2�C�^�bx� �.j, d�,e/��������<���)�!�J�L�}E�EZ��n��Ǿ9xx���Te�0Q&���%w{Q���:��W����@W����<��xH�������p�Չ�.��t-���Br77�d�L�e����#y;��H�Y��*m:��T��ov�����_P�T�W�o����=�g�]�'�P*X������v]�s9�]�%�X!�{������W�1��H@)z�3BqȚ_/@���hm���Q:zbX7N���}4�3��-f(tV�<�O�R�H�v��m�蚷�'c��n�f�����#6��y�R�h��%�n��4%���(����Fp�z+�<�v^��Ɩ�K��{�� �� ]�T�Ow!'�C!M���{����sE���'g%PX�\j��)��]��y�d69:� �����f��M���i��k��`�����'�О$��t|�$ȸ\�-y��Ν⥝��S����`Hw�T���[��0��/'��A��~��ob��b,�4��S��k^d�u3/3)8 q���N �ìb����3�rJZB!��xW\�~���)���w�%:�����^��������M��N�-��x;�FQ�:�F�r��{@�K
��K9��>o�|�����5"B�&#�G��j{L{�3�5��T�V�4R��˺C|�[����5��Dw=k���S���#����	MI��(Ȥ��$��ѵ�ǀ,*ɉ��gB�x u7�L�Ȅ���It��ݙ3.R�UW���S�}�j�3�m�؈�����V�˔^��L ��N]s�(�N��+ߡ���q�����V~�&�٘��Aqa���{��U��"7~U��ɮ�͞:a��d�G'-���t�j���C	+U:��76�`�c~JΖx�aXos�����ڋu���"&������.H�;V�R4�
F��А�n=_�G�����n��[�+˦jG��r[A��E1` �0����4y��1!���Z��s^1�l����O�V�5jZu���!ʁ[�!$׏�T:/��Pki��x)������>��8]#�e�4����Ԁ��b�MP�57L��ꞓ4�2�����
�j{Ly<R\�*��P��0�����c�#a�Oy�nCx�KQE@�(�]�-�g��Zj��g^����W� ��֮_,���W>Bk�T�_�cd��\\'�|�! �[�����|m��ޫ*���B]��V`Ѥ04'�L*Dk���W�)Hf�w�'H8Mvm��1�u�Ɔ�9v1c�o}x�x�q��a0� P�AG�̬�n�}�r��=�VD��"fF�6�޵[;��ϋ�GD��pAz����^������5[je2"r��Dy�d���̷�֬���d�|Ci�|CwvT��טC����"��|t��_E���~�!BK{(J�,u�e���FYo�g�uiv����p�N�3���U<!�^<h5�˗�,bP����}TV��oA4	OODY�%��;���X�������-GL3L�L�9*g�Ş�µ��P�����F@VD��ݍ� ^E�z2�=t�щ����
�i/LM��*��>��Oafj�N�N�����xd?�оn�t�b�r+7/����y��g�2n½��
iB_�j��4q5��x��$��d�9��X �/�#�,�8����[,6/�Q��3�8��j� ?��d9��Y6���~{�k�r���B[-�$:!�2.�P��_��5ȓ������=���k�t�e;[򯉠z0QŖI�ӄ�S�!��?N2���֓�n��/A���`�����(A�����nI� $sT�"��9PU5?W��-м���	o�k�ތ�u��=�"w��^f�$��S�f�άKhG���] -���F#/����\"�F�����j5�m�J#$
����^���V���S�5UQ	 ��߿�B�4j0�H�S��E���<���"n8���"R�Y~3HeyhW�]c޲V�����Ț�A��T����H(IQ���a���n�ž�ؖ�)A�$�F����8��������JϮl^h�[�)�H�;�������D����J`�>[��J��j��=�����aw��0�dx�����V�d����@��Bi�^�����,o�	d@���53�-� ����Wmٰ���HZ�T)����k��_�c-�РQG`�[�|.�r�o�(�Q[��R�=k�U��vR�\�#���:��Py?\lr_%�i��[/�c��?��*G/���t{L	w��>�LU���ˢ"��r����ļ�\Q��������)��x���+ݾ�*�`7UA���kN�5���N"�������bk��x�d�1*��<��gd�.Q�������3�b����tD��+��lG lK��%��{QfC����p+=��k�;�-ps�c9ms�#4��d���}s&��L��D�(�S��]���P}�x��37����Xh��A���x��i�W�]�\B����1`9{�d�kLk��f�̣��AUwEAR�/�d�ꔕ*4��w!���߭%���0p�@>.�s����	�\k*}�Wڳe)�v�*F�(z��P�M̮9�{�Sk`�\ҏ��`����$YM�	a�Ї���k�k��<�S���_�l�6\p ��G|����Z���0�	�ߢ���%���za�3�ݧh`�5c�l�	*�אi� JD1Pi���wShl˲���O\m�[c�%}'�j�,�!��X��%I��>�}?���:i��>G�gw2f16�����/�kF���� ���g|7@�j�z�0:�||��.�.m�-a?TI1��?�c/���Ӆ��Yѧ	2l�8��K[|)�pk1����O�)*�^�S���*�#W�v��΂��%��Mp;�m?�\�&����������1K�kAx!1����"1Ӡ��JK���//�ƽB��3Ǟ��"&H��Ȗ���N���PҚ@~SU��Ro��2�_��|��G�r���QP���辕LE
Lh��URUTeLR��&�lP:`�w4����.r)��:XQ�b�����{�O;��%*b%������P�{q�E�U�&`��T�`|� �;"/E���5�{.�հ��I;F�1���d�N�I�b����O�s�����%�����e�.����qg�N�V��=߅�������x�����~f�Κ�g0���:��PP�c�B���J�@<p��r�0�u�	�Q��Q1��΀�d���� �[T������WkѸ��V��Ɯj�v�W��Ϸ��֞Ѽp#z�m�cm�ە��s��yiUr��.{�
.���0".�����ndS�1L#���
ruN�n�� $z�M�\?�mHԸ��W���k�Im���❤����{�1I|7�E;��V؞?\� �� _iiת~B-�e����=�R�|�:��]>d� >��Jc����9BꯍA�yZ��1��/�{�$ګ����Fa P�Z6(�� mfF��� �F��fGt�PO��wE�#��l��e�$ۧ����-��NFض7_�ΎM�إ�X�.A���kR��#�qƦ�r*iDȂ��̀�c�ɶ
���K�tC�,3����ӕ�����F�A*�wZ��iS3��hip��A��bd��+��<����w�!��FS�+�҃hߚ�YTgϞ���07c��UP gu��H~�x�ws+���pXQ��s����N?�'��ѢYc6��E~�����3�(���H{��9B6��R�>�aF�fr�B��/�r�l^\����v0�����.�2����K��N�n�e����N9 ��"xH�M9n\����5ۆ:�1L�Z�~o@a�P�5��t�wFM�o�Pl�W�WB��Z\}�<��{�1:X�����=Zۅ��-b��3���o�>�t�/�➘�E��?[g\g?� S�BM������w�T���BZv���4�60��y�½[�ڟ�)Wa�6v�aH�{�ʖR2za �-8���J	\*-"���!h��Jr�'��3'$j��NR����D�X �v��_۟t���K-~*���(���ɤh3��>E�<%	%��P�_Z����J6?S0Q��z�����?�b�݊S���l��X~�Q�$�yMp U�#R[���Ni�"���։Ƌ"����Rd�c���3�x��8)��+��~a�K�������"�HN�t�M�2��:����J�&bOځ��)���:6}�C�Gn������<+���>8��?��9v�?ضhCx���z�j7:揎��]0�=`7���l��p2X��!.�0�i�t׃�e�7���ȎG���F#S=�����D7�'5�o���T�/]���I"ΔX.>���Jo��٨%��{��Zc�g�s^�,=�bǛ	ǲ2��͓8��E8��x�^c�_��O�x�8�W�\ںHwSR�|ۮ�
��X^��Q G��Ӆ1�Z��+]x6�ύJC��{�Tw�Nq}�XBp��23�I�\.�1sha���	/�2�4H뎽�Y����ؿ
��� ����	��Ɵ����� +�Y�;�ֿ	q'��[H�P�v��Z[��p�d�|��{\�\�d�I����f����
����I�6u@�Ԭ�	��LI�w����g��+�lB��H��&�j���UM�%f��e'%BY9�
�
;{��P1���t�/բ!�0�+bI��JG��4�[�G�A���@��+A�[H�������:���w�J�U|�b���Ôk�����o�|i."t�b�q@�D�v�X^�J={�9�\������T*�~����.��v��FS�2&Yծ;o�X�h��x �WwĽ����-�����`
TAP>x��� �kt���q�����eg��c�'A� Y#L�C��C���F��k#�fސ�M����&�����K�����_���|��q�W��:�E�6���`�=���+�3{b.mXlrq�h5<Aym"5?�V��&��­����;�G(�Q<�{��),� -�R�<�5�����ӁG2s��΀W����<[��:����Ac�d-�Y]%�/��E�C���ʁ�@j�$��74@�nĶ8�
i��LE�w��X���i��Y�zh]c��F;��W�E�r���\N�p�j��2|a��j�y]�1�}���n����ӭN� �����>���0W��]�Z�Xi|�� �n��T�B���Ary�4�?��!�:�DN✎���4-F� ƍ;WdF���s@�7�4FK��T��0��h
�������m����^0�#��)�H3�� ��͓߯�|
��uvv7�"x=)����p��+������n�(^�-Į;��3o�_g1Pot.*@b �_F�&0Ka�!|�p���7d*-���+��%�̈́m�LY����s�v�����jR��k�3@1S���O�}ФuAԀ��작�����j�����5]\�韹�@\����P&Wq���cr�җ���(w�]�)��F��τ��7�<��Mf��z+��k`�Փ� �(�[S:����2�s����,�6b�R��5~�V[������y>�����r���J 
�+yG�������9& �Oɞ����鬓5=���l �&@j����]C�'�L2^��x�Mw4��ʘ���TE�v]Դ���A�.5H�:<�`�r��1Ԉk�a�w�57�RkoSk���	��t˩���T�6����.��W23ZX�ۻƸ�|Cl�h����x�t���'~	��CB�d�y5z�*1�V�o �A\���I��������6�ߙ�=�u թ����H�C<������U5���aai����C��\�����#7~�������U���Zw�0�{��c���-��
 �u$�H�9�7��y [ M�����u�qXk� ׋d�C��aetމ��Fw�ܡd������@���&�k�Q���YRG�y�w�f$mX�Cjܨ��R� �i>�tiYb��h��+�.�F�)&8���4�L'U`�����Z����BO�2����F|ݾ����h�E��zբSh9�u�ǫ��`4�X6�_
�8{a�e.˶��]��(&�ԛq����_�W��j8�	#̘�`��Nz���VѠ�����)y&h[��G=�h��	'�;r�#����w��K���	�3cb��*� b��R��?���e�%By���v>�/�n��(�_Sǧ�]F
]�5�4��^ǭ��;�DOo�zhrLi�l�+��`�r4*�i�
*�=�K*����L%\�b@�V]+�ܑƲ��(�5�Y`���y7l�Qܡ4�M��\�|��UN�R��yհ�/�G�<4�$T���E�5a�RhV�c�2�H�{�r�s��&3�kv3<���s&�W��*?S�:F���U�Q��L��27����p}�A\:sIxG��<�3�k�9[Ltw�?��?.����S?j������p6�yl�}P��ҚTt�qK���3l$증!d��� �ق����f�O�D�In��Q���>l�qq!�R�� !D�z����@Flw��)[C��5����v��鰘&������ ��ۊ����-/U���A.5��A���P/nG�W7!H�a�2>����~Y疱T�&a�X�{��ĳ4���ngR��:��|�RߟZ�U�v;�s����h$/��q�����_yc�ǲ����# [�G�95�k:n+�	uE�����
r���!��I_�#�a��hq�&�A�gg T�1�z�B�*�\�#K�>u������a�h4�5	�B��`�\��.O���b���i+��q��F~�8$��W�+����$jZ���h&̂U-Ʊ�\��y )��0�&u]�]S�v��#�Ћk��-c��s��-�*��k�7A�3Y�I��y�]>'/a}92{u�R���/���R��F��� 4�D�`ff1gRN�^��ځ����BF��ʧ�r��T����4���~�Dk{t���g̙	��j3#��1��Bܝ�ޛ�C�ǤՑ�-�M�
�l�&M��nv�d2B姬���o�긪�8,���w����y��A��5���CA�
� ��(D�4�rQ̙�	8�z&`� � �w��觝��M04-�5o��S8�w-u%��}��-��a���tR������/*0���O�OʍPв����d��+eH�J}L;�-��j���]÷Ut�g{\'f�w��T@�S�V�W�ަ�.�Қ��6\J���{ �[,X�C�B:(��;���dO�����Ҙ��|��]��L: �%� �/#E{�ha��%�	�&���vmgU*F�s�\�q�[58%e�3�EϛA'��/��L\�P�gT'c2�%p}�"<|��u���h�)^c!���?Ց'_�?��A-d�W��=��#3��4�Z��T��{Sj�����h��E����>��dyxŪ���vq�~E�!Y�#�rfd��}!M���$��m�YJ>_��!��A�j�K���v��Y(��z9�<NPo��6&=� =�sڂ�Ƚ��=ΥCu�ʪ�f��%yO�(���s��u�ؕ?����8�V���,���[�$Ƴa.b�NY�T`�k�`�/(Y�`���xvye�\�r߾�+���%*�u����~u�<��X���C��Mٍ�S7�D���ǣ�O��U�E���^A�6�������}��(u+��FP�x��iW1>HJ�I#Z��ۗ�j�ju [g9듬|8��(��+ʦF�̞W����kAȔ1��7f�o�&M.>���^Vq��>�yoeoz�q�?\,�*�'�n| D��O"p�F����|��![�ɲZ�+�1�~�q��|�h�œH���䦹����%ܙ�)w��VР-��f�Xk��Q{��Y�4��������^���U���D>��6s���$~$��3�&�UQ�>|�[��aٓ����(�3���9�/�`a��:P:�בz��Ck)�ď�F�܈����3̑O�&ơ��*���	�� _QG�6���s�$��A]zR��Oó�f����A������vA�y��`������CS��A�!��C���O��3�へ��?S�`AJ�G�s��������]ͩ����?Jޞ*v�v�F�,��h)H�bՈyY�K	(T������Y��E��D�i�kR�����~9�8�[�]�NA��i��z"9U�9sμ�j�sa)_���j��2��ʐdi���\�t^�`�����G��ݯ��ͣ���ن­i�,��������<F�4槌���`�j���;è�*!ίSy��98]�k�Έ%���Y�I�A�A8�D������3o`^>�<(�]kLε,�Jo������i�����>��:�\��½~`ɕ:<�_�i��tU�Y��`��V|���:ܛ�7�c�h�e�+I�a� ?9�m�s��F�;)Fˌ��5� t'�;�je�$d�|3����z�n[��b�Q��F��l$�~qQ�+�;ڠ3ԩO��ﴼf.������]]�?���t�Y��e�S�B�e��س�ȋ9�����x���Z	͸X��	D	h9�i�3p���f{�m�4AsꞠ�,��1��d<#�~���|��� + Y[�L0&%��6m8�Gh�f>� ��y+�Y���44گ��f����]�~ <��'-�t���`�|[��:(FJ,2�.�1*	�����8q�Ѥ���9zfcC���P����(;�|Eg��j�r��d�ъ[�>6vJj+��MV���{��	:	r��g}^�%�՝1��GO��Ոr�9������4�+l�����H-z
O^p���N�wn6x_ˏ�25�SKO�Q���5���\#G��[���c�
��R�UČ������%������ �x���,�G��|y�W#�n�ꬃ<��8q�S
r�Ȗ�I���S6�*��Lj(�N�����!��D���R��T�j>��M1��.�C�%A�_g���Hz��c�$J�'�yd˅-=u��S�����P1�RP�?v��?+����po��s�C���ta�f3=�]}R����a¡�p��τp*|4$�ۛ�s̅ �ь*"Oy��\��\v��.����\�Ż0ӹ��M�p�]���Ad���|F����%����FC0W(�~�=��3s�N��Z���3� �Δ�~��sh���i���)��Z=�z!럡sWڄ~��/����x�f������N�����t�C��7�s��+��>7�-��)E3�����]YLA�[�;�g��e4ҵ����+v�@�$-(H��x�F����ǞL��+��jJ���ڥS�OS';=��M�h-&�;���ј��o���e������b���@�`�ʅmi�?�@C�M��{��f|E�~\�-wk3�)�����sj�3=�v�&���&
�'��J�^f*Υ��f�=U��c긃MKg�X�dwx"��?����Bq��z�1w&�:�J	���1��ek��N�\CK&�A+�{��J{�k
��K2�o2��zLVx��ݲ����<�S�'��V�+�:*#�)��?�Q�:S)�����GN��y�6�Kw~YF��[_ќ���i���,�Ӟ�la�8D 9e�Q}pe��9*ut�)WT�+BS�FN����H���'O��5�SH�K�Q���V�����t|���PNfT���ƹ��P�:� u���%�9��W%/��{~Px'����9m��j�YV�p�_��JJ�ǐ`;�%��_ʔ_7:�Ϝ���d�˜G�"@V������ĭ\�&.�sJ��"'�Φ�J�=�a�P|�}}�;���;�/O� QF�Ar1�~�H��3�����ǰ��#��9����~k�Ϊ���.��5 ÎTɱi(ZQZ�1p��x��8I��2�)��g~��g�W���A��<;��HW�܄X�,Lu�VӞ{�T���_�a��:Q���2�\�.Ĵ�;�R��O����7n��U������<##U)!�,y��|}���X[�ڞ�²�6(%?��o�d,�w���1sk��%X4q2:P��e�m()���Y�ы?����y�*u<k?[����EJ�B-�EG�`�M��ɸ�}~�2�;�M��`Qs�%�!G=p� $�YLO�/n���2��u�V��O���2�Dq	��<�w/+9XD���+�VҺ �>�,�#�mk�D/��T�G��sՀh۵C���稯z2�j���ij��>�פ*��п�`|�n�W���#U���jH:կ��w��j
=D�Z���XR�]��x�`�6$�o?bX����?�6�A(�c\#�Q��1��tT!��<B��(�O�- �D�Ǧ��:9�{�A"p��!?N艮ؚX��sn�{ϥ�cI7�|���5*Q<N~wgX�aX�?:fu괨���a��D,��J`�iN��(�f��|��'�F2���{$���бm|*�>��-"���nS��*]"Q'	�[��we��_����^ ��R�x�(,�t�����\=�#v�$��%�
	��%G<�L�?Z#�����$I�(l�j�;�-{�Hc �I�g�-W�122)���?O���.��g�:?�쒮���I.y��j�L~�YhUlN�#X�[;&"����Fh9�%�Ų�����<N��;���'2����˃��x��awL��3\��޸h����l"WrЫ��P���d{L��O�W���� �A�c#�P#4��+�|/E�Y�VE��iDt���6�JJ�2�JT�8��d&CPv�G�$%�7G�Q�Y�Y��.
�.��-�7䳚�#XN$� ����������0��� J٫��X6~L�ӧqG����d�J�8�����:��ڍ#�VdZD�{�89�|T�Aת�����`#iNAo��=#�3�];e�+H��]��z'#+����n�즢,��K���o�=N�gS��yq�G0��.dDڿ��zsKh�j���h!a �ªv����{����MA���obۺW҃'�T��ȥr�ъT����Qk�:��v�C��?Υ�w�2�xݏDG�_A1�yH��bQ�w�:�N���]����$�Gb"��
�Yv�����Rr��GХ&�V+�����n�F����_�Dk�05Z�,����3��5m'o��:�$
�  2Cr�R��S�+����?��Q����;%���!,��?.�i���Ce#��i�8��.)Y	:Q�EUq�`$��_\�ʲ�����$��$pu�2�P�8ʁ�B@�G��f�j�f�����Ghm�%ے��ǯ�^ں9�� _p�j+Hꑄ�k� 3�sz�hr�pR^@V��d�$�l|و��Z9Jw;��4I|��W6{f~�g�+꿺�y��V2eF��He�$��%`լQ�d�;�Kp^���������t7.FQ��y1>͟��hn�/k�_w��y�q��1S�@�E?* ��S.[ҺZ������t��uje��7�54�-"���D)"'e����1�)�x(�2Ϥ���}���&,G����`_��.3���]`Pz΄4]�H�g/�è��U4|��h|���7�H����+
4/�?��[��q�wE`�������kW�f�Q��}?Z���t�ᑺ<���YZ�ϧ���4� Q(K�A�q�z��ʝ`[����]�f��\ou<�t1G2_X��s�E����{�3���*�t}�>"��[�:��5N�0m��
�A�'=`{SO�h�2����/���{�����(!�cg�l��o� ���?�׶�M��w�^��L�g�H���oL��S�4�%�"ўCgk�t�ˡ�`��O�d�MQ���|ZBy��;h�1����m�An�~|��Z�%��f�_�n�C<ׇ�X+oY�-!�)]�mF��x�0�M))x��vMF�:�1$_(�~w�ݦ.{4�.t�ôd|�%��j�^(��@�[U)���������������N*8Zn�C"A��謕Y���]8�x��l|���k*�c�/[�݄�ECiϾ��wTP�':vKqqb�|�۷����eN�+�y�H�z<͜��eW�;��Q존s�DH7}?fc��<�ĺ��A���L�IN�В~��� [6�s#�P����lei{�c4��\��}��D����H.
����	�nkD�2�o�-���ʦQc�݈?��}Ӗ�_�_ڡ&�k�z��˕O�15��8��\ѫy?E��ZX짧L�v#�EC�OҜ�~$�sRUWX1�?wNێ��� �� ���f�9�&i|w2��7S�,q��kȗf�=�5���N>�`�!���f쟠��C/�X#�Ie�U~��ek @�ۼ�[��x�l���nV�pqc��jIZU��E�#Uc��f��+#�����1s��&$�<�oVvg*�එ��ϴ���!�Y����9�qu�� `�ɲ�?�t	��흊t��2r�m��N�;v�쮨!f�k"�k�9�JX��#�Ԙ��1f/�،n���$0�6*��9	z ���P�����f�Ӝ}v˄��+��������w�B�o�樯��ۓ@#5�<�dww�`@i�2p��Ϻ׳��fn����x���}d�Û)3A��&H�b�2v�:Ճp(�	�1��;�<���&�,$K�Y\�U!fQWw�N	W��Ff'��"�,A��rٖm �MFZ
D"�9�O (¸���h����gB��\u�yi�{n�A��c��M�y��;�d	JXZ��%x'5 �z@A9^��R�+�{��V��!���y�k96lǸ���\�E�C9�ǯ/����8������|#:��֥�,�֓F�:��VWH�ͱ��V�߻ynw�/��>��2K�Q�+"m`�ɛ{"��&vDo�~ȵ4��,�t�%x .���=2��h>�n׫��r�NxӔ��ſD;P[�.���X�;���K
�]�=�YBjm،}S��=�~��Tf�����Њ@�������1d��_sC��o�v.�g�:j�ӾW���g�9]�g�� ���������ۺ��'��h^\�?M�@r��#��;����f���_�Z�T��Y��=����8���g��\vN�{)��C)v��J�v����3aM�_!ƺ�(;hR���Q�#���<cE���EҎƍq��9%�z�悶����c�ğ=��m3V@D�܆梔� �z����
���=Jɳ>=�����؍@a��^�t�*�S�ʐt	�K���m�#�9�$ U�#�jSb��ɦ�l���!y�� 2_��Mqk��\$nA�
��n�%1Qe�M���>��H��o�<ꡒ��"����'��z(����e�^Q�|/�;Ş�Q��H?[�{�J}Uug5�7�K*�JE2�6��{~��.���AI���'�YF;�Q9'I���@sG���+k��~�lIL�T��=�����]�I��~�B��PK.�:�1�)�n�Ţ����'��5@����lz�!�������S,klSut�V����B��e������]����K��*�q�Yfs��ۘ|��;�2Z�Z���`�c��$ED��{��,�߱Iǳ�����H�"��K0iS�4�dH@�"]J���/�>��dx�_e���J�f	��#���PFŲ��I_%z�N������ByL���������iW$XX����,Թ�$1?�ŦkL|$U�@��L�۫�j��$oW���,oW4Z�Z���8#��D��
94�*�Wf�c��N�@]J�*a�8�l��IFR[��mf?�O�=%b�o�u�`>\�Z��(�,{`h��NnxV헡LW,FF���y���fIKTM5c$����Q��g�������������=�x�Pl�`p��r}�	�tD	'�[⍴{'_��5��g9w?T����Jev��I���Q�F���H�z��Y�� �+�f6��^��4X��n���ގ2�,�mD���hcf�!��!�z���MX�b)�N_��tk*6Q�|/�q����2c���-�R�I{	�F���<f����b0'�<�W;���K��(�/۽����%�������^�lps~�t�=3�v͛!6�|��r������th����9�T��_1ʅ��P����{�'r�V]]6�P��t�������&�X�B�T�G�&I�����91A{���5����m��BT��,Ų���Fg]0����<o[�"���.%��cx �·�3��e =582<�k?�e�e��m*}c �j�E�Ȓ���%�*��^�]��/��.��	z���
FǕ���2Td5� iZ�L<k��%{�n>D�}.��]�zazUQ��o���y��\w�����Ĺ]�Ǧ��|��V�(����e��P���R0y|����z=�W��.�Q =u�˓����L��J݈/>upX�#hy�UO�f+� /(M���ZL��U��>��a��)�"u��l.õ�(]�
s���lC0�夳�����6��z'���k�E���S�O�����V(��������:���:��9�A%�\o0��]����S\������o���21_*�m���v �m�A2ǉ��L��|Mv�y��X�Fx4e���f$���%0�5�].��c�7Ɛ��tQ�u=*����oB�Gs�~�R���l�M&/����ד�Х�Pحp�}�~�Eثaj٥�qⲣ͋G5���V8$��JJ�;�[Q���L�a+�D�S�o��xB�%Q�خ���/����_�U8����,�#kR�򋇘��$�07��f�hዺ ��	~;(K];G7L��L��30]�R��R;�D���!�緹Z�e�Mr4ψ��Ȣ�E��0��ƨߚ���N���L��Ec��1�G�_�Ai�D�m�{ZJ���:A{P�'%����]��5u*�A���wfVzlOK�i,T"g ����������xlSs쉃��x� �-��0z����4H>���vh��l�]���0��	�|W��FDQ#��s`�����:���M�Į7�b/֒ћ�Bv��tx��Kz����M4!��C��/=��F@~MR����"�~���v���ְz�s�qd��*�^�5ɀӚYۥ��*	�gR��U��T*d�̅)���+����� �0~���Υ�7�����V�?y����I�$�'�}����d�q
DN�)�8:A��h�$�ʗ0����S�اSW��W���,�C!�Lw����c�\�`��Y������hd�n�4���i0K�S]j��%r��&��B�W�����n�-����iy���=>QuA*n�,�S�6
�l��T��7�~�z{�|{�:S��g鰌\
�;������7-�,S
�	fguy���W94��ӏ�9�|�J�lnr�M΢�ND�Ϙ�NSY��%���?'?���E�6i���N/�� ����M�vG �\K�5�u��8؂;'� 5/��� �Ԁ�<.9�1c�f��w����F����\�m�a�/�.������Fx��|55�k��6��ǧԻ:FG>&��j�n8�	SOA���B(DcKݡj���0����Pk�c����saӀ^WI{�RIl�Yn4��r��R��e����ׯ������d��ZR>^��5���9�sns�)Qؐ�˅J�&��X�a�7B���;��|��'%c-"4��$|"�I�����su|d�!����W�������\�ٺ�L�	=K@H,�S�"%��qJ �����s���"C$k����{�����<����H�B��o� �uV�y���|i� �yk�cx�잣%��JK�74�Y�s:�6K���� at�y\��CR��ŗn��R_����1'�˷d��Vե���lU���|��ȅP}D�C/TU�>�	�;Z�{{�@̈fR��`A�F+ә�E4��$�ښ%]����Ȱ��I�U3)�I���O�$;]�c�p1�p
��)w���lQ�QW��� Xހɚ�]�j���s��Dݲ@�8����?��A�]���ѹ�����Ru*XQ�Q���=$H�+1c�U��uM�,���c�g�v�Z0v��5 �IV����c�4ܘ܋潙{�h���(��P��|�����2��\���A��!�ؒV����9��ةƻ�h�?1\t��$]:D����K�h9U�4������i�^7�,_���j#]C]g�� ���Z�m���A+&�?��,+xq�&�F�o��b��@a���J�����6�"��픕0s�3Ofu���a��Ө���gƑ����� �_��X8>7�� �VFU�'�::��:��r#w�v@?�r)F�B�o$���x���C�vzߎ,}nN�5
��p�W"%���݄����>r�ӣ2p�>�{Q���������^7UC��a6d�1�;0�ϡ�A%H�c��aU�'���|9����8�*���;��9 ƻ*����?��n��3�Kmv�I	Byy�b��+޺V�R6�;�B�Z`$I�B��5+$"�aF�.�/z����SM�Gc�%��u��b,j٬�+I:f�:���m�:�I�{]()�v�$BQ	�8/FJ�����w�7ڛl5h�F�I��Za��AQ�WL?�J��1�w%���FN�ti׋����,{�~{�q�0���nq4�S��U�?�oD·;e)N�1����x��;K��t��u�����f�趗b�w/�0�>��g��7�B�̊ g�U��@*�#3��M'_ �t*��l&s�\����P�f�O`d�[�\i�Ӝ"�z��]�.-�������&E�9m�p@�*�����nf߯C�<t�P����B>�h^j50����p�� ��]fP�Ƚm4�Z�.y��e����˒JpH�35-u?�?�'C��&J6�0��$̦�f���%(oP�����o�̮A� ��hN"��p��i��T�r��mD'h�diYS��h�c> m12����,���}��s�v�h�r�� R��T,�C�}ᮭ*[z�,[�0�%AbO�B��!ѯ�!� �������3�TD��|�MH�mǃ�t��|ͱ(�a]�P�F1Ss^l�[�|��]{K���
u�N�0�������2��=����$P�"s�l2Y�9t	"�/�C��Q���\QGKYp'�Y�/�m�V��!�m�Ѩ�Y�5����2�6��e���8Gb����1���~�2��/1���b�|\��922�,:o��ֲj���<�c����  �!�T<|
������ �?s��]����M��lDA��
����bb��i�Q�������}E���6�O%�x3R1��^E�(������bX����S �ǡF��~d�b����@����1&P�M�LDf��O�adR���v��1�9��'�A�����T)�H���ǘc�6U%h��o�ɥ6�j���j?�[��RR7ڼ�f�9�i9�$(_����,'������|�!�_+�/e�!�rY����PK��P��Z������iYz��
N�\��6�&�r}�q��7�d]..Ƈ�4,8�<f��
�1/����5@�Mļ��O�v-�|a�E+,ܞ�@Z�^	M��f������;�6Df�oa�!�}���Ce�;�@{BhAi��Ɲc?Q)i	Ԟ�lO9��,���H�D%{��Ⱥ�9<�45�FrT�#]���>m�o3ڃrݛ����<�Tv1r��F��챓��L:q	79�a��p�ʌƅEť���?D�;�W�+	�a�%�K���w���]�i=�g#MQ'_�Ń4�Zӡo,�|	�e�?��ub���j|��Qq+���h��{>�tC�L�]u�`�l~�DfvZ��y��!��d����4D�Mǵ���o<�l�X4�|���a�?�	���PZX��K���^и�BW��.��t�����#P�q�RA霥�ƽ	���p�*���D�F���C�_�_��i��_&�B�
{,��(!�<���c�o��y�����r��Y�>���u^UJ��YW5ސC�a�����Ց0�k+�?Ί���^���sЕ�������.ɾ�ZL���<�?$ӯ�����,�:����]T�l��17��S�K�.���y'� �e�z��G����c%U� ��T�5��,��N,�JvK(B;�2B-��O~��ˀ"yUX�,z�Ko�ӫ�!]eޏg��vO�"�`�C�H3V�V�#&�b�i?�쁳�]ٜ|�+Φ`��=C@/"7�S��Ôhbi:,�n�*���ruu�t�8&��9���9*���_E y���@�[�h��@���������f�#����H���/?�����r�H4V������~\�#,���
[à�%"Xs�C��N�]�/����b��<�5���Qb������̔����ؕ�dkօ�p��M~�u)�QN~	�C�ݥ���}8`�
0�H�Fgb7�����z��L��h���q�2�6~(�g�t�l��9��ȴ�5�vE`9�-�
�Z��^�2 �{P�|2c�&�J�O�Չ?l��v��u��Ů%C 2 �,ĒX������L[��ģ�gi���#�X�D����b���)@
~`:���-UL%p)�!��'�N�{MbV��!�i37���8V]�����ٮ�uR"p��MI'�e0N��^$��_$�������S��i��Xu^���&��ײY4�PQ��a6�"���f�a��˫�O�k����K̓��qv��S~E�fL{r��ހi��(�ɟ����2��Z �-��V�]�8şJ���g(v�1��\:?��ϲ��gx9��%��U�}@�	���2ܢ	'M��>�+E��:��>�*1o��� ��Wx�6��{��v���2&�����j�B��鈫_�D��>1�x��Jtר��%�
?�ΓpW=��{�&��dm�@t�����q� �TO����V���J�\&�r�Q�<�λ%�_��m {6�@�v������I��Y����8��@�`Pw�#�;T��־��R �a�%���z3�ĕүRRrr���I�kEB��ϯ���ɦLな+�7dMJߐB�c��	�y�l$���3�5Im�U2Q��(g���)��ת�B�D���́4�$z��<󧏙W,(n󂏙�t�O�l��Nl"x�eü�9p�J��(/lS��K
��-E�x�����(�?(�ϢT@nY�/l�4��N^�7JG����d�POc������#�UĂ�Dx'q%ˋo_>�f�Pk�rDHy��(��Nl�u�ϴ���ew�=���v&��}������H����������E	G��k�rޚ�!|�����p������Y��cA�T���?ӫ���)P����$�8�g�L?�Ц/|&loj�	d�B<���0E!�Σ@�dI.����U�R�L�u"��x�� W8 B�<��DQء�cb��F�C9�f
�3�����9�Sʊ5�l,2���Gi�#�;K��s�tr�:�m5��+fݖ��� �L:�WW�p3|��=�}I�L}�x�En��<�y�̍�%�-y؜I�k�*������Q��⑟��]{6}�f%�7�	;�H��b�&��H����������(�g�]�͒��ߎ�P�XVSȦ��֊9����pа6�dzĕ�d��+�Il�����'8քh�Ĺ�&�5,#�����ѣ������yrEQ��-z��a��	�aV"|/���q�n=P	UH�~^�Ί�X�����Q�~��Q#��`XR��$>,'�o$cV:�[/�K��#�9�Ov�Zt�ve��]K� N�qÜ�\�<�5Ujh�G��)Q�(�ۧu�J���$ ��*�8j���X�w��+V���f��U�O�j�'+��Pq��)]�M��\V�'��"*�ua2�~)ܷ���^2Y��71�L0���-�^�&('�R�vN�H��� �G�����^�WN��S�3v�bםed���:?���Z$g6#]��s!�4"��y���j�TUk��>2'7�f����D�a��fYUH�,�F(�MO[(Nê%�\M�v�IN-����9� ���u
��P׭�V�?D|X�k�R�?���"�⋩>����񱈫z��F��j�F��( ��NuHI�Y�\���5�����/?��I�0�}������%�J�}i�.�l}.4	wIN"b<�ImL����{Hg�p#��o��=��;�����'����-٪\{��(^��]�/�-�鬱G�����{�?���SP��m���y��u�_��h|��;�κ�R��-�^���Ԭ�%]�>�� զ�[!Q!�������ңd��T�����G�8�B�����s�XF� �J�B0k�Wg��b��+�p��UryÿC*Y���ByP�*��uv�KtWy0F�w�q��O�ݫD��J=`�w�����y˽t�Ke����Ϋm4muZ��%M��Ղ���*���ci�k[A����Ym��>is8W�[���J��]9�K'K�j��[SMN\г���*��̟��/�,��jt�M�8�
��^��#4翯��>3mEUMyez.K�`�DƐӡ�O�/%xk'�7#����@��`��u�����#��K�낤9�	}~�E��?����U���H7�g�P8��X�A��R*s�q�i��8|�a_�/���<"
hn�J?\�L�4)��7Y��zU�]��cz\�5�����(Q�F����'iD��Q�Nf09���c���d���w��_�!��+<S40����v;����׉p�li!��a$�i@cH-�T}�#��@��>+>�W��iD�Vä�l�����?Ȉ��gj�ֲ�OȲL�R+[f�Km�e�G�=ܣ��wRi���i�ҢTӍP��XJ0�t%\w�IÁ��d��O+/m8�z�Ր�t�T�{' �,
yb{����I�igb���	R��|�<X.����i;ms�Q�D�,���7	.�tҩ�C�Q�ZD��ᐪ��	]Ehk���kd��4��~���Ԛ:	,�O�Җ����0w�X����ݗv���\Ӻ�1��#`o\5k&.��Ҁ��Gl��J0@AV����J��-��`y���`�);�9 ���^�<gԾV&�H"�
T�(t�+[d94�{�jf�Y�5׎�g�j�L�T+��p��J���S>��)��4	9i���+nbs��&8�$"��t���PJ�k���Ѵ�N=����O��W�]V�����eʶ���Va���Q��G��aaD�3_���cԢUMm�iVHl=ֺ�},���f��k�-�zDz�ɟjX��V�U1�&ӄؼ��_4��e��W!���H+�p�ܕڜ-q��=Q�T�� �I�? �q%�r<�"��^��l1l�gC�|k2	��Y�H�2N *��/�4J
�!��w�S�%���G��k�%^�Qt�z�����Hs 	��(0,a�݉Ur�|Ƶ���O�]ۛ�')|q����6�8���2�� ߦʠ�x���!��'t9��6��������/�*��)�!	�-N�Z�7;��5p?��]�x����$�Ŋ��Փ�b b��Ot�)��6K6T�a�|���ʘ�#+��ܯ�o��-5�,���[��zZ#���]_BNw<����*���g���F�֕�ܒ���v�ŉ���nϡW:jW{�N,d�u$�µ�t#�kBg��n�A��ݒ���
a6�{Tjg��N�����j��B\c�Kl�w�����5Y2
�H�k&������d�ż�mֈ��ƣ/��#�u[���y\��P�Ai\+Bi���oC~�_�@�,V�w�I䌉�~N�NK�u)����m@aԣsB%�=�����L���Q���q����l��<���I4�$����,������o��vՏ��/���嫳C��\�~��&/Fx����6tH���:�b81]w�����O���ap[�ER*�8'�R���G��h���4:�6FwZ�2�4�x�|�Nlk�'�7��O���U����M��d)kp���8'��Ge����}�ޱ�c�Sq=p�q�����q$�v1���(�gΥe���~B����_���mց��8�I�7��B�yNf��O�ka�>C�r6h�T+�{3��4�v�+Jj�Ԝ{aI��z
���p�5��"�;;��s��͖lǊ%4Ų>��PI0��r �EU�`�uWN+hj���%��A�P8�>�㣌��U��!����p�����Č�Uz����_���wײٝ{�j�\z"�����������;BK�P�bñ����P�� 4  ��:�Q���^Ĭ�6���a[:qz5(>�"j�l�$�:��\�D�o�ǝ�&����z�yu)�6��L�?� Ql�V�Mw1�<�]�<RIʖ�{�����sѯCȢ8.��_�e
�x�`���fnCW:����>FTQ���^Y�{6|]�:E�����d1	�� �6*�|G	疆�������dm��mpyag��8����m�(MU�IbF]���
L��J ��P��>��Ά����5��G#�7��޺��H�fq��qL]�MP,}u|���1xW��4_���V�]�5���'Vt���Wy+fp�y���b"(�é3N�*S���8H�з��=S�5桭�����K6(nB�|��?"��`��Ac �汅�����(1[�y��9lM� ���H��ڕ
|�WW)�d��1?�ژ��I� f2���
R�=� 7�٭u��a�a��A&(�Ē����f:%k�0$F�Ja��e��y�v)�#Ȭh�Imf��D�bW�{E��lWVr�t�}
Ik$��'x�� >��^�f�{?oōb������lx�'��?{N!�:D�#Jf�W��ƒ�%����?�
?"IХ�����-����_k/A<�#�y9vZ��d���0,��¼շ����`U� �a�^�c�"�&r��	���v6<���}���`��|����
�/,�<��Mҫ>U�1M�r��ЃQ������cୟ ~�P[�Q�4�����U�eL�~iҐ��O����$�4Vҩe�$cyM'6���XO����V��L`O��H����[*��I^������jE
4��Cu&z=�Fٮ�U	���������NУ1�C�U��Ѵ\Zf%��J#w����M���N2<L�u��S6�!=-��P�tkVy�<ANe���na���Bl�[`���@��i��L�I������=N�>�^QJНh��-���(oM�o��i�;>	�Z����l&<��EK̲�CI ��Ŀ7яn�
�U��6��3�����]�S���[XZ
���k�la���'��#������5��ep��( ��Tgb���'K)��nbenN�8S��y�Zx)��~���y���x�`jy)݊�<d�U �p��Oy�q(�q�p,�C��G�_��h�-���8�OHHB�jO�9 <\<pv<h�S��HJ�ϲ�`��a`p.��LX#��y��-р�u#4�}�6��1t�z��ƯrzQ��Zp)o��K�է���9��kR��W��e�=Lܬ�4��ϑ���CA`OY���ATg�(�]�./
��y�
s�Y�j��Zރġp�%����	��¢�ҳńU#���;����K���c%����y���o�u2&S �?hCx=oL3�^�Q������L-p{J�@{@A���(��&�/�}�'�Y�k�����Ul��F����;�����iz�Y�FC�����џ^"��}1�%.YǭA묀�"�X�����_��w��dĔ�,�ű�g�����,^f�v��Z���!���Ka�:�?�Q�J��h����Y&��-�vh�m��c�'�D	��H}���g.yiD~7��5�f�nq�����*�� h���.��D�4UB��v���RT�D�M�c��߭�� �=*�ƶ/o�V�!��cW�uc�����*c���e:�bI�B칃;z��2~���!��:�>�5�_ ~1u���e~K���Q��C$ c��fN����o:F���;�j�|[~�z�� ^�̀�ܩ�(4�rͽ3�#����Sҿ�'�ڣ���FdMK�b��㷿 ��1K��W��5 dB�c$��%ќF\~{jଓ�+�V*QO��WH7;�a�[9�}%��V^δ ;��Y���b^4֮�e���B.G�Q��d����m�s�Hn�[�j�녡''$�O�
m�Q6�f݆ ��xk�7XP�`D���r��|�~��z���Wuۗ)�|�,����B?:�l��t�� �:eP�q�[6�7�dY�F}����ygx�ۚ�偡ζӆ�\�cl�d�uq�Η�,��|��i���-��ʭ�<5��!��I�>;}Z��{��X��b!���TȭCa��-�I���R�,i��Su֡urB�V��h�4�%���tL������(r��r�[l�塞�� �bl��]-�Ϋ�V�O��Aj<���o��4�,�����XTf�3j��70\�F4�|A'��<���v����Ɖѓk�<�d�j�m��i��u�#�=�X*�s"	�%��2�����^I,^,�*1 jT��t},,ߍ#�꟣�,��Rp�&�Q�*�K�&&]�}s1V�cT��SFR��U�C�!BΆ�v�����nb��y*�6]]5���B</ׂ�0
���r�܎R7�z�h��_@��{�+Ģ� �]~ �6$|�?�D��cY������
&�7��@� �bK��O4�I.��Җ����ƒh+��[̑%tU�Y8���M:!�K��c�x��r��0a����|w\j��������vK;57���ۂ�]���4)`d�eN���o�:�n�o� ^,2+��=8) (:̛��t����'L����y>�eqH��>�a�N2c���A[�����q�k��A�����/�a���Ȉ�P���h�zfv�3��;mY�N�>:��4�1��P�y�B�������s�(��gk2٠���7����≗��\��K��t��rԧ��A����U.��t��m�i,���6y��0������/Y�J!�����ɹ��\�]�����q�Ik��@�O_��3P���sЄ�L�@�o4�R+97q7���p��f3�΀ �HV3�|ߔ�xM���f~K���J�ͤf(�.���;T�`4S4�����[�	�tz��w�榐/F[SUԯ)_�h�ZYjbp�,��Us5듊���۽���F�'�����-q�H6f�H*�y�t��ne��
T�S)�H�O��S��?�w�)i�0�1IBd#�b�c��+9�*/mF#F��[��Pl��9@�cX�����e���;`F��������s�$ϐ��f�|��)�h,p%��ө�0�V��J
vK��v���Ă�cq��+ry�f����/D΍�tV\%d@\g��6�5���!�����U �Κƶ� �WW�*�����D��X�b��Xn�B��Dr�D1MssF=�,��5m`=����X�0n"B�\�9;�F�K�Md����d��TfQ$O_9Vǻpqp<xkU�t��*ٟ��ى�"g��&��tўJڥ|�bS{� "���A����n)?4���ݫ���u(��tT7�2C�K�2��m���\�Y��G��/���Y���ڛS�wkO�D�=N��+ �J�~�\e	 b@�(���b�/�`#�(����#i��R�h�^u�d�y�Ӄ�I�+Rp�|`�L�7Q�~x
���]*��r��Y���2�i5�*�/ϱ�qz��[ʐL��~���XU����t#� 튦�q�t�7�:��h����ʸ���v��!ԋ��9k���� w$�c���#L�����[F������^�Ϸ˕�x�x2G[�:N]�C�̯���"ʷ�(Q��|S�po�C�a���َ;sb��}p�t��d���M�D�]�4c�lx�z����6���n�Hq"�SЙ���^������$�3�n��ZJ9�v�.�-43n��.	B�� M�*E&ˎ-�e��;A{�l�k���I׏~�,E����2m4��Wb��N�|��x���V6�0�8�:`-�����q��+�U;��~�m��@H�v #���ރhoM�}��5����?�Y���AvK�f-I�-��Ĭx�vP�E���#�Z>�8B=�pp��8Ʉ}�B����-ߞ�dk^�EO��y�>@���/���n�秂�*j)(D��I)��N/�E���jB�j��Ώ*]��0{	�2<�?��[tv)s������d8�+O���6�R8�#.k����p
#`�򩬤��k4ت�I'��{�_ɯ7�b~ �����J+�}Hu�W��W�_�J{& �+��^�0���Pt �
�4�Ό
3�Ο�{6�-� ~�f�7�Tg��꿢��g���$����%X�i�wue�W����72���ndHd��~�ik���i��]o>®L���:�2�cG��F�?âN�6�3�o�t�$�M�cV|�'q2�y���w���"�g��DX�ų��OGq������i�*%�V��΃��g�c=�r#D')H��(����&�Wm�_ni��fgw��vv�� ����ء�����$�='��x
�,^g�~��ԕ�GW���I����n��ӔDK�HA�
w#��x[�"P	rBn����lJ�].�)�So��WmqR�I��tK���p��>����n
h������ь�˻�g-7`a�WT��5���Q�;>.u5i�����@-�6�V���n�` ���=�n�����QM%J��8��ޙ���� <�%�ў��\����okTH�<-Y�@�̈́����z���Q�@�����V���Q�<Rz7{����4j���M�������-�,�P��w�l�'��zd|��f(T*����2��Ci�vm������)]����ǃ����v�UG$���.����%����Uc�����_�D�K������_l7Nfy��ZSP�@:R0�r�	����T�SԓYi|�r��!��p�`(G7����L�n��;$&!�ɤ>+ ���*�`�6�����3H)7��n�!��������NƮ�� :z@D<`���I	G�Jl�c� ��[u�W�k�R@����X�)��*�&鬡�mMA����<�_.y��@f��W~�G4�5�xqM��ep��grR�t	���,2��!?80���^�p��*!�{�?n�R�_#�z�x��W�Zm����\Z�X2k��N�瓌ٖa��a����\?֘��?n�ֵ��@��������Os��(Ȱ�v ��D�Ӊ�y�B^{Q�.��ʉU����z'mO�v������Ժ�o�W_e�N9;����FW�:/w�p�wsΫ�E����N!�З{�zhh���\w��N�~�x�'�E��P{���8�T��'R��ʑ[�����N�L�q�\c����DDĊ�YN%�%!@9ç�b��7�w�5Mr
 ���n)�g6�;��Q��&�
R���1��4$�?�g���*w�I��nCB?� 309��������(:�Yةc���	��#H&3�p����䒿�d{x�YI]��{���E��,u����?�795V�"Ӱ�D&�+��<��qE���B�m-Z�)�=���p��s���2�sP"W2����N��+���
���M��F���0/���LDO�n�G���3j��O���84�;'F��Zď۴��. �i7;Lb��oo���/�"M�@Y�EQ�>;a�`��䇉�>=f�L4T�S�~�>.��w���J��'iH�7o	�Z�2�V�~{yN���\Z�G��?�3Z��Q�mH��8��*��ܐ6sI�ބ� bH�Bf�KP���@_W2�ch�7��!���h ^���7�B��5d��!��f���y�h�S ��Oٝ�3���`�2T���>S6(�̳'֑��<��9#0	c�����ù��:��7<lC����ȑL@���`<�X�;}
��-�ԗ�N�j�V��aF�>�^ւ-��ã�'Oh7?٢��+?.��'Ir�:'�bw�c�ؿ%QL��u�Z9
�������m����J���{��^��淡�"u����%�|s�d�M��4F���;(J'L��B�QjO�jF}�ˍD|� ���B�t&[��,ټ6���~�4�ɗ�5Ar2O~����(��݂@e� ���b��I�W@�4�
�N��v��z%r�f�����ۈa^#C�s!;����V<�C��aEE��pA����*��V��p7B��$�W��K��9]׺�,��u����g����N>c�x��̴9\����t^*a q۶������?P^��}]St�i���85q��	y=���f�9,k��:�~ڦ� zgZ���S��]����%�\��ݴY��b�Rj��;��x�C��jCc�(�,E��	K w��q�&��(�/�'b�����Q��;a�BA��g�Є�dVL��Tx�I�� W�V��O�����.���Vt��.~=,Ɔ	r�h9������X��X���"LU��٥�<ɒ������_�7�2/�=�ڑ~�:�q�C��7��Y�0�A0��$���KU8��7��{FM�_k�f�l���5�m���hK�S��^>�@ĥ����XY9�b�'��I�)0|ͺ(����}=��$h8܉��8^7ׁ��½�u� "��D����ҡ�];qYd�;D3E1{�[fc9=7 �)ѺК\w?&,h~�?�L����W���
�x�|9Yn��+0���Z��+T)�<�O�2h��-���Q���[0]R��~�kA�7?;���
K�\�6�у��ˀ|1�P����K��t�,F�đ��Q����bC<�n4]��ԙ��f���8:R�����=�������Q��̬�88����0ym��NB�n\�����0p,����л��sbf�0�8�cQ�ͽ�h���g{~A7A<�"���Ke �Ɠ����S��� ��J�4�K^�-x�	<���⹨�w�b:�
&VE}���j "3"m]w��"�7NE�r3+�%Mu�5g���qBAO���CD6���)����
���q��5ы2�]^����a�!.�x.w���~h�1��D?؞K�JA�w�h{�z����zf:?n�)�f&U�G���xly����6���-��kN�+�!K\ 瓒k���@X lV���a��8knw=c^B���pп#��2n$I���Sw��Ƭ@"�6���Y����
l�UK�&
�Z~��:�h�P˒j�'��l^K��I�0����|(�Z{�����0�3�Znƥ0�[c��Yu��-��R_/n��^�	U��XYD
�Mh�Y-b�d���O��5�8�,u..e��g0�n����*��H�jT|�T�ߎ*BH�n'�:�A�nU"��@Iqm�Maf`��#��(�>#�խ�� �ȷ%qՖ�0��H�,I*(rw���bm�/3F���-G�6g~Va~jye�Ck+�>�����F���g;�Ks��=��VO��q��)�h����0G��P�j�������'�8��A��wPqPp~�W��$���OQ�NĊ)��Sd���5  �L��h�Y�ɡN3�JX= ��(�9� dnhY�DI@����'h'��B@'S�w��J��Աȼ^��{��4�+-��?u��D�_JYDI㛕kͫ�b���f��q$���֊)(��~���@T�b�l�x
EBB g|;���3*$�<�jӤa���;�r���g����c�bۅtE���gB�MZ��Sb�Z����%S�r�|*�
>��E;p�J<A*�M�^%��߁��W�9���n�y�,������
C�+c؏m�dЦ"��w	Z,u'��=��`�T:���6��(p��Ŗ�����8�T�k7lY^�:��W�ϕ��Z�� ��U��.o����pP��Z�N�ַ�.�����nnp�ܼ�#W��)t���=5	�N/���5}A(S�v�pv�0��ˑ��
�.���0�ūc���K�	-N�r��ת6��Cq+0�j�U(�Ob������'R�Q|Q�H���{/d%�A�;���O�T����r�+�z��y�Jl��rM��M�^���I�!)��X1���:�	��@=ݻ�ZE;��sl�e��h�0�8DT�/��a�ţd5�9T�)�`b�z�+?��}&;���7.o���Uz~�/�T8I�:O�'0��wz6�0t&������Y,B�)��8?�7��; �Y] 5���k
�ɀ�`��pJ��!���=
�ݏ�<��s�Z�Y�*��&)���20����BO������͟j�;J�����5-8HIy��YۼY�Mk��y(�.y!g�����J�6�?��&��S\���t��57h,�#^��n�;գ��x0!TtJ�0C�8uN�pvȦ�#����(��茯DA�l3�_i���z
�	��� 8���\u~�`�i��Wo�gb�I9<��<����y:�Q\�~ƀ~��m,ݙ�����`�-P�S���&`�g˶H���)M���ʗh��=A�� [�'M�%�B����?��D-9x�y���YH�q6ɭrf�3����5p8�A��=�C�%��uE�hS~��!�}0��w�1ψ��2�����_�	�RV�~������-�C�PY|���p�딄9�*K�rL�G��=����O��|������DZ*���0�Cr��wR`�����q�v
3g�K^{������!�3��P%
Z���8h�������D�"@���>
��
�K�f�:��bҙ���Fs�#S�{�Vs||1�py���,)~3v�膷5{���f6�X��7*��P�}���)V���X�d,��B�h ��Zs8�'f���*��o������/y�����.�٧�(kd�V��P^q�ӀG�vF�
	��C� �bn�"��@�:�𴊰���P>�Vۯ�f8,��1�o�*������}���#^ᾡ̮���X|��U4�g"�� X1\`��{u�l���'��d&4G7�I��|S���d;�ty�RJ�P���S�A�~ʢ�To`636͊�^�C����Z,@��5Z ���u���(�	�R���<�U'��a ��QBŜ�r"o�s�`PL�mD�XU�V���^I�@��K��J��Tش|�16�	��գI����X�u1	�;?QY��7,��	&�,��aΊ����$StD.Ǵ��6tFj�t@�l�*M`�����#�`H��Zt�RjYL�X��D�E]��L���]>C4�q�r}<SyQ��/_H�����yA��t\�x��H.U�'F��ی)�u<�S����\@IxTc!\�Rqu�h�����F�m/��!O����AX����R�˭a�C�����#w�w�b9X �e�+��\~Z�L�RL1-�;�z/M����KP�e�{��gq$���Y������;���-�{j���Cc6�&	g#���O*����&k��_J�8V8n��\�b��Ear���b�$A~Ue~6�)gy����Dơ	l{'-�g �����a����B>(���sD�9�iW0�YX��������x��|�k�h�G���`~ΧjO3�0�z�l%��O%$>��wc�1,o����
J16�o#�U1�8A����^��X�����C��4����w��y�A:���pK�����"���c�B��z�ėXX�Cl�lW�\d7����>~�RQ�2z(D��M�?eH8ru�C�o�y�џ��E���G���ݬ�y#�F�;C�����Lu�Dk�Rs�T�WA2ʄ����h�F��?v4�c$s@:/1L��О!@�cW���Y�m��S�S����3v)b����L}Z����[�[����Q�]c����U|����Ly�f����x*�� �y����(f���@.�N�<����\�mm�XK�;ʘ!����z`;�H�-�TZV�ʜ��W�Oy���G��	��Kl��T�?j����]�;WT����G(��8�#,��iR���$�]jy~2kBI,�PHi��9��"�A"6�8����Xk�T~.�'v4���1�,I�m�s[C���&P혬"<�(2C�w�i�Q��H��7ο��BOw:�P���������E��zI�XR�6#�̾%u^iO1��ɮq�5���N#�4kHR�`}}~��^)l�N������lx{�u{��Z/�j�q	>�����z��H��!�M;Y�6_s@Zfoɶ�#����OЖ��WS(�:Ayߘy�K	��O9��n��D��a~è�/W��[@�7gD i;���%��et�T�
���b:��| ����&'S,��:��A,�9�AqZ$8^�Xs���Q %�7L�K?_���������=��� ����¼sedSA'�ԲTZ^��b���C�]�Y����/��?k��b��[P�ک^�N�2��h��v�m��ne��t��4���VVx'��օ��1���:���4�Ї���¸R|o{@zk�}�_�F#��8w��/�U��w�~,I��k�r�7�*��Tc����8�n� e	mK(�#Ca>�Xۅ�r%����k�?W���>'���^2�({G�I�HQ�	�~gִ����;����}:�w�ua�v2wq���w6�\X�?
6����Dsa��l~OS�J|I�<�D �h�.�%F��YW/��L��O�ct˯	e��G�UeD��GU���c.}���� �c�����]������D�
X!�?�P z�.�U���۔�j�B�1�j`����I <�S��
���k��e��N5�x2R���	�=����$rY
�����E��&��@��8Gz'�&���_�H���z��NM^�����قqS�Dݕ�r�7�A�$N��ڼ�細�v�hhQG������6�-�o�*%�}#��_���*d�����*�=T,޵t<pqVƑ�ҧ��SQ��͑6�(S3�1Ї�f�G�{��`��>C�ڨ������p���~�S��7�]��t:˧^�_Ik�ӈ̑�%����~'��2H)�T �·
ɘ#٭+��e�$� ��da��^�L�����b^� 	gd���_S)����$���w�[�@Xb�~L���~m\jy	���_��1pM��C�U�E��i��2�®��1s�����<����E ���z���?����U�)�K=�t��r�
�i;����~�.oGKئ��D�͘`0�W���D�[f`�DѴE��V@�"�h<ќ)2b�[���`�$�Q�K���^�ۄ�7�(P��6�(�Y\�CT}<M�Q碸�̨6L���n�}#r����#�ML��d`(�p�BT�Z���L�����[·�<6�]D��WV���z�j4�:V�l�J�s-疂M�
y�ҸWWJ��G�>�2��88�x�������Pܙ�Z�CDd ��3.�%LCF��CP��'����ZK�u}����Uֽ����
����fU�ȍ���?Kͺ	��!�S��}��U�:W1��_fQ��)�[����-���ވ�/��q�D��!��Tx����`%r�3�NK�����.u)dH������$�>EǺ4������P��a~��//eoQ_)@���\�d���|���%q����0[��nڦIU�I�\�@�L~�͟��t,�J���$D���@��st��HCc'�<Y�����J�'�U� yv��:��X�����9��Rn�ضY::���<���j·��l�{s�U9Y�I$�������hR�z"��Z��[Pޗ�F�1����p��ƞR֥�>�A��t���������w���̍�.��J!�tŕ����C@DI�'P���e6UN���!��me�ެ�� >�m/�T�VU�0A_|�)��q�����~��A&m�0Eś�T8I���;��5��=���T��n�}���t�,h@��u���^�Sߕ?�
�;v�O�[$���fT��l�Yg_V��d]6��^��w{L��n# �
P%�+�e�M̟��?/]��+�Y��JnfHfB��h��a�,L�C���hа��W|Y�lsD:Gv��I��椿ϳAG��T�}4�n<��vo����5���WیF�<UX�_������1���	�}���O���5�f�7��@4^H�٪���~_Vl���sr���~pRAg��TG��>�)�,nl,m���])y��	|�������`���`���ꅖ�����؜�|�>��  ��I���wG�'�)��+��ٺ�-�;�A]���=f�4~B�%�#�P�6�YO�R��y"�J�o�<����֯H�K� U�>=˴���������$�.}�&���W*�@VU�]�X�}�a�8l��'(�.�E�3!�����_���n��eXʖm"��.����E��j��sz�����s�Aǎ���{�ɕa
dS8A>���� �^q�l�Pq��������a�,�ysI��%��A�t^���~i6
��~ �����\z�5w&�y����kդ�����2z�1�B��߹0�������N|���S������n4�C�O����(l$�m#X�p�ndI�\�!i)�o��V��%Rl����=�[�MM[�Z��� �;����Bg�ۥ�5����c9���ӣQ�q�_k&��D��=���J+^	��b_��R���c���m�A�x�+�m��>�gJ ����Nݵ�/�Z��ϥv	�PQU�rb�Fg��â��c����u��j
��h�>�2s
�'�x����b�3u�īҢ�ѱ?�c�(�t,�G̢��w/kÎ]���)G���a�G@H%���/�RD��1d�Y�7����JGEV����ˀ��[�$K��wxQ�I��tzN��&�,$��̢o�����W��K6��G�6�Ou"Mܛ�^� �)��	�3���c/"�=�D!�"�-��O���W��?���c��*H��	Ew�]��]{;��t_�5�"��ԗ��!�X��(��ׇ�)-�4� P#n+/FtV���cձuc��20�10~S
 ��jgP�'<A}&��ņ1�l��h�w�̍ii�� q�B{�%d?ܡ��iC��;�%M�}���������6��5���l��z�7W2���c��lD�e�}��(B�!����TzF~x�=~�5#�5ڵȮ;�P ]Ř�8�@5�כ�p R��7W���>ّ�-�?fRY;��}�Ь�*kg��t���XT�� �[�fi�[�h��wy��'9�/��ۛw�h���J!��ô�K6'z%���@9��B��9���,�>�_���0�e?�=$)��Q�栜���m�����7�t�
���y�1� ��<&u����U��S.����S[�b���]�y�	��E��ﲛ{�<���TJ�9vn��� �'D3��3��� (yF?d?���+R\�ѹ��v���u���%��Th�Sr�H���ܼ�"T�=��oq͏&-@<D�T�&�@Ї���|���j�����%.�R:��OT7��F}������S�̚���6H�G�&x����љ9ɣ��;%�x����"����+�Y����jB���Q�Qx���ݵ�U�rG��b�S?���<���	Q)�KeY�UU�ֵ���H���a�&�5��ҫə�e������Jkh�'�����%����'�� f�ܶ���P�P@ڲ�t�AB��E�����ܧ"���ॾ���J���f�ϰe!�h�	�����rN_��w[�����ڂ�1��k'��hp�ɋ{v�~���m%�Wa��O�����AU�)m5"A��R�K<o�}��+U-�i
N7ʯJ]�@�@��(��k�f^6���2�,]	i`���!D�ʓ~� �y�w�!�YO�-�HVhN7��6��[���-�a��䖣�`�.���֐Iv5�{ �6l;jM�p�aԏq0�K7�y�|�Vv�'�f�5w�� �v��[y���<�[�qt����[`_����A.xېt���I�Z���M�a�)��݀��ݚ�����
I>�Q��}�� ۿ�9r��|�'�H4P�b�lG��5Spu@۵ �2n�7�t��x)0>!5Ĉ��D���C�#.|�2�����۞�9���|�HZ�|�5��%^���8⦄E�2�!A.�tu��M�(G 3Y��_��NI�m�,�<Ϗ��1��;���_3;ˡ?t�$(�ix�A��
A���D�XA��e��񘥊X4�����p��~i"��6�]SO�� 	m)	J�}�f@ݑj��&ge^�X-n���8
bPm�;�\���Z* S�
P�������Ơ��e�9S��-.FL7Qݓ�a\zEx	Sa6fc��R���e�T�T�:\$o�^=Jƫ�r}/Y�`0�d��v2�Hb��\���>�h�3���sz��(�J*��U���P%��C�2�C!�&�f�.?z��
�y[�ժ�Q%	�?�����,�Ȱ���9�+ �<!���'��&�Ĉx���(�3��/ң"r�1Z_y ;O���t�^^�X髋7؎�K���Nf�T��Ya�t��:LP
���s<U�,u���L�@!
O�����O���`3�â�U�
��R�[�'���䶙�������8��u����0�A1lc��9SĢ�+1D������i���*
@�r��er��i)�>%�W�Y�d!��<�ށ��%��ZW�a���M\g5t=��L���F'=K��"��^�Qd�V�Y���t�B���P�s�VVC�٫�TG*�;�����^\&�e�����z[���y��]��Z�J�X-;G�}��,�l��Yݠ3q؏��/By#~:�(3��k�P_���7=�U�Η>h�d�ָ�r�xඎ2��c>?']�=HQ��L�a[N�teN��o=}&�N�qhc�y�݊b�!Q������g+���[�<(r4�	k�3��Ɍ$(�5�mF2��:�>�@��AU×�R1�VP1�K��r�h���i�������]��u��E� ���g�c�b��z�D1o^�W��6�[���|��x�[T=5���ءTк  ���a5�Q"����#|�+�K��Z7��E�����9Q/��j�کR�p�i-��QS��N�Э�4F�����ϡ�|��F`�+�3�w�[�7i�p ��ܕ7�eT��d���Y4Ԏ�{��%����z�4N�F� �'�.wp#\�jkR�3��$h`QU9���U��,��i,*򧵯r�׃ʼ�
W��A֔*=na��x4�ퟶ֔��]fI��j%�� !�@8J3tV�|�_r�B��$�>Gd�N��Ծ��:�Q�6ȡ����`N3�G�;+t8q~(ѡW�U�M��))�|f��b��t>p�R�|LR�1����jn6|�<���e�m�Z#��u�en�@ҕ����4������	鮱$/�	�����W�_2R��e��:��Kj
�i��ֈ���`�n��p��̹�H>v; ����2��y���Ԗ8D)s�7�ew��?��;���'F�i%�� ���tr"ʆv� �@悥�p�E��ɔ��I!��>�Swni�.���yHh/+{�*�� �=j�ގ��7w���h��F���}��5�6!�g�(�MYT��w\%�l�hAy'��9Qi�N�5�v�X.Qj63g�֋��%�x�]"��Ķ�$�u�O��a����:*M|���� @�r!u��Za�T:�ؖ�ٟ��1w�B���C�X[�(�>��W�+�G�L�z`��0E�z�ĺ���!U`��9eR'�xtܶk"���F�P&���.�� G)]:�,�ÿ�+]�C�e���n�w)�r�RǏ������*��ή�y0nC��<.�Y/�t����@ˬҠ::��0r�7�$��Wi����� k�t��-P�?.��T��c]��ow�RÉ���9晟���N�!ҍ�8�dݸQ��9�Kث�)4
K��3}��xjЏ��򟹈7����mYT��
Y��,.�#������6̹�F�k��zw넬��?�$:v��Ђ����u�Q�W�j���E+E��g>B�LC���q��n�*�0
�E
W@�o6g�}Wo)_
���d	�t{��� m�h��^�H"�\�6fO��@�>��J�M��0�_D7���{@ ����O�W��M��zƢh�{VQv�|�G5����Q��j��	��w�i�P�y�o��/ "��W'ZQ���Ēq�Q��~�b2$�l�=��v:��6�q|]��{/͙��_ϿM�ƹk�:d3�:!ب�%����T@�;�U�J�� Xi���Ǆ�����U���M�3*�r�v��;�?>�l��j�]c|u��vf�gF$��Cwv�A��w�� �5���xئ�d?�Um^>͌'�b5�?��@��\��w�T�CWc�b���`Jk�8vi��=���D��ｃ�t.�J°:ʌ�F~�鼝�<[��C��L/z��
��T��wXP��y��i`��d����ss�vɵ�6��+�j�J��>����Zj�<O��\;����M0?G���5I28������u����V\MΒ!E���h�.�"#EJ�V�Yvw�v�s)���)n�d� �C����ni�U}�\� r'��D��2g�L�T$�v���z���d(�����CD��fX�t����N��`��_Îב��ƀa����9�!���pT�!oI�����z���̷ϴ���$5>�	�n�q:[��6֯���7zFQ��C��>A�kK"+$�I��sBJ�����P�G��l��<�E�V����Ӛ�R���7�m�� *���q�e��j���V�P��T�K�ܭ��Wv�
m�l	w�A����xb��C%�;%�瓫>d���Yv\G��J �쌓`�T����9�Ò���������Mz2��Tt_/L��mz����0��h�rU3��a��W�f6K�T������'T�=�g��^���9t�
���X��KV��,8���2h�qI���?ѵ6�&6&��t�{D�oZpH�N�}e��އ>Z�>�MI�XNȉ�����h�#%�T^I�e�
�Sz`�N��V$ė;C`�����k�LbT$����G�HӐ��8N+XP���4c_�E�j�dө�5e��&�b=\'Y���6��$����9lG��j�[�����@^�b3�J����ȁl*���Ӿ~L3��4��ˑ
j�m�(��، ����}���m0X��Cq��ˍΌ���=��k�Fb�H.'�E)|���l^�<�N�6�����X,�e�&J�9�����{��dV�ҟ���������O�8�%�\�b�mkC�-���E64��t��v����M1��;{�>����Y�	���>iV]��Tr<���F"6覅�,W��A�7̮����eH�����L��B^H�?��D%�̕�|�ta`��d?�CY���i�e�~�
w"�����o�Y��>�Xv��r��g��=k�t��p�&�$��<��P.�s�2���@�ĔI���Ӎ�?��܏X�P��k:`fߚ��A���j�#)U��aV�[����.��d04��V0X]~�tW�� �+E�B���:rpY�`���Hi6$�C�w��秌XQY5�y
]6�ns�l��&�Q��L�_ZW�� �@�V��2z�K��,�8d/���^"`E�'���{Vn�> ��p;��Y�ٸ��rF"�V:`04�#��A�P�����6���&��ٿ7��z�3��_�ː�up>'�Ǡ�"�S�|ۙ|Vn���!ґ���`Ň	������Zb���#d� H�hk!�笷!�D���U��b)�o�w��f���)�	|��1�.�ӟI���}�Gz��;_�7�gD�!��֬EqoO;���Q�=-]t��Ў�˿���aR�_v�����_��%�0&EW�ٱ���X����*S��H�h��IM]e���z�w*%��xjW|}��]�����ւ��=a��������}���KP���^�hp�*+�E3<n>�5�����r:�=�^��\*�8� 	!Q�&�W�-�dTy��[�~ �~�xUu�UC�!\Л�0BP��Y�[�����}�4�P�/�p�~��9� ��6`�m�o�?�}s#5T:�df|3�`$m:��7�F�ǹ�D@�3�po�P	@��� ��#f__|8�/f
]�����s�cjc�z�xk��T��5�n(F<
�]�h]��,MBeH+�[-����	.ʅ�Fs9,��Ce"�㣠��+��y��~F�d�G1���Ie�����~��[!˶+:.`�*l�Ѧ%�D?	i��^�T���@I����`]P]RxQFnx�̲��q����/&
���hʄKṅ�Q�tl������km��B��(@�!K4G�ޣԧ�{���;�F��R��ljelm)����4O+@�%�F9S����ҙ�=��xh��}M��<�~Vh�O~$�q8�o �W��s��:��M 7$��'~�4^iQ7ӭ��l�HlT܌<(y�eʩs�c�̕3i.��8�0j������n�/3���DDJBS��C�d�W�o�NϬҁQy:D�����9��U����a3 `��F�����(��­���TE�2c'�>6�5?$R]kf�~��_��(�/I��_e��i����_rߑ�z�;zN��#%2o��+��Ҳ�&!EK =J��1���Z��8�H<��?I�Rʸ�ث�9���������G����ݰ����"7]#4Fм$~�~V3�h�`�d0?ԇ��N��A=.B�Py�k!����%힟s/��8����.г8�ၴ��K��&���6_�V_�3�w'=i�Z�"�����!�}��2�k�� @O�<�z��Dn.EJ�G%��)u�z�G�{�c-���U(��{x-�V4-�o�����-�!T��v
Nk&?A�r}�-�����C0׬�s�WXŃ6
eC8�Q�Ȁ�yu5�m�=\�/^x��ڗ���\����	e�3 TwC;�I�?y�/�ǈƸ�"�Z���]�� C���ڛ�+�^r���K�J��̫p��T�_6����;u6��ּ��������R�8��Dz�=a�%=􉿝����7`�U��}ԃ��nC@о7�wϱѵIf-��,xr�=��[�,�KQݥ�� ��N�K�9�*]�!)>CeyRD�����.mO�ڶ!�{A̫�(�I�L!g���
��-���i`)����}GҼ
|mJ�I����@��#��f��L�(8�>n,�	�L��U�%b����&�e����N�������_h�&Z� Y��~��Y���4*����4C*�fnGW�s��C�^|��Hҕ Y K�N��_�晪�$/W�p%כּ�)`��J�fU�h!i�� ?�W��<��Ct���9�^�=w�;�H�v�f#��&.?��	����w�(�+�HM�Q�_�v�i�>z�q��d�W3փO��.�<Y,�� )�B����YK�,!� ���v7�X�T�*,����M���ͧ��D}��/U���X4�E�+���fz0~<��*8�%��;���cE �E?joJ��2�$G�A��a��9��T9s9�D�#!*b@�c����P�6�䵋�|y��at�CI1z���x�l��.[i.M����p��`m����_yFX�m��T<s���f�G���s֬|%�/��u���oֿ(z�sr�Z�3;�A]-�C�Q�9�/�+b�hg��O�P<7�e8�i0��H�A�+<	E�q��5ir�������9%/"�!�����s�z_�u⊑LNn��q�q����-D��30�,���"�6��:�}�Ǜ;��2:1{^�e)���om|A�\�˶���OS�܍χ�P���v+^)���5e��'�Il$�{�����'6@^�u�����{W3CB�I�e���[�$~�֝R���(����oF��d]ͭ�C����Չׂ��d"y&3�D˨���X��?z�ܨئ$?�z���Cn���H(�-�:��g���l�A����T2��
>�ċ���������c4����c���|���}�@cٲ���L��x���Ҭ�a��mi�K��aj;���j�%�����˘fT��^�B^�g6�S�H{�t�_�����|S��:x!��pe,��� K����6�m�����qF�]��cb���^AZ,L������&N��K�x�hn��t3˹����e�\3�c~x�W
G��3U�x.��Z��o�fT4`���ֳݞ2[m�AtefzC�"���M^w٢��C��߶J�����!}kEh��`�6����L���S6:�W����?|�)-��E����c�e��7�)�Od�����(���1��=R{�ܐiG�X�! �Q�4A2-.FTdd��+5��)	��p�Z+8�g!H�}�ok6��<G �ޤ�	�j6F-g��- N��:����ߊ��d[�vd��N�Q$�o�䁑�,�ڮ���f�0���d�O�,C����r��[EC'Q�
��!+,pY�1��"$C��iy���/H�c�3*H�b��A ��[��)⭤�4�]���(�����Wb����Q4�5��/���#Ӎ՘1��!>�mq�E}!����9nS�L�c	��h�i�����F1�I%L?�o�׏�Cfr�C���n��+u��j�������\&.1e��|Xmx�f�>�v�X���h��Ӭ# �?�J>PIsݥ�;4��ޡ���m�f|W��d��2��
��|Yժ��Wk&NSND�Qk�YlX�֬:Rڞ �W����� ��d՟�Ҳȅ�]Qe���:��˜	���P�	RG��bj����X��!�c�������	���tkj��>x�5����E�j���H��%^��jY����9��������?��N����vk��'I�d�cd�����)��_;�jR�;�MI�T�F��az�k�N�Ҭ��9qj%��Ĕtv3X���eݷꔢ�١+�tAM�8�I���N9�ͻPU�(硷{����b4'���ߣ�m)�~+���;8%���+Oe������K��ޒ���qې9�:D�[Y��$� �����ex1���2�K{v�.����kp�߳�������&�#?��f�y�t��Ig�����׌���m
@a�w���L�� 2���?
��I�"0臨�S��cUS<������{)����4�:~Na���s��E�S����s�h��c����j���Ic� ���2{X�d��1������O�d,��՛������N��Ԛ
v�֧��/"|ϐ{Ԯ�^�[�<��E�����Q(�16������b���*,��k��]$�_:_5e�7Z�Sٯ�����wF#zr���\��A�{�l,���\���k$a�N��[`��=l���y�;�4Brk�7z�����>yN9)<��G<\/���O�b�a�}�)Zt��hSכ�`��,�z�᫬���9��%F���|qi���p���(E��\_}6C�QF}����"6Wo��W��nBĖ<����qV���%Q \E���\ٻ��[��/��"@�D�bPF�f���qh�sn�s9�. ���bn��"�f����k�G����8`v��Wщn���z���n\�sqp�(��8A�=��; wo@��n���mOAcx�T��IWTh�A��ڼ�?N>o���T)YlKfnr6I���)���<}���~�B�s}�H��x�qM�Ɓj�m�瑭[&e�:�I�8@L�]������T�R�=P����𾒀C�3L��Xa�&�ԕ��{c;�Y�u�Zӌ����:WG��:f��6�=�0|�Yy�&���{ƙ�5�P���Z+�׸h��g�LLcÚ��c%�IV��J�Ka�F2zʑ&m�l֯�ǜ�l8��{�~��+�<��x�s�8��6���K۷�A(H���K�1^Y�����%]T'6��y?v���F7#�'mI4���6w0�z��}f�_�����&.)o/�z�Ԅ5�HC��{��ᄰo):p�����<��
p�4'*�/Sۖ���&%j��Z(9�i;�1�u�bj�@�oK���@��F�3
G��]�e��o+;�~qtݮ;�0Ө�H���>�jR�o��}0�c��ڂ>3>ﭦ,ۙ'�B����V�׶PI�S�{Ej�,y� ��^'0��*��$y��<}I�x�}�P�y[���>�B���t��@�͢1��%_.�;܎���q#L����G@uh��6��V�W�x@�y�9�S���&����A����s��ٷ"�u�=�>��>�4�.�*ŉ:��|��KU��f��<���'q��R;G�kʿ[J�T��0�?��<#3��:-М�5�{���>� xL����1�)P�@T�g��w��=T�`��k"��s�IEv��r�@�`�Q��gm�-�%]qR��F30Z�'���y�%�����D�(��1��`�y��/ra'��)۽<E��.tfYָ��K�l'�-�������ռт��D��{l@�+��
�u���0Jb����Y	/�b�ۺވ�K����59}@����WQ9��~����Q>ǒ���4�i��TY|����W�� �U?�����.4�H��	7nJ����ɞw�@����m֌��]>��k=��B;��=`C�Wׅ�n��Ϗ�g���Y����~���2#~��;"� Ag�
K�h�ﺾ�z �����HT���s�I���g5��p!��\[�����hɼ&7��+�:wZ����@����ba>�� ʯ�+�>/I�H�;�[��D	.�˱q]�%��)��H.9�G���u���O7�S|�k�#���M`�ޝMZ�E!9�N�O���W8��VۀU _�O/���;Ƈ���t��!��5�}���wN��h��d����>N�1}_n�E�!/b1�{̨�:O�������(�ݴ\N�E�N�l��ԓ"W4r,��	05��VTj�S#S���ZkwC=!��f�r����:#�벉�EE ]G��rB�%�@�ൠ�V�L�Λv7�g� 5ɚ��wW,�	���,)���]����Q�T���蘴�9`�W� 6b�
,	�~�0 #�%��ІԒ$�2e�r�9ӢF����Hѓ�q+�H̸�1�\U+�f���ϑ�7d��>�蒬\l~H�����.K���J|�|��צ'�\]�ԑ����kVJ^N��ҟ
����=���u,9��A�p* �mӤ7�ާ7�5\)E�����Dø��Ɋs	O|�`����֎�7�ScE�$'{�� ßr��Q���9������]3*���h4�W��R�@�u% pNZd�O`K��bú"9k�50�{  ������Xv�����o�l�mJ�ꮟ�hB����6�x�j��%p�b;β(c:��@�Pg0��O����87�9�~�cs���#<;��,��o�Og�ȣK�m:�ۺJOBk�^g"�����ˡ;����;wIVM~!��/���m�q�'�{q�i{~{�Q�=�HLz|�r.+�xwA��p)���7���s8�3�CZ�cI��{�B��. �* �p[���_�� !<��W�s��0$�t��YTu���fx�6��H����BeW���
�p��Kջ��~�]��]�2��S+"?+S�+Ƿ�퍲j�[�E��qS�1��UÝ�3>��3m2�O+�&t�݄�i5W��p/}U�oF�r�U]�$��ӾA?�¨70��#�$�Jg�b�F�d*�
����6��	|x�'y���S��?�tL�d�.�wO����Ҿ�{�?E���E x]8�����*]G;�sY�n�b�r�hQ�*}�%-1EC5�&ߦ�O�����b�%b��ښ;��|2�/��#�����xc���Þ/u"5����@E*�+$����L��%��r~��κX�-wJ��|����AW��&.�F8�#����C��;�����&��<W8��)1�'$��l�&� ��U�>1$t�"+��+D�������g[Pӟ)�V���4V��س<sòE����~�F�ȕ���*y�(��"�R�w�۠K���������.xJ�g^5BE��]�Ƒ�]o(��M�UL����(�-9:��G�]}�k�n�T�:MGz�ǻ���匹�/偂���i>w�L�7��e��,fUh��z?���'+]�#�DQmK|�Lǂ���>���(�w$�#Dr�m\���FͨF�'�?��;IAl��#`Ț[7k�jyle�PO�������Bk��*V�=�C��K�4�P���,�'	<,���WS�~0���J�)mr��MlJ���`��t�I���)�@�Wx��Ƶ߷�u�ن��r¾�<��Y�ۜt�3_�O�d�>��M-?��dpe i��j�b��:ѫ���6��3႞��N%Y���N��A�X22�[!�.��TgT�u��UO@�TM$;+�%Vݍ���I;��)a���{o`��#��S�n��D��c�2�p0��N���Ϡm�c�fΟ<{��Ď�`M��pXM��l^B�%�L��G��,���R�V��Z_�&u�9B��}oe�0X�[��!c4����铻w�`FTSO���M�s
k���3VD��-�u{��J�1|��L���R�t���@Ͳ�q*�u�o�$a��%��$I$}z`�Cx1rH5��?X��us#i���k��� �e���H?z܁� ���*��_��`r1�;h�m|��Ś��Ѽ/O+X��w��$��kp�k�ں�*A׫@%U��I���\!��b�EG�7[t��mJ��uގ�s�� ����O����H3��W6�}�FrK��n��m�g��� ������$�g�?!���b~i%=,6|���goY�"Na�Z�$C:��XB�fU���	�0G6qVw}�O;��E3���.' ��R_�J�d�"�Aθ�б	�1q���t[���6>.m�5yS�ّ�m�:(7�x �G#�V�4��t�%K0�F*������x����`�����Yv���a���ɜ#�$���D��{-{l��/�i�]��QIsQ���9dg�,o�Ԯ?��L�C�F�gp��!M�h��{�Z���ǁ秦]B��8�A1=nϔD��É?WY�����B�f3�e�Be�՝�
azj=�-�;7�������D7�t 	Ҝ���_��q�D�^q&X��Gw��X�/�7�b0���F:�	^\A��U�V�&�3��^��lp��U9G�(�m�Uvn�*z�#�@Ɠ�o�����i-��ăU5<������z�c	�Y2���\@�@���Z3'U]�O���y�BƸ��{MU3���ޏaU,��
K���桕0R���B�z[=
��T��Y#�ӧA绋��q��~U2Z��$�A��D&�#j�Ը�'�-���κ3D\��j���S���Flk�y�a�X0.����{��Ψ<�Z�����]A/H��_�J�ף`D��2�9�˷a!h_��_����������,�O�V��h
|U�÷GN�=Y�T���tl�*<���o"�n�����1�"��)oe�@1N���L_��	cRǦt�X��ڱ9��VOcG&�Y*���n����urYM��@$f��;�p�?Ȃe�R1�Mda�H~���h����J��J�:�ְ`�Ȭ^h4�\����@�8u��ߒ���v� m�bq��Ή�x�|7&p�k�N�an�M��2~�5�Çb�"4��n�N)� �����.�x/��]�X�@3�L ����X�4��Qt�,
��cۊ�;�� �.)��'W�����̉^i���� ��t;xS��1<}Rm��ҋ�[��Al"����W��P32��3��Ι�9$ov��x\Z�e�3#��k�K���B��{4�>CV�g��
�\�2�~��[*[�����`B�5��R��6ژC�gNpie�م�X��L�����[]vـ5�E���_	�<�K��^���a!q��@���%3s����.7I��A� �E�:�����#�����Ɲ��N�"���� �1pr|*1%Eb�I�΀w��^���z�z <$H��IX�@�N�{u��X��!�6z�*A�,4��^�:�>	B--9 `^�DEn��a�|��ޣR1�U,񇬵��������-�~-M�rJ@���N8�a�k==�-��;`�&���TT|~#����A���f-��p����fIW:��zx�r��i��ᣕ�e���4���H��k]=��4�Xw��@(%�p�W#ڞ,��U���1�䎇�����n���27��t��ܤf�x�2�Ӈ�c)ģ}:IiC-�h:���*�� W/(���oMXg�ER��-����^���EQy�$�>���W��ǅ���{�~O	;Z�˽��0I� ����6���U��T�N{�g#��{��T|gT��ԒH:u��a���jȡ+o�|)���}�v�;���_U�gOY��A�f>�����aiU/f�R�g/>�t^��+
z�sF�5�l��ʑ#\��q������tw�I�ѧRw-̦RsX�/�C�wy`24�bL�6�����6�V%%@ �k�����j�f|���������O�En��4��!+7���������%��$�i�����~��¤�[F�[�]y���N8�,�&���e�K�Z�����V�IS�{(�����j@�?<�;��Sܾ3�91��j`��E�ԅMH������6�o|N§��~>�[[��^��p��f��gF��d��`[xv\��]���9[�����+���/�޴��g]��0R��2<����Q�#���Dm.]��_ 瑠H��E;�H��E���̂��Kr4�d�_wk�N�Q����W�\�>%�m���Wa|�[�}S �����զ��� �A�JM����������H���zn暦qf��!������AU���b{�uwՍ�
O/�@ ��K\�r-�t"�x"q8�kVC���4��b�k�(�:sx�p��wQ��{�,k�.V�W��n�.F��T-]�ĩ�ӗ-�OދV�k^9׸��ۏj�v���d��l��kbV&��L���MO�x8S�ј�2�<�_�\��������j�|���ʽ
�ȹ�=�@������;��+�&�J�٫��n����	]��a9�]K��K��+�o�EzD�� N��.�+�h����E�9J��y7FJ��к��b����N�*"��k�K ���ii$�σ����P6.�+��9�v�+=���V%y�&&�Z�Xz�`%��d�X��Ar���F_R���sv�T��ݨZ+�Z:wdX{{�c�سo���dj�G��ZY�cf�����Xq��|�&�ˈ1C �]�!�.�@, ��x��55�^gq�"��-k��o���&T7&gn�������2 �IEiW���Z�q�-�	�P~-���;ۛ&�9h��-�� �����-<����l
�;�1�jm5;�dr�nڵ��x�]��0�������F�I�6�v+�c��*����w
�i�@����zq�ŷ�⹣c:Ü���2o)��U:�O�^�^q�7yp��5Ep+�2l�,M�p��
,>�][Z�gH�-����\�dŢG��U-�;H�n�M��NZ��8w��t�W��9H�`��4m&IOCh+2�oX4��2k��M(����7��3��}K	���[��,K>�C�gxA��FC<8@�F�?&�1\�C��܂�p�R1 ^�c��r�[vq���j@�8�Tfr�`���<@m&"DjO�!$��0b���jw�s�x;|J����<�ʞ3�>�d�%��]n�W��1��ԬǦ����H�A
���x�n\��Vt��t�(J�e|�����V�� }�~yT���'4���P0<�]zKX�1țڤ�j'2zdT�����Nt��u*D�=�Ujߐ'@!����
��'���CR�"lm�d�c%�B�����(]�q��Ӄ-\,�*����Ց�����;�T�(��q��4�A8�X����x�	�U�Y��P�q�. �4'�q�ʙh��f�\3�8���{�X�n�Þ�r�9�#M~��S�1B�j;�����	�W21 �	C�a��_+��I�M2-ɞn�w6u�?�he�x������>PB~v�t?�ڽ9+��S�����)�T�T�9�l�x��v.��#��������i�I:UǙ�	����7"�JKG پ�Aۀ[�ǩ^��MRJ�C��$����6���,����+�@�.�M
~ܦ�;U�Lj�c8��t?�*�N�����UW�K��8FBI)4��?�k!�%� �"�%B�Ӏ����p�ic�N�1m8�&�u�2a�/�,	�����p�^��H0 �pk�@>�ۺ��N��>7'���t�U�Ao�;�������w�U3��#���eX0�"&$�\j4 ��0�8�u��bv��Vܼ��u�އ����a�M�@G�ts�	��vl�4N���LR��%�ٰ�w�(��pg�Dv����DVG�b�S�VتN2k`;~�d'��b�>)�QK���b7�& $Vq����>Oه���������Q����V���s��w�[�Ƚ�tm�u.�
B�c�fd��zv�;ז��VŦ�c#~���T����O�rFJ��7�L�����SHk���xe���Ρo�������s'����.s�����+��)mX��Q��`���T�вY!*����Cު���Cj�ѩ>��f�����Ŝ#F)mu͉��0 ����mH�
Z�Z5J�o�r2����hv�~p�V�H�eE�VC��[�T�a/s-��zpFyH'I�)�����Va*��q,a�eȹ~^��2 �3�z�.0��ΐ궙^rI '�����ޥ��K�����]llu����?6�&C��W��r���&f��n< ��R�ٮ=1tܿ�
G3R��PM�>hi�1�����	K=�rW�����j������!������7���v ."~
O�q�vxxΣ�I����"�dՉyt��0n�H��K8�t��v�W�� ��X�䉯8�,�-������q�����.hk��4r7͑{��Sd�����:�.��X��Ej%�3,�����5P��
�3��Ѵ�t\�}S��V�C����y�aj ���4�uv�K�ڡ���ʭE�� P����C��|��Kǰ��[�@w|ߧ��OB繬N?�Pۦ���:����H�����q{�t.��C����F\rZP�d�Y���
�����D<"Hэ���ɲ����^�D:ѕ��Lqjr1�Q�j��̀*��߱�}�{6���
��'Q��Lt$N����e&�<b�0�S�͂�%�н��E�:C�ADƐIfu
��-�V�V&���a[Ӏ��,$�n8��L��F�35�k�zUz�JZ��M+��L1P"�?�>`~hL�u��8��U���u�ܙ5��Z��i��|�N2�'��/Y0���c7�J�S#��K�I�b�� �Ɦm�O�E����~�>�����.yb0�.��ʡ\��{��,9�%������rg+�#7TT	`���Z�B�|�ID�Wǉɠ�'�5�`B5M-t��3$:��짔(�t_��V�C�d$�q��ܤZ��C�gĮGS�*f0}�Xn�_3C���up�1�<��v�X$8b�BՃ���M�Ls���S��K��f�C���:7  �D��~�Q�d������o`}�]E�)e3�(cFC��x��Op8I�I�rPO3&��C_[���h�f�< n��h��Р𯆐u�V7��X���)ȅ���ެm�s������A��=Yq����SD�z�m�W.ٹ���.����HI�����r���g�lXR������)�I��6_��;�_�Է=0��۴d�������<�ή����.���ng���d�
���a�u:$a�{)^����>E��fAV[t�;*�i�k%)1WrD�������s��p�svs�-��wr� �a��oY�g��R\o~}��eZ%�,U�ꆼ���}�c̶�ui�p����osA_A�׊��/�]j,����/A����_�mk+�TB��Y��G��n�]�q��ff�k���Y�k�eŘ����N�(ow��R�����:��km�R�[d��J�]��	w�B���T�&����V�,�א��M"I1����*�=;G8�/���H{�T���i��W�ٿ��C0ʃ�XU��:�=�z��5���EOB�g�����~_u�岨	�^]U��< �N\� ���:e3I,9.Ka+F[�;��j���g�,%e|�,��^.����d ��>��ςv��O<���!#�:�*i_v#t�շ�G�l����'}��
�"�G{M�¡���۶�������s�ټ��-J��,a��K����n�͜�*���U-��uW5�U�Gf��md���+���	�cC:�2�-�(�лw�B|�l�4�}��m89xY�0��+{g�r������܂�*�-������g�a`�QR�k�e6��I`5��7&P��A,q���}�����󳎰Tl��n�cxE��],%�,�!�ԍ�e!��"�eݓ�|s̷߽�����c��ٍ��]3�9Q�&��<p,DX�7O�J6o�nb���5��<��� �]��������0w&���]&}{�9 w�l��8�
�ut���n=��}Q =�lg/��Y�rr��߼���vx�Y��-����MjoO�9mۥ������s��� U#��u)�\��vRl����h	�E�=z���vEs_b�'�}�/H5v��iVy�!��J��)�c��y|>YbN�����q�+`ɯ��u��D{���J�vs�mߦęuw��ƌ7�,L�m��FҀ�00ϟC�N֦5��l.��ȣ��s� ��๕L�ę0��.��1���6/��P�*��^"���7ꀫhy6�K�t]���46{UV9����+�zZf�g�>=�>	�t�?�Iw��W3,��ophL�`d�Om�`D�6X��)��?%��������(n*;L?^{q�]i����з>֭��Tu>_툣冶�&�����խ�e���K!P���9���fU.tyڄ�;p��k�	a+�7�	�g�|ģr���+�|Fc�44 >;��yvݳ~�OBZ�����m�����ڞ ���������a=��*���0�t�u�+�,��� ��gd�c?Į��VQ���u�?Ƚ�C�*���%�Z~� �鞶�I���SQtf�ؒ[j������%�����ÂW�t{�j,��_����A��N��%��"~�zϨ�Y=����V�k�j��>� _l��l��k��0�Hl�%��'����:E�c {)�+dZ���v����42������������w�Kr̬��7�S1��mp��x��\��k�4ܦ?�
,�Zʟ�	�O��O-�F���m�����R�~�Wh�7:��5P��4ߢ"T_zL=��T�ߙZ[Л|\~�'P ��G����;J�\����PxfTT��V�
�lK� 3� �vF����f����7@��׉���]u[%X;�5�(�↊�D@f�N�R�۶�3,e=N��Cfl;Fd*:���T��q$<>�'�P���"��-�7�-����,�q�Y�%�c�Q9=25E��ĮS�n�&x�s���6ld�m/�=��&�-���,6��M�tt��A�פ����A5J��)bj�?�Y�h���L���?J�e�܌07_����anT1��c�����{�ry`'��K�i6���eG�\[�<����[Ԇ#��Y�AIq��\t'8O�P�
^�8e��b�د�24=��>Ze�<�}�Y3{����:9�~�v��!灍��1K~a*����n[���6�T����d����.xG]��3o2�vUrK!K��?��,b�z58�)��\�^آ�X�)�(+rK���Ȭ�7iuI���)"�;/��Jr��4b�R��B9�<�lT�Y��i�EuoE�5��|����b]�rc?ɲ��&=����V��3f�)]�Gg[���M
p!���b��C*)��I��4��k*TH-�������DR�,�C[�?��8])��A���d�j�ҜOjfr�~�d�r���\�6����bK�\3mr^E�*'�~g���?+k�1�d��0���`��!�2Iܲ����Qo,�h����^
sٰ��[~�T0yM*%��=���P���$�<+�q�Zo����	Mi�4[^�{�-$��k�HI����gR9�����~�X��𺻮��Q��"a�|�%$�	���(�.5W,�nC�H�������éK�A���]x�E���&����}��s����,lY2>����)��ͭ��N�l2An�U����"s���h������Z�g^pu{�Q*��%����A�2�g��[=�Ӱ�X�I�9H��{ i��$��m.%a�ܷȱZb�i#�F���FF-9�d�-83���7T�!z�Jd�|��q��s���2���<\GY���#�(w�lpt0 v-u�L����m�oC�k1wL��r�*�����b�Iփ����M����Dt�C��9Bv�7@�R��~[q�eP}����u���"X	�M=��>D�iC�1�ϱ|{�OE�jM�)��V�1�5X���ke��o@MVN��_$�z�M&�����X(P7ϚZk?�<�d�lܵ��������6�!-��ߤtƟ��$�em��-o�>��.�ci%t0Xf��M����#���қ+���qZ�:�H���Ϩ3;�:�-�#����3���+7](�L��vsncyb�0��~��\�'9��Wtd��i8�ʊ�C�aJ���r>��@{-�/��+�DSA�k�W���v�ϟSf��U��<~yu�@�0<%�߅��C�phE��1�|J;Ȟ��_b	J��.���2�����9�V?b>棑�<8!�$����c��~��BK&�x�3��A�e��GV����L|��d�w=fD����'��ܔjd�*��!�#�K9��:�D� c���&&>Lq�b,uۃ_<[Aև��f�5Bً=��ԁ������$$�I)��fJ��p[dBRH1�F����(z�gb���?�ɔ��3�|6L��	�kq#Y߀i`��d�Y��sH�&Ե�a�Fn��F�s}{�ZUf톴I��� �[9A~��A{��Z>���SwҸ@	T`���c��-�`�XC�
�� ��<�U��Q�}y��PSG�UW�h�tZ�T���C�:�{ie�0e��W�n���l>6�h��QS�����_�z �G��4���lg9��cĤ쒝ђ�y�)#��e;v�4�����u�4Sr��q�f���SR�O�l�k�C {lq��p�mW�g8㽄{ӑ�D,�����9���yX�OA��V�8/��%�*�3��l�͘���Luȝ��o��?�ĔΫ,Y�.�}����k}��<X��@�7���w���cZ)�X�z�
��@��؉�*ڀ��� mm_lN��w�Yw�)��Z��0�b`"�|z��0�~�ew��p.�Շ��)�����l ��~^��	@��J �,+����Wp&�ӛ_�c%SD�.��U(�*#�_n�)��aS߬Tq�Z��,	��#x�a�� �iq�C%����u7b�%fGl1(�j����w���ul��$E
�5ƛD��y�^��o7����F���Y׀&o��z.jtlꠏin������3�X~5���>8)zx�jv�-{Q6��-���u�y�$h;bZ�&��n�s�;n��U{eq6��L�T�E8�p	�_�}�_8֋�@��_OI��!8_�Z�lG�jRMQ��K�O�!a�bqg�MtXa��=quw6��@FI�ju�����:�#���gm��˹�.��,P��e�Q�f�D�3�>�_d�'��1���$���2�3%~�'g�O�0�	���(>TobqS��^ Z?�z�:J�H��x�R�oit�Vrj3!��2z�#�~4���9A�rx� )ƀ#bFPh�	�#"$wv"^{~ ���h�������ޛ/���ņM&p��-��Q8I������&pF�������_�P��޳�}�S������n:W�D(3�ܻl��sŠ��#c��l����
?Eu��~:�6ޮÛ,����r�o�{U(�Y��z� ��R���tD�p�l�K�tXX�8��FnxFoK�^��o���5]��	�mt�����swPPS��6���lyx�����UY�G�E=⁗��#�g��2�N9��.��Nk�U��e�U�/�����6�s�{���-=�Ҙb����#��0�8�	h�01�$�[N�Q��U3ܴ�����bV�u#qe�s���qǩh�����m�
�&��r���L�RTi�`����k�QU}9��{�*O�+XoE(�#�';��w���V�cC�,�'Rv �#Q��jh>��<Q1���Q���N��)8m|�hO�q!�+����7�:�s�N��;���ߪ>���G��G�����wR�k���E�l�N�A�
>��x�X�������/���0���������]>orF��e����E3.l"���(�FG����������\m�V�����[��żk�-Aǁ`�ͪ��y�Xk	���.g��mv!QJJ��xR�w*�R�	���.:Ί�*C�dϟ2�X��$��$WL�m��"@kxHÜ]��ê�^^���i�u.,qq3�hdAU�v#z�Sў�D�ݯ��H3M?����O~n���/��~��6�9ٳ���E�Q�e�����&�X- ~ԅj�מ{M/�
|@���t�<߀��~� ���;�0�iB���ckw��&�J��0�=Ol��k`׻H=iȕ�В՚(��)�2�o����Kzܪ�L�&�L��iM��l��%+g_�M��T6FN���=�K���g�1h0H��ឲ��h�I�΍�o��{���1:� MiS��Y�s�^�����M�7+��@���K�ȩ#Ý��.��ӱ�+��� h��gcؗ�ǖ���9���崘�^&��~d�x~FKkʝx�y^(�T|Q� g�_��?y���vX��x�»7�.e�3��`�]�.��Ή�s�(w@���x'X����q�#u)�M���jm!3����k��\��o{�J�~��>�.�RڣW�����5OIń �h��;nyL�h�p�]U�`~��S�Ј�Z.�= �΄�]��!�K�76�I�8�7�a?�!Vu�k-5-U�����W�|hL�d��OR;'/�e�شWI	Mo�����rj����c�J�a9��3@یiYX�;���uZMW	��:��4)�sX�4�/�4y�y����.��o�,�6x�M�u�`͑�c�/�]N�K�Џ�I�M%��x\������ �e��lK;e�6�߂���������%Gyj;�a4Q�N��3/�gW�K�^Ca��'�K���T2�� &��e��d��k,��2�Ga#Q`��;�-Z��OY�'�V�+��X�$�F*��fϮAf�\���$�\�%���9��B9� )ٞ��	\�2�t�#�i��.�u�^�֭9�	�;��:E��]��a.�Æ�a��-Y�{��=��Fj�/c#�������1��|�94��N��:����?f_�qb ��}����Z���FL��ړ�f<�j��o�5+̢e��Guݞ4�mx����C~?�F<U5���D�p�����H%K�Q���)���g_篙A;�*ד�����C��wfJwlz����VQBy����n�a@:�}N�zV��G�����9P��Z�kl��B�ሪ��j�)Μ��￙z���)��f��VT�g ��7�9�c��8@�D(1?��&�9����l>X���TV��t��s�,�k�d��MZ���ΐb�y�ug�I���K	�����U]_�����Ћv�����p#���������s[�5^G�,�_�U&ڷ�"F�6�����Z���B^�1�:�%�7����V����߶�i�<ZC--���&U�nu�R�;�1���a�'%uMtQ�i��K���b���dDi�կ����W+B�'��DݔV�������k:�!��v�Y<��y�I}֋��u�6�(t�8-�����ߑ��Z��3�JVra�������FK�/��j@��k�c��:��Q'`|��8�O��3W�l{���B�$ƭ��9X����_����������N+<�w����0�q�]]I��ZŪ8z�����ډcF�����ցQ]O]�1��W��䗃c���5<�Op����LA]7�t�ߤ��('�g�:+1;N'���D�d����אT�f��l�NG8~��3��dVvKti�C�mM��%k�󄞗bJ���q-�<1�l���1I�?C�8_�*P�>���������p�M���LT�Bc��Ds���H�a�9�ź��P�&s>���l����ؔ���䏡�$*���'�ؚU��KgM��(��+g���^�e|�ݿ�ʏÐ��5[�:�zvS8Z��nAʧn�<w�p9�>�d���u3�DϦ��/��4��#V�σZ�[��9!��aa!��h(��OG��[l�V>�=�sk���ɖ��u,�ạ�	����jf������F�H9����p.+����������Fz��E�IY8*w8�c�.��'d���b`<�`�i������(� ��6"���:����k�/a�R�nm������;,������7���;�u�e73��݈s��=�6�*���tRܦ��6T�׹�\��	�h��G=L/���g�0�R��6�}̵8djQ���I"��ݓ����F����Pf�n��}�{[c��Y;�nQ�l"Œ������B"�&fO���M��-�v@��y���w.�K� wB��u�e��Ru���� G�j�]e�לxܺ�\��YE��5�q-z��	*B� ���bw��&���`V�?��{��!ߝj8����#����S5g8�x�����l��d�S��"��"vڶ����t?��S�,-��HW�E[��v^�����_J�V�E�1by����%�)A�2l:<�����]������}L�S����8�c�����Ve@hr$�٢͡���;��:��^�*�]��4s�H��ҵdo���GP`݁Y�Y�jA�Gc����Ư�H��a���,��~���G[W}`	����O��Jt���U�"��X���s�`�\g�X�!�sz�����c'UP�]铘]��A��ki4����W�%��j��[>1� -��Rt�r��G�/�J��x|G��F��r!{QOG�VCy�g^�<��C���xM��ҳ���:ow6�	wu�K���TIۿ�8N�m���~a�7��h�0hR����{������U�L�-	!}[�x�M �G���܎m�^�� �q��|���F�|9]�\�Z�[������ �m����/�/;�X��`i~��F^���сƷ�l��0�u
>2W���(�l)�E����myа͕�o��
�`��tW��;�N�T!C��ONm,�ܭ_�4!���PI���%����Y��!��W�J#�_�`�/�:���*��y�	6���ܡ�͘��l�A��٭��aу��%��Lml�
�	��\/�Ȇ^}�eeJ1�15�j%�>;woA-���@L�^[�����b�*Q���N��Dc*�����g�
��i����/B����6�?��K�v!Ў�a#�{��s������0��GȂ8����-Ʃ1�r2S��05��~��LG�c�񢽿�k��67����׵t2+�#
�����>�����,�1��cy�����ŻQ��9'G48^��ev�)���4����/p���f�\Qk�={p%��sgk�?���+݀�w������k��Z4���dL&���D%����P�J���ߍ,�ܷ�q�����V^��+�M�E�YI��R_K�!���Fh
J���c����|@s�QJ�>�1�Z����	�̔�����|�c��~��݇��:���22��)���Yt�pOl<X&ֺ��B,<Ys�Sdv�X#�o��,��� ���v`r�b�
���캇��6�W/���0�e��yF����	7�nqgSݰ�nw����Ҝ��L���D��9��w�vl�kb�$6�["	��!��r�X���l�p�ᤃ�,�X����׮�0�3��,��#DV�8(��k��dᒚ��q��� ���)�9�
�s��	��3NuŮ��P���ߺ|'�h@mQ}������!g�B�
����~if&z�v��* u��X�8'f�0��i��LȤh̎�T]v������2]V;u9����W��X= P��`�%��YjS�8���o��zU�"s]�)�^7*��3�;��D֝=�̡G-���_�d�%���An�2ܦS�+5E�^3lT|��8�h�$��	2Qz�4�<�XA����`�����&�5��%2�!0 &��$�����u~=,��kۭNB�`?�ȓuDDV���;�(�[�	@ �fg�v����<n�N���U���1
�5�Lb��s|X%��,a ������1���e]���Y�_r<�{$�.�GF��Nwl�/W(�x�@Aˌ�!�pSU��J!����?��Tx��=�e2o<B���pT�%�O��p�0b��;��"��b�4�.$+��1����~�*��߾hQ�_����w���ci��D �Ҵ��Mr���P-�	6��ŀ/�n�����bf#�h@b��%�BKE?:�=>(�CZ�Eө6��J���Nz������JF�F�y���FW����Mǟ��ǌ�g���}A�����R*j%TBo܏�@aP��4k̽ʂ	A%�Һ�-D�o�h�N�w�6�}c�bE�
v�'x�M�#��y�8�.�l��14�F�xV>&|��&����d�D�Ǹ������e���)��dt�"�����+/Zx�C���H�mү����=]���1uފ�C�r]�AHW@	��!��Vi.9m���?��|��Ioą�N�M�5��}�s�+�NRo���qV^~]3����ݐ���N�Xқ����۪�W���/��hlr���@>��v�bi_GO
��9�5�Ep����*��ߠ'�����F�׼�*֝Zf�T�㔌�;:c �с��{�i�����f	�X�E�c��Y}�9~�$�q	�1�I�bt+h���a�T"�]]Ch0?�����M��m�d3e_�LW�s$����MBvt~� �E��L�c6b�+WY�Ǝ?,A���|��Y�]�5P��5�-��������WP��u���qt���/��RVVrwʠ��z��wD�ʆ��ps>]��a�|��(Xt�tˣ�yr��C���u�FJ��͵F{i�����&��*БU���|J���C��Gf�����%z�Cs�ã��9ʏ&��Md	6����e�q@BA�9�&�����X���`c��M0]HX���un�����#�=�l�[�'�p PWn�� ��<�ޞ�@����Ѱ��5����z��M�dk�;�y�P�����m�Ռ �v�+Ov�yGdYU�ߜ�K@�����;�
��cw��=���̧? 55rT���������!'�GZ�e�s�k�2�7�g5b��:ͩG�u �r��&!���~�괜�s2�AÆְ�m�	KA(Ye�O�w��u�` �XPǙ�kcm�_92!�v"��
��Ӌ���y�Dnj���0<��LY1��vn��*�Y��ReC��oŇe	K=*9'��^�b���/߭ܺx�(� �Z�G��*$���;+d˂��>��5tl�+p�IK혥��N��3Nlg}Ioif=`����:��r(�'���-mlR(�:��7L�A�<��־c*R(k��5[�ߙU6H���^n9�޻��tj:����2Y��x
O���o�lݙ��b^L�����گ���J�`=��,W3�{��g:��B����9�0�P�'Q��Y�'2���I�~d�?SBދ5�e��10|�R�F�#�h��x���q'-p��b#�I�gjF��8"�ȓC.,LSzV�z����l~���Nr���ڰNB�ghFN��ǘ8g!I��z�'���P6� .ֺ�>K4����H���F��� N��d�0{��®%^_�L��;8	�DCz��mt�|nД����<�u=�(��,��xj@!����,��D���%#��t�L|Ř����%�96q[�i �*�����Z7�=��/�A�Z% ��Z�0e�j�*�=h��'Q)��P��=^�
N�x�tE�n|6c�W�ٳԝ�ؔ�e,,�,��4�4<mF�*��7(mPW�������Ž[�C ���wŐ�Z�=�d���+Y2�BBG[��qCh�oP���o;�\��aP��IG3�����w.�`E��;4�5%��K#G��ǽ(sz7�������M>���=�Q�����|<���
���;�U8ܶMj�����-�֗������{�v�E���q����v{�����dF:}\-�So�j��L��<���i�d��5p��
�����!�(�<����8׿��n��+�P$��	�����a�?�4A�YQJ!Ӄ��z�~H���sUO��ٝs�l�Ӏ�RǶc ��|�G�m~��K6	�~/���
�B�&�|��Ռ�W���=��Ժ����IK��WV����g���g�����Z���A���]$��P�
Hnk	��yAe;�_���\0pIniig~lؿ����F���"46yw�Qy	Py�ْΕ�
_��'�v�E���~�	.ʅ�����>�U�Lyhx-l�w1q��eA���F�E�舂��$�����;�yt�`s��o��Sr�J���XܘN�H�gsI/_�_�Sܪ��=�,��T}j���	[@PD�E��"��DG�G2�ԒY�`?��d���I01���0��̐_���#����$��h�x�1�0o��ɱ�l�X%Iz��2ǿ[�jU�V��˶��� �ՠ����9g�En���G�g����e����Hu"m٥��{uy�\�U�L��X?�d�aT��/u�|i���֜��JQ�:Xz�E�����N[��c�<@g=r���{䗾�C�˔b�m�N�~^rm�3 ����������+��j�+2�3���<2��0d��웩�qx%7���'W��w*,��77|�#���誨�����S5�b���ϓj�ar��c�89��b�XrH�hpA�H���"�6E�����xp"�N�_����9�22�@&��{�p�h�W)QT��fP�I洫��r|8��	(��*�Tr�?c��9��^5�>���R��XH�qhXye`SxAW�7�W�k����������7:��k�K��_t��f��AN��@Շ曐�P�ħ�jzw�g��T1�e3�H7˵Y�^��m��Ʀ�O�ClY=I~�#w���3��:<"�aٷV�o(�n�[�ѫ�ѹ;xd��Rd���X�:>|z;H��l�\�'8$d=�09Fؑ<M�2��{SW�ὧ��:oG)�N̨��)I������QYz��)�F�'�܍�b�?�  s��RBq��\��|�|U�[�'�rp�m)X3�͸��Acl$�e,{q1�F<Y�@��,���?	��Hv ���P�g�G��EV����������S�r�|}ƞUK�s^����7�U9]���Թ��=װ�\P2����jl����9�-��E �,�[�F�Y���A�m���8��� $����l?�N|A�+@VRH`v���2>)�H��5{�O�y�����+'N�C���Zϰ,~�tn�̱�f�C��B������� c0޵c�� ��w�|Ɔ'J�b�1+����BR���8���ɘ�jv�3b6^_rya?��=/���Y}x������4sM�+�\(P9�=�����)����z��Kd!����F�` X�^X�Y
a8����}DD���`6N��J��e
�P	<a�*���9vix6"���UWM��`�s�s�b�u]?�V��Ee3['��
4��!�W>��34��b/�K�xJ�����d��u��U�]�AO?��N���t3Δ�D�N�> �����{vC� Z�/w�!z�NZ�(I|8k�֙�_Aoq��rG�KUoj���Z���o{����W\ʎ��HXB)$8��PK`e�4�1_=�_vѠ�b��~�J��>�J�?ѐ\�K�ތ͡��U	��7�0Ye�wp)�ä���݅!2,��"C�&7Y҈�G���I����KnJ��� /zz `�2�䏢#f,�0�w��u2���$f����CUj��z�氿�*���Ѹ�١2�q��8H���9�����n�
���Zz���V�Ρc.�'a	�|�q~K���;�Z�e��^�ehV�$e�A��&�%����CY‽�����W٦�������S��q4�(�-.׻J_c�{=�7{A��9)��K�KS���İ���%�.\١TT�ˬ�� �_�a b�`Uw��{���T�9��]��N�8�jW��z�c��iS��&���ٔ_v�{=YE�WN�{��	&�΀SP����f�WL���J��P��Ʋ�+]L��ƃ8�S�0�Ç�Ma���{C(L>4�
��/����֖���n�78�����M@�6Wa������F�D8~�,�Ǌ�H�M�8��q��|E?����� G+�,D6;�d��V�{���4j���;���M��,�D��-��^ޅ��{a˗�����Y�x����}�)5@�$^������U٠�v����:G�M]) ��6�h�ȫ����)��{��zVQ��x�I���U�h[�dk���i�l�����H�>,?u�UI���t�)j��e�~�/�w݉0m=}3�X\j�����5��Փ��nl�ʁ�6���4�#D폾D3^¿�N ��O1�r�4VB�^Hc-���qԜӺ/�j��L��#x���ȩV��&��.������9�'���Ĥ�gp��)5�O9�b�ȑx��;i3ܟ�F���	E�Ω!$����%�/+eB=$�%�K��S�[��q���"�V=���#Q�J�2Ek3�6��QoS!�.We"<��MjU��(?NER��v95�)(�����EXsa�oEo)θcYJe���5�1gJ{vY�B�D�*�*{9���ֹ5�����]Ý�[��}�~�'Pg���Ej>S9����p����㻉�{X8�"�E�1U�ak9�R��1bH ���0��wJ�[!�<�3��_�9��3�����ӧ:];�/�����`���_zm%�[���ơx螕]f9�򓚧��Zo�A� ��֤��\-8"n6�g+j�ieI���u-1�i�
�J^kA>6\4C��\~�n��.ׂ:iq�ȅ��΃1��=�4̗֜��$���د�����?�N���|�<5���`�~�a�ȇ���j������8=��+��PE��m�E}�e�br��a��Lϩ��T�֑k��g�=�d�Jp&�`���*�'$�/�6�Cu���EÍ�N��9-P
�� �Kƚ�C�ʶE��M_�j��$��Z���G�*n�Z�-^����MۥXMf<Yf>��I5�\�+��tq�5������IS1Q�4�,���٧�N�j�MفB��;'j&>WaP zM6Cg�"'珖��d��V��=�w쫕��8m+[#�t �r1_�4H��#�,��x�OX=}|���uB�K�m�Vl,�D���.�8<����驹aAT��~4��%X=:�l��S���Ձ	VfZ;J�;���[�&7�ΪU�-�L�1��L�Z�r�Bψ��})��Y��bxO��SbUҔ�X����,<�F�EH�mS���?{�`�HM�$�[��G2��`�[�Z�ZA�~
�*^�s��fq��h<��Y"�>Ǽ�h=R�̮Zz�{F̭Dau��>ݎ�:)�s�clP��H>\����G�r��(�9ʵ(�h	wG��(Xj7�^��H��CVD� �}
�1�!�j(A�=��H6@�&���bL	���V���;Tͻ��1��=��JL�����(?�7V���e�L�f����@&sQ��Ά�v2np�S"ᰓ����.�T��.{MJ�����z�i+80�/$\8ܳ�s7f����D �NJFQv5p�@gR����R����MAo�&��%d/N��Ѫ�`�}�3Z�I� lHiK�Ѕ�����R��Z�������q�ͬc��UG��<�U"�6��
Аڬ9�v0IX�0�GH��=/���m�"�D!�OjƏ�\nuɃ��̠�Ц���ǖ~s:�q�fA�IM��Or:N/�>ad�+>��M�sΛ�����$��)��y�v���!��}O�+]�T�X��w���uk��RR���n�h��)Pfqt��J��>f��$�t���sf� (����=B0 �����#>�w��?g�2���Z����"�������4�O�Ѩ��'��d^�%2	��]H]���H���1�o3jI��DÎ{ρ��N�n����"
?%�ZeO������L��7'�\Fl�ͨ�P��^I#ɾ�� �n�������ͧ��L\H�m��W]�Y���M��u�4M�c o���~�N��� �T�hCAn�,F���d;�U��iɎ�����i��#ℿ��)]-�=�q_����"����&���(N��|A��M��vQ�`�o� {Rɓ2���7��lX)�D��3/� �v�E_nQ����It�<�h��UA�5^*\v������m�V)�I��P0�pQ��o��5f����P��s��In�x�ď�l$;1�<�8�J6�Z6��#_�ʫQ�W���_c1�q�sUms�ߴQz�r�Ꜻ	����NP�ԉ�N#�7	s��C����N��V���T��p��ޯ����w�����B�Y� �x(�'{'�V�#��z۞(c��&B�c����3�}T^�Cd�z�4=���_S�<a��$[y��`S	1���� �м�"%�����Ҏ�j_N�_C͡;Tcp��@��Nklha0)?�H:H�ʅ��|�=�ǎ������d��f\��0�gz��Y�N��%�;з=F'�#k����	�=oG��L���X�Ӛ�m��8�dR\2,zg����6���@_��m�S������1E��CN�
}|}!�c��^納���D���E�GYWl���r_�y��6������z�>(�Zr#@p<��~A\�{{�q |<a�L���v�Iz���F>o��3�<A���}	2�SSwy{_7�ga�5/RF";��^Y��nG��Gb=i��@�*V*�yX:-?@�G�:@��k�Ồo�� z
� .q��yJѓS�񯴘N\~����9���( +�A���)ō-Qe��0�+`,��a�k�1�x�? ;�� ���N@Э�P���|;��y�:�k�����.��t��>���f"܆��k*����<U�9]�;�6~?��T(���}���Q��Z�2����8���X�k��ކج��D����p�k_��?5���A�2t����������;��T���,ά�����&������������*hkp�������G���}9��p�D�o�6���ж0FQ�� ���6�5��{���ۍ��I����D,�LY��3o�%�;�yO����Q�Uo�X(2�\l�l
0d`V��5�F��3��W1�2ܐ��T��$��~�aE�O�3��pK�`�O�v�qA��iG�RV�Q�#��ۨMއ���)�g#���{-��߼�����ݢ��F���Wq@�4�&����B}�^�����UY{驿3�� 68�[0��ٌcN䒷��+;�f� ����H�ސ���*�3�𴕙�sf��7��B"ޱ�p���@T@F�s(oL�}�����fʾ���4�c������ƙ�ь� �@��	�)Sރ��qǃ�4��U3����BT>;��I�b1�$��gtnz��%q�r�ƭK��P�j ����TϢߺ�_U��|o��m�w�m݅q�Q��L_*��3�A[��WPo~����Go���[w�2�X��
�c$R舐��GK��C1 �{}�Rbd!��4��p��h`\����3P�Za�d�R����G|��u��Q����@#8�$ T�]�_T*�bV9�d^��� �Tc[�^�);]t��=O�ףs�E�G��fb�Ǡ� �����_��5,�#��_]����Jźl�0hk%Nde���Y��z�:}��Mx��.H<��6��(t��^�����qĹ�N���7�c�ϛ\�9N���;�91Q���/Ir,����Pq��#��P<��9C�*�]�YP�k��-����Ϧ�rE�l|�dU��$�]��60���޴{���ǓtRU��r4\���.�R��#�}�$Ϭ%7�^t&�$�� �\@�N5bsG�gJ��բl�>���/��[��S�3���{(�3�_��'e���TPזw���1��+}�� *����x�s/���ti�[M�GB��ޕ�_����⡬
3f�;�6zF��T�a?��cW2���G�˵:�+�׹�Jذ�L�k������Ϯ�\��*t��59�{1���h�5Q�S��P�3�>�鞑�Cwׂ{�|�{�B�d���,����r_S�
�pj�賒3K.+k��K`�<4o���Da�*��/��,��t����拰DkU�t
2qh5��G���9�E{%(�������Z�����X�"�˂1f(��N+���KuA����[��ŉOA1u��O���5^�ˮ=�!6PZ m�S��f)��-��#Q��'��b�cW}
L���@��W��hl��p횯���Dϖ�k�8��X�2(c�T�����}ʂ�PEs-�X����	Ɗ>?�<��Li��޹�fUW�>�ⷨ�,��w�ku�K~k9�Tc�s4jom,���\������'�	\�.qӺ$���B���<N���c�.AI�c���V�AU���~����tP(ºv�ǖ�5���G�8���_�fkqnR�dǋ���^��+�0��������W��P��k�VN�m ��y��q*�Q����oQJXh v�dT�5Yl�*�s?�j���>�����fI�|;����s�,�
�:!��Go�Xe��산���ڣ;ͱh4�
�ގz�~��_�,y��8�?`42T�	?3jK*y\-	T����Ų�����%1�����-�b����q61k��Q���<��b���?	�x�֒C�i�R%j�� �&-<Y]�˓�mMJ��?B?�����E�������l��!����Q\y�9j3���I�s)u�m1�DP��/���1��������v��x��z(���楕e1�������	,I1Vv˥��6Ӭ{.V�Pv�P��A��n��m�d��`s�Ϣ8�uX����8 �p����w����Λ���%�\f�0��VU��h�'<�%ݸ{A*@�����\�wd��}����oF;���UOp�҆B�eV��_h�
���`a���!V�>#�&�d}3�q���	ڷ�{h��P�_�G� @u-���~�����6R$�L�j3/�,bxoa���͘l�9���T�3}�}���ӵ�u�o���Ω���l����v/)k`y�N����1�pCb��[���<��́�T��C�w���r�-���؍��!���b�����Ѐ+�0 ������%�z+
ƘN\\'/�H.����J�B�p�����z���	���䥭L@z���X�e�s�ݾ���j��~̷��To�� D\�_�P)8�A�#A�g�+brJ�Ef`j3�R��_a��M��;�?�%N�Y��M � Q�.��� y��.�5��ٝM���
���%r��N2�O�mt�9c����B_y�FX
tzm
��@Yy]�����D�v�|:��[�&� a�ҳ�?��Q���Gmu-���H	>,]����B�f�s�>��c���8��^]��&H���R�ќ'� ��Y�0ն��D�Ijq�'nM��+�Ǚ+_P��pUX*G1���\Փ��PV�K�Y�0�fA��'���)�X3���<�ي�{�{�﷿�l�Y�����#�?l�갯���c�=9�m\�q�t�5)r�{�i�Z���Bø�ͦ��N�ߡ²�ً��6�HF���A6����8���������oPf��NtT\�D��y iK �R\oi����z��w�����cy���^��sm�+��5��̷S��2�!��l��������|\�)��"��:у�C���t4-G�ie��ԁ4�:xA�T.c�ô$+#��=i���f�����v��!�{~ѹ�#���m�,a �z ��!�=f��L�k�S�����A7O��o����Y�͆l�?�����R��̾�ji�S|���Ҁ>�����t��3:O�_ �30��# 뗾H% op����m0.ږk�ܴK�Sj ڊˊrQ��D��̾�+I���ݡ��ofa[6���<'�b���ѫ֓��2�:P�ؘJ?����G��;s�8#���w�'E3+c��������,(62�%ۋ�TT�c}�h5?-��f:Ͱ�F��x��y��ڊ�Ո
9�J���.	�����Np��̰�{*���;cȢ40k���d f<lX��?/�zC,ҏ�%�(8 �6�@��6f�F�:0�V* �:1��b̓	F6�~͈�:j�Y���יx�:&��	��A� �A�\
~�~���M��p�tQ�'(�ז|M�/Y���O�o'��**C����D�+pnɖA���^��JQ�W�*��(�O��h;ѣ�2E�T��vW�,]��w�}����0e$w�)���ϭ;bʪc��Uv�-6˅d���H0��� ���d]���SuO���\�vI��,�3���w'�� ���ؕHM��wъ�p��l-2o��/�z��Ӆ����/Vwd�}锾]ZM{׵�,]�	Dv��׎�ce+���bg��4��R��"�&��^���')���\��8g�BE�����Y�1�T��Ѹj+Jɖ"8��`�Î"t�l�V`!<�&��DT�~��k�6�'�*I�	^e��{��d��U���o��L�B@��ɯ����d|��CZ�8�^ĔB�5�����z9���>;����T����|p�a͘�j$�vx)`��ǠKnĔ`�����"5���u9���,<3��x��rag��suo�a�e��גU������B�eN��8��l2�a���� ����rB1������Oڪ���y��ŀ��!ܺ�w��,���OS-#I8�8���|{K��(�U5q{�� �X��w>�(X�&�֡+ycnS$T�� ��n���nG�������)��|%���$A^ݢ�E�k��x��1!���e�
�����JE��e�_,���ߵh�)�9aq�IR����	N�T�uC:9dQ�kT�1p6RJ��+�$����������>�Ǧ�L�-��`�V���%�7R�P���K$�D�|�qm0���FkQ�&u�����"ճ]�I�����R�±����L�F�:hb%��
�;���!��,C��秝�)*���:;�h�2ڬC�&
�������������hK��u��k(�b�rZk.ܕ2����� a�m�Ͱ��w��=V�8��q��ͫPb&�7�a�V�B+����4�����?��z��`���%L�[� ��]0h�Jt�t;�]�;9#J�R��c.�-mk(p5� ���7c�*T/'z�ۆ���qAKpux|���$�S�1��k�Wd���C��7m�'ܝOڠT��/ޚi	'/[�q�_Z^�x��N�1���S�.�RӦ?�
��Ib]�S��j�[���˖_��;����J�̏HG�(�O�5Uoy��V���1�cP+*�>B*�8���,�dԠ�&l��]�}�_�m7ayB�=a}��|sOJ�{3mc�%*B��U�kU%x&kn��_����E��ׄD�/A�[zAZ���EO�9�2=
;'Y��g�Y0Ϸ�#�P�|�bҭę&�M��tm�63���ʊ~�-3�Gv|��@:L�z1���	�Y��A����c ��	��k�}T� gߖ�s�=-�����t�r�*]�ʡ蜹w��j��*/ߎ�K�e�5|O��I��Bd��5��y���AU�;�:K�1�-op;5u߳k��f�^5؝���r��35��Ů�)���	&K�=HC�N��K*$_io�k:H�;P�*@{� f�K_R4��Z_!����Ї�(@�I�Qۃ�����W��Z�+Ϡs��7lz<�Wi|%�;��K�0�M���!+9v�>B�ٙ��2^����M6��{)b�RX����g�#�M��(N�J:��%��䞓DD�Sg쨢�	Vg�("� �<�~�N���vl��N`,8"�`�z�0W��o�Ύ�Ua �p/�-�}m������������M٣����tbu�|����f��=��ୢ��D4$J�IN�KRk��/�#s����&���W��C�Io}�8�<r�-Z��j̷��¬���<kX��͋ɹC=y��"��e�"��iŰ���g<��g|D��QVY���NV*�(f³j���D���y���9�Y݊�Tw�b�W�E�D����@#����C����P�S6+�P�:�\W"���	�j?�:o��m:�M�X>8�$��M�F��(r]��Cd����������X[#wh�[�U���ٙ�:�(�F:��f���W��o���\��1Y����Mw?�B�����<�~xC�IA�+��4\���Sˀ�
������L��.�Es_���~�x�P�w]�7nd��"[�R�K_��DG�����d�3�D���n����8��u$�jZB$�"����؁��9��~j��vT=Mי@��c4%n[��ye���p~_��yy��k��\W��`! �fi��#�Y{

 I��j�f}_ºpV�w�|>q�Ѽ>�Uڅ2�7�W����_�-��oEJ8�JrZ�S2X��d������-�T���_;����ovLCBk����̱:����%2ϻE,�e#��!����k/9�R��_�ƽOJ���YcFM�y��B�sȇ���R�����e�ȃ�U(�a�r"�%�Ne:�I�o0��ɱ�!R<K̗{II>`M�<l�9��t��-	��e�9a��}��T$�2G^��?���/'�_�|&�ԋ��/fa�>i�e��?����w�53q���%j����C��X�� e�]֘�P���1��s��ua��TP>��g�1���y�#۝��n"��_���x��`T��q�`�Ƕ!���(rke �p���	����n���E,*�<�Q]���p��\ ����у$ eN7N%��`��K[�Q�j5����V��-��÷u^���]�!���DOv��α�V�0����Յm�iT"L:�|=�k5�� �*ǜD��q]�D�-�B{e;�VEkd<�sCp��Cix�L/ܘ�RYMw_ś���r���X3�¶0:�ӝ9gI���>�����G�n��>z� �'��59�A�:@a�>)G�=3v�y	$�^vP�1#�0����Z��$�y{})��r�Cap��7��C=�Q��j�����>���(W��Z����X��9B���<�ВH.�!��*&e�Y��i0g��B��,��Re��di�B@����)O�4&������d?v��P�+�	vv�"����t��&�Mp��ȹ)\Ge���Z��Y)�Bo���&V��P��	�c�����_	Hz�~�-�W�JEt�twʽ]���	8B��P���}�!�O�0��ʒi�����c�hY��m����K*�m�E�P�N����ldX�V!n�r���:*���w}�>)�����{@E�%���1��J#]x*�ˬ���E'J����5R.Y�����RnN�z�6��ey�Ĭm68 `�D*�#vy��+�t}�Ϙz�����k�]�4�=�o����������fЉ�\9�\₞�˂�],�\���m Q4Ѿ��q�T� qG��q�xo�1.z��KhC*]�T��-l�S�2�j/T�-�ش�d,��%W���,,ZQ���z�[�����Z=��ed{����Ǿ��g�]c�j��Jo��fFFO]�;����u����^PM��3b�:�6�v���lw�y�Z�@�K�����И��*���Ohށ�O��])���-i�1#g�I�<}�E�Of���W��y���J%����6��U;&�:wf�l�m��559�/D���)"�"�,�*,�F��º�!��^�� �*����-�U[ųDl ����T���~f�k5�m�G8��D�{W���F���D`Z�A_-�9�z`f$8s�7��!	�n����`��A��$@Wh�|��Y�=_4)LG���
]�����T��φ����k��?0Ȋ��*3�.��Fw ���(�p�; �������{4�Q�������{�I�O����.r�X�f@�Ҕ�]x�{��y�4;�%������v�����K�Ԝ5�s��c���ױ��kY��[V��bF�*o#A<Ղ'tL�4����:�s�%����.�ϯ�>3��K�<����Zӟ�$jޢe�d�ꃃ�^ �(�ݹt���A[���BK��3�L�����z��;	���8QR���=���cg�`"�oR�m�.��=�z���z�DVu^V��!��>^��������s�=��xsiU|��z��J��atS��6cۻ�eI.q�v�'j`'�����Z;X7�t8�ʨ���@�*q֫�OBfP�*����6�4�N�yk���Q0p{?���0�v���bV�%B��Y��M�hK0 �UVЬ��s"ď�V��AG����&��A�NFq�f:T�,�k�O+�me S'C�ށ��3;�ͩ�%���_�ga%�允�L^�j�;FT͈S��nD��q5ǎf!����d����!O��l�%3�.�| �̖ �1��-s;w�������g&�����my�t�2�4w���_������'��JX���U�oA�b�K8�vfO��2ZZ�愵�#�l�xC̵A�/�]
}����G��Z"��OP�5��+Gh���ޅ\���Gb�.'�:�4�t���W�� `]�ݰG�K���C�3��#� qF톿'f.T\�˭����8s���{�C�E8^����!��0� |����f�Ni�D�.n�s��,�y�󇳳���7���6`d��mՀY�r�c���l������7�57�|����;W-b�ϥr�#q�`6��Lbi�Ԍ��⻼�QN�
~0�}�������t�ĩ���U���� 2�}x����8N�獏�1)RFЎ|.�AX�s����l�.JJ��0��0��/g��v���QӑsU���3IL䔫[hN��0�4����/�A,�*��vmg�$�f�["O;���<Az:w�c�E��L�]��h��2�O��],�`_�������Z�P�F-.#��7^� �j煉��ss*)�ϩ�ĄM�BHV]M@b
Įݾ1o0�r�/�~Eo�tz�@���Nt�]�&�pػ�S:������X�b�4�Px�3��ۭ��<;�*�IB�1�k�+t/��4�뀉�gbi,���|k(�T��X��I�;ϓj� nG*DqK/v�"6=����f����l���IN�ii��3�Cs�S�?�Р���y�e@�W���&�߶9���)�Ң�`��>ߦh�~�W'��:���*��Œ�,`>)S�ȉ�>�\���k��հ��>�n$�ќ��q�g�渑���]�zxu���q�#y�P<�;F�Vo�����j��^D��u�$r���8T�L	�(Z&����Cwd�SFM|d���Xه�=���E?R{eq^�΋I�雚�R�P������|���cK_^� ��P��*z[<��I�ɫb:�h��G� Zy�� �T!!�1���96��ɸ�r���S@j��l�D�6:��5�m"2N/�Z�-t뺳���
iK/젴xC��*M�bQ��A�$�_y��#WrF�Ne�|ܖ� S&�E�����
���H�h���������.kG@H>��
��_V^NE�T���U:kZ�\I��:�5�����e"_9�>Ê��꙾�+M0,֔���L�
�K�j���ġ
�yN%V�O��d �m.�nX������T5+��K�x��c��1G�e� r�����g0�c�5�����6�	���Z͠�>ϸT�9b�r�����Q"��ѭ�.WuE:}Q-�+��۾������v�U���׌��S���p�Z�O\�\�˧��5#OQ\A�}���H��iz,�\�5S1�@9�Ph��Ce8��Y�g�r3� V�V͊*��D����kh��0R�����qѱ��٧���l�F��ƌ�� q�vi�z!�5���-��܄i^��Hd�k�c��3-�^�u�!���;�Ȅ�D���5�����{^�*�(��t�{ǳ���{F�K�C8D�Q��{&r���%f��ܿoNp1����_9����xjFq��g8x3����[��k�{by��s��J^�f�w-/P> ސ��W�Lˈ1�~�	��bq�.�bA��B�P6�����X��(;a�	���R�}3�_��<��(�Pd��ݻ�1�m��D�J PE5�����.|{Ţu�'u��O�#'W+���V�<
}H�Z��A��D�-l�C�����R����<~�ҏB���
¤�Q���BT�s�k�v���Y�i
�|���qh�l_h�|Ѡ.�.��o桃��Qh(��Yb���,��N�:���K5Bj����)d���(�|Ө��ј�OM�������iB�����W�8o����J~u���UE>\
�S����>�y�#�JЪe	^.���.���o���L>�K���p��ͻ@�TA��z~$j�����{R�W.��w�`R��2�<N�Q����� u�Fd_��U��2g}^J�e�߄F-g=t i��mfZ{��d���dٵ�\�"��LN�۵�|m�N���:"���8�_��ye�\겖�I��#*��h��;>�e�6�T�QG�h|������I�Lof����2���a
ʒ����G˥+F\�I��
g��7���Υr�zsj��r�;��rF��kr ���@Nn�Ԉ�y��Y&d&��+���bT�̪ �P�����g�·�;�ߖ�~A�,$�k~�/DT�������t,Ya�F>�����+�"V����8A��hhQ���W����ݢ��E��4~�|�<3�+�0(�0B��x��{5�I�5�ϕ�'�C��J��)���i�c����x�	?��C(��9�`�\4��#�c�-W����/���f�k�_s��S�e�@�'�z�/I1fy����}]nNeS�~�[��'�#����\;�����t2a��Omr��*h�G!R��~�k�vRz��׹6��:P/���N[�y��G�ݳ0�������5af��I�u���j�m I����tvE�FK�j���"R�VI����&����xt��Դo�b�~�Ǯ�8D����|�<Y;�=��n*t!�Θr���	����uZ�g���|�P�[y��}F��b���B���9�A��g�C63��Q��c_᧋�n>��!OW]��&���I�Q�ph���P��C�F	�c\� ���`�B����"��8���8c�R@�l[�A���~������R�m�B�h��9�ֵ�%0�hV:·I���~e)f���e�:��X���i$�駚E�֭��N�4���A�y�I�+�Y��-�|5�"y���g��ڍB�e�;y�:���� &o?��Z�E<}�G�h�ܖ,�H�5c)���l����#IF݃'�S@q���Zq�0������V��p�h�Ǵf�����R�5�{[�M�^�����TE��l2N�i���1���F8�	S�Ҷ���d�P�Φ��3�<�"exP����}�� ���C�aW����~�}foо%Ծ�3y�k��k@��} L
O]��^M�=��C��^�j�R7�� �"�v����|(���G1����>d��h$E��0��u�c<0%V���I	NN�����tw��=��1o�1RW�O��Bk���	A�$��{l���U1h���]52��%U�I,�h8�MjR/E٪���@�4�(�i&Ƌ��QYce����)n�$aLB>L��5�pAQ�-
���*b�������q�����ue�!�\���η$��LE��#��Wiy��&���ό���'��\4Yͮؿv�.�r�	�`XȱI���8�#|�8n�e����"�,������������!�ޘ��n,}���5�����|z�-s�ΆP�"�D�M�Q�u���� �dSMO=����[u�Ti]H}����M�ں����+V��@��O+t���/�qڤ�L��Sz�r���ɇ ?���r�j<���@�I.�	��dEf�)`�d�v���A����?�x�(��6k�{p������#�E�����F�LrqRhgu��p�4����ۜc[���Zd����do�n��U0KŁ��&ԕ�3�YlGL�M�
�WK�0���X�nM���ٟ
��bI�73��Gr�h��^No�~`�V�E��-B�d���,s��}(����I�@��Vh��G�����N3?O.�\���ȳ& �g׸���E�m2� j�,o.`La*VS}���S���h|�H��^��꘼�2�C?�3�ԟ��0�OeS���*���: �P�!�&��)� �\2��^z��tc�̆O#�3|U��-t=�o=F^?��X�_}e"�`��}
JG��~sb6��{�g�%ZX��K��]{�?{�a���a�h��E�p#�ҬR�5K�75JZ��+[�ЄQJǅ�!~Xh1|������Qq-���+N^w�S�K�k��/Ѡ�F���@�m~u�˦��;ncB�	Z������{F+/`r&Γ��p��۔K�U��~3�Qz����Ɗ��*qB��{c<?EP�_��4Ŵ\"WPHe|=؅&�JZ�����i�k)���� �B+��u��~gD���k*m�G�u��.�[�A.,6k:C7�mD��A���1�(�?\|f\zƍ�=�!�wo����cN�8	��mkF���R�}��Z&�7k��p�ae�t�xv�1�NxC��ӽ��v�H⡖L�We�Z�*�y@�E1���mJ�S<�7���l��KǑ=	Q�/v��c����.��<�y�n"Ҽ�0��������H�T��#�#��Q��J�`��,䎀8��נ��Ϻ[9�R�Fn���M�Gᨑ�v�@Z��lA����� �����k��[�Ym]J���2���q������w/�bW�e6���X�1��f�݁� "���Tl��T��'t*[�^C 5Q^�;jn���.Э��'��?ͫ��m�H��
�:����c�V�f�\i�����h�p�$L^�3M�~vk;��'L�e>Y�n���9�<�`��y8�h��o|7�ݺaWt��0V�C��9�ߊ��Oy���ٞ��Ɏ�R��kL���S����� ��{_�b��9$���f@�σ�&�g+�Һ�ʜc��-�p�C�Mb]�IPU c
����#Z9:3'�0���I}&H��ۮ�Y5E�XQ�'�T�B��{��n�ut4(���k���!��9�t��KmQ�NF�M���h���ݼ�!��$<gE�5����S�I6�,���$Q�87����Z�7u���dM�w8��&���Ί@|���$�&��^w|��F�m\Qw6W_��㙻��K�
&� P��^F�//�h�� f�N �,U	&�=1}�P��R�_vP|QVh�L�㊱�s�W�鼷z��*��X��:���ut�O���E~(�U�9ܘ3�np*8��b��F��G��+-��>��p��=	�y�t�wN��}�Y��/�(�[�`����e���p��D*���pc��r����g����v%�+堏V_�G�z�|N���2(��fo�d��6�'뭕/sGc��%i�~��ى)2_�������MAaG�$'��rm	���R�l��ቯ���I�(M�7f/��I�0Ǽg��!�v�":)���c(>|���g��:�YV��6�rQ�Ƣ���uc|8�^sq��ϱ{����Z�͊�>�Vl���۱"�F�di1�i�Z��?,���	���/����M����{��Q|`���ƶ�0)�T�3��CO,�C	��wu2/��U���z�i�as�o�~��s�;Qmks���x"�=����5��c����J�0n�7Tx'�G�!�h�o�D�l��e)�r`�.��3.���JOr�j�U{4;�O��Z ��w,�Ջ����Χͱ!7�+c|, m��AR�� K���� ��$���w� �7�SL~&�X�LK2)g��0����|��!��(���c���|Q����Eu���.��5���hA����	��E�$;Sz� Clz��x�ٲ�-�t����7���jJr��0$��7��o�z�)0�yS�:JΆir\�,�����	�n�+�)fj�������rQH��´
R���>0��:& ��XRӯ��]��
���dOW����0<q2p��<��!&R+2�/�ļ�8-_�p�NWL/�y���M<�N����V�����.:�f�Z;�f��m≄�.�SX��x3�%�ȼ��e������z.���i��sE�0�Wo=�Vf�|a�wa�YU���i<�`{E��NU0��k�W�0|U��7�>l^8Ėj��1��X��Q3c�U&@
is�o�8At5G��Ix39c�P~XS���v�M�T�D�wC�h�#���vq���@+2	.=s��eh�NUH��J�em������[[�J>(�Y�Nm�-Ϩ����#�ʎ�z��J�_ٔp�h�< I�ǚ��}/�'�RM�9��� g �Q�}�k �Y��[P)�^(�A�QZ�
�Q4S�_�y
� X�J��ڟ,XE�%�g�rb�T�޻m# �NX&a�����Lm;�uvH93�Cn���\��u�9���*:P����8�I�ə4u�uYN��HV5�=���s��d��}��Ճ|6�4L9�Oh��J�B�K�\��M�7�W���xD��ؐ�6�"���G`e�iu�=r��r�3�?�S�&|3خݻ�v���n�5T���͂��V���%�5x5�-N[�����z_��6�e������{>}G���n:*��� �5vV	�)f �݄��II��H������m� ټ�E�/����(�s�1%6V(������hz�KQ�i��t�9�,]��[݉"�$��Y�l�z'Xh�?wⵯ�����mks�d+&�n��L1JYOt��oX�oM����`�!��*I؆B@','�\[�%���/#Nu%t�1���N�Sj|a��,�v�o ���ut�"�LN�z��%M'��^��ߓvB��+(;�z���8茩t���K�.�\��s��廚;�̀5�leJ# �Q:կ)mQ°� �F�*$�F�����HF��ߖ9\�;W�P���R�)�m�z�%L��V�D���O{�5+�Y{^\	�+c����G	�:si5ghC���z3��[���es��Gݯk�V�]���?�`���<+MJ��
y@5��t��hh,B�y�藆n@q��
�1��sl��i���L!������  ��w��b;�MM�R��p�SE��t�7+I�i���0��RQGc|��p�B���
�JNp�}X�)]����Bt���E�D��|��>&�����,K��GT�>��Es��� �$o�m�4�q��i��T��2��[C��F�8L@���%� z�di<n��DF���b�R���O����v0Xp��Tf��e�����3jЗ8v�@_0��:��Л���	k�)�?��qPd�Ai��@��s�XH��[���d>���Ҋ�H �@��s��}}��Ⱦ���g��
��� ?�ICl���6�֌�������0&@~����Ed�y`�1�n~J&G	�g�i�D���]B�Y&������O;�����Eup+n^阽w$����un���h�n�c2�����������D�>!��ؼ�2qd̻������n�a�u���>��y��	O�
�<���t.В��osU�<��挭fRSA��m8(�$��q
p[��Kd����T�������'ds�N
�	�lڡᖲz�>)�`8��c�?�_���s���d�M%�"�7�R˵Z�"[�}=�v)\>���;;M���@Pt���Ӡ��}�TP��k�mlO9�QְA�E3��q`����ڱ�G��e�D�I��~�Z��:BI���(�!!����IQ���r/
��(�@�iӔ��ujc�^�.^���Ճ�;����Wy�q@+����%O(r��a�5��_"AYx��pñ|QA����I���p��O�~��z$���Β)���s�LA5e4E�5\��ؒ\ԖI3�-뀵�Ӫ�x�)��_�چ�k��*!w�U�t�ml���s�~�rM+-Ktr���Q�_����'�1�Gdr�Y$�6�D` g+{�"bT���e��UX�P�?d��>��j����ZX��VV\QRkKz_��R,F)�el#��IB�H��vP��~MЁ� �ڮ�uE��#�f�w&MIYܹ,P�k^ڧ����v���p
dg �y��hW@�C`�x-��G�Od/�إ�j"����.dm��dd�s��
�$t~eyk���̄����R�	��rV�}��ȡ���C���6CS{>�0�Y;���r��_I� � Ƌv��흈?Z���bo1uhˤ���GEkm���*�:a�@]+�kaI�~�|�h~�(A�����QG���E�Ɠ�?� ��e��x!9��i~�7��Sz/A_���zY��4H�rvZ)
sn��EϕIw�l����Wi�2�F��U8s�V�MǨc[&�u�p���_�7��&)z�G�J�B(�SKt�L�@�����N{L�w`��,�7FN?��W�$K����R;�������l����W�Q��م���}�.��J�1�VlC�C U�+{yٽ ������̉�H���U�Hb�ҷ����*�d(tQ�P��D?��:'0��u�u�%�݇�.X�_�d�'x��m�(�&6)i�ήc�6Ч�>%�x5_�P�a��V�޹�:�zm���6QID�M�C�*�V%ɦ�b�b�W��=�{���U��PӋk\U�vkV,��n̨��HZ�o"hؚǫz�����8D*[��;��p��3�nݮa��k���p<mu]0#	ID�-wmDk����q;���s]u�GVq"�{`3�5�j��s�����"�bUV��;���b��X�x�V�˼�.2�/D'.[3֙N�0 �h���ṡDv���es�fLǰ�y�w­��*�?���+d���3ԃ�A�����R�}m@ΖHN�?�t�w��27�?
�lj÷�?.̪�4��!�i�>\�?II����<�0��g��;�L�����Њ�g>0��5���q.S������7XS�N>�$ ���]�{���h�g�i�g��P@Pܻΰ���F�
b�4�,\���W"K �������j��8�HYd~j��,���ɹb�.C�!N��:���R��m��w����w�d�T�8 _j�H��5�'���D�ꑧ(���6���I,FU�G7c��ܽ��Ƚ�Y!����ˡ�G��(�f�^��=E���P������&�Ç#��j���3SlH
����K/
C6FQ�x���8��i�u��/����Q\�߅Wԝ�2�+{�u����>�����+�k��$BX��2Rvf$q����8��x�?B�-d���3���Mk �2A��H�t�>�5T�!�V��{G��^ܳy	�V���i/��z���nv�L�|�ˑ�8�ءs�.�ǂȸ1�ɤx�9A)��s���xVG�$�~&�w�T4��U6#9pN��[��le-��'�@�yN�İ�����`^�D�I���$���A}�����Z�Fzĵ1��G2�f���H�#�D�x�;�ڕC0!��T�?}������g�	���ǯ�Ʈ��.ѷũc�q+��6v�Y.�U2^2T�o/�W$����k�&��4ҬmVڦ����}�b�IƉ�Ć��b5_XP@�\�~�qoR��_c�� iU�8�B��2ChI%�h�5�K\������Gլ���G�k@�ϰ�B�pR���8)2@�P�v �ս1�|�,Oʃ�[�4x�f4M*�Jq��q"vQ-�:E1syϿ-�����c�'���hkV]�� ����#b���XP����z���T[6�u�nCk���s^��6�MO3L�?j����K�x���,X�l^/�^�g!�$���7�f(6�H�\U��I�p(�~V��{�$��q�=�\�Q�/�7�d���I=A9�ϻ����9&���y�GW�kIز��o���di�	T�A�]���g�K��!���n���UkyQH����|��iLd$�����]�E����_U�K ����
��e�2�%S͘��d���Wt�[����;��r�X���N�`?��` Y�f������c�|�~u��?�W�u��c�~���[�3͘�~8ct+�$��;0z3N�H@l+���(����R��?v��Z`m�W����
Ǫj� �`C�b2��W�;!���|GT���iyK��zJ/��
��w>(��3_Z2�ԗJˌ?�/��a[�;�U�F�u�����9���(��:�7+�	rf�3�@Z!�� 7���
��[8�)���1僄ʴ6�N��6(�����U����3t�������e$�T��cLY���WO�(��{�/�&�����9��p�yHȰ��z�: X��p⮒�+c��س.tp�|�y���'� 7'��0מ�j�Imϋ�&|���+`Y��-U71:g>�x	f|��*��"�� !&7	o-r�c<�>���8Ed��o��F��)��C7tПGm,��*gy���-�oP�(W�X��X��J>���w�%]�j�OH,�V�>t��2&����cN�EL=�]�
>��D�*�rHbr�4��P�H�]��Q��0;<:����Sn8 ��֣O��B��n�Gl|z������A�)����d&� l����>r͡
i�x�k�x=A���H�5͹��qP��,�҂��Å
�	<��H���}�sz�H��^�St�;z_�57FB!04k���.�*�_�0v���Jp����?�pm�A�ϣt1�<p�n�p����1H�>���=~��f��|�C*�2�B�q\��)�석i\�˩4u�S���wx22R�z6�[�x�ig�8�'�z�z�A�
��@�DHHc�|�3���^�:�q �����"��\��E��O4@�{d�l�ۥ���y2���GY��F���0 ��cF?`v�R[�+�`�-���2���X�l���`�������y��	j&��$��q"~���l|��I�v��+Ӯ4'y~�x����"���#D[6�}���9-_&U]�[а5�j|�fH8a���4����i��{��H��y�M�Ya	�\���dKQ��n���d�{��,ޝ9XU����ŕUf�R?7=uC�/�eIn�
���z�!KT��8�͵�H��!'��$��;�<j�y�4�ļ��#��#��g��\%y�`��:��/C�ϰ�PT2�^��u���,t�ª���/QӚ�QbamZ-�I�_0'���߬f�{ �] �����:i8s�(��O5�9:ι���aK�pN��T=�<���@;�<n�s*bU�=�J{Lx�?�����J�h��hl{Y+, ��j��\���"G�<C|�0�<y�(�~�3
�xs|rm?psf
�W�9������?���o@D��U�g{q@�J��w���h�0���j�0u9
Cֹcuݤ�wyː� �����  t����:0�)1(�>��WH��?�w���-�+ߣ������%��X�Ȉ!�G��YR<���M����ӽ�K���G�	�cJ,wF�!��fY��8$Bb�S�gc
���@�롹W۷tՓnǵ�CԏY���8
P���LJh���?�&�ж���b�f�ꈝ��k�E~zI��[d������Y����s��r����}��̢�l�i���ߘ�w]���Z��R�,ZSJP��4�U渵ۆL2�[5r��(+���>�����	�z�y���j��Q5,XJ�H2���K��a�3��{�
�5@	(��������jAT�q�+6;�df�?�� ���q�bj��?���g�������'���ݥ�3���-'��y<����:�ӀVKo\�I�Љ��3�oKD>��M�۸��Ee�^�̂�1HU��E�]�Y��&"�ߧ-��d�BG�@UF��s��I#�P��^tg�X�_l��VJ��_��g�Kk��i�\�m	+I�%P��a����O�d�H�Er�]�%�C���X��o�Bq�����r�?���꺔�H?7����Ra5ֱ��%D�������_CϽ:+�����֒����+�AQb�r�P!��C��G�^��v���(��o��G����U&Oq9�h�#�k�?
&J�sb��K���hg<!�p�w�;�j~ ��� �)!ž��j~AB�W��q�,��V�~E�`��{&�=�zP+O�ɟ�;��ӭ2=�8���)bAEp��.y)c��n�sQ���q���'��������5}3�Z����ޯ� q=Ȇ`����0z���V�Il3���]��Pcj�q�L�B��D�҇m�(ա����F�J�u��Jv���
	w6T�6K�s�!��-2�'��k�2��ۋ		⊛wgKS�H8��x�pB�
u9	-�*�g�spM� �1T�W����8 �cC�T,]� _��A�nu�M���t��H=y*�f�_@��7Bs9G/��=��
F�MM�t�`>F�Kt�BD�����wJ%T�pZ��%ú�aQw�~��W�(��4)+�񣘕���%)�h��X;@p��##b���Q)�@�Z���3:��X��/*��~JU�a�Ĉ��*J!&@_͝p��$H@�Ad� �S*���5�eo�n'h�
iZQ���x,�غ�1:��q��a���4����p��2b��Lb�V=�N����<��xk$���2��/ίhZ�bk �G�!����KS{�T��MH'��n��G��H|�Ї���ӽҕk����zD�C�m���Q�v	��O3{@;��R�^�v����b�G�N �h�T ������]�d�����v� X�q.[�#�V؞��>C���>�9�Ӝ$�ڮ�'Wؗn=$�O>? ��c�6
�8ڙ>;ܕ�4zѝVI��n� �M�b����d�VC��en�v��wU�{�&��Q�F�c�ʗ{��B�	V�'�5���3�r��l�[�ćM�~��(ۤY�R��#kv������[�2� ��k
 ��';/Z j�3�Ͷ���� ru����oǽ-B�Sz=}IQa\+�ӌ-m}S.�����al�NO��u8����af�R�W{�#w�+���C��f+ ��2�Q���o�O�x�Co����l"_�u�2ĞS!���yA��ː�\"�CI��b9dC~N�=}?�(�}ō;|�9ۂ������)ΗE�7�Ax^I�������Q#w���r�H-z����I�5������D�*K���<hȪKh�l���ݔ���{��ZE���P�6���4&��[y�̪8"�	%o+O��E��z��>	��z� ���=��� V�߾���VV���/3�}��̮���w�$���qWxC-X*k��%봏����;��2��Б`e�C�z���\w�h�G3s��!g�'���#;���z���-ᶦ*Zx�,{9��s:�v���cܟyC�˹�	)j��d�k�"+��Y����H('3Pg<f�8�A���ȸ��󇃮�۠�m2EX׉aM��6 ���O�wӿZ�FX�Ӎ����[�ۆ;2�#ڧ�@/��^z�У��~x��  ז��+e�Hna!>�$�uM�Hc!�RSM�=�J����п�{�9��ۍBϠ�O���Q�>|�W�C'v��X�[���&��׸�⌸��a���	CLej�0}D4���V2�h���rV6��H�l���P5�ʖ�m�2�Հ��������p]I4VϩS�N�7&%�^���k+'��F�J'�i��|���^�����2�6�?��v�L���:Ļ�i�	��0w2�pҥ�M	���9���5�]���Nd�y��Xpz��@VzX�~/
�X��>F3�4�cǦ�&�,�ⱽ�c5��K���7t�16������u"��.-��%��l�h��]PG�.�{�m�?@!�o�|T|	��뷴7L�Y�8o�!��4)V�:�M��'�\N���4���c��F��������c��ޠW���~!��n3�6]AVُ�&NB/dH�U�==>ާ�
HxBc���Gg���;�J�ޝ6c�[�&�n����a���ۉQ�m��P���fM�Qԣ�ysO0�t�q퓮u�\�K���ˊN��kkq�*�R�����U�ȋY\�X���3�w�I@�&�o����C���uP6Eŧ�Y�>��_C����Q�8_����j�I&���Q��`l����q�h�O4����cjB�U���串H���<5X	�m�4�����on�ݱ��{<�5�t�]�n��}���U�|0���R)Q��d	@o��_�0���i���K����ԯ-�^>m�ABN�[��E�� S����/�� ��������ĵ�4�	����m'��� ��VM�KVKT'W?��X�l��L ����Dʫrp�0�CQm��>,�{[��W�_L���]SF2�!vHa��?X�8�c������W��|�h*Po�X"�ͼ��Pi���Or'{J�?���(:m���ϣ.����c���'Z�Cϩ�f/;�_�Tkz3EP�Ą�<��6{�I�T#��۴~���֌5�bXG��$���O4iѠF�8��($��H����M���n#NB�iFh�/��>:�%�H�JǛ� �ԅ^`	�@��@�U)�}S^��`jq�-����0 ��DQE�?l6,���% R��$�]�����4וR���@�ƽ�c?��Sȑ��$��ڳMe��;	S�a����Ό;E#��N�b�Kp�c��h�0�)�ř�l
`W6~eR�& �������Y��
6 &̶��F�I9�߯%W���*fqx �^@����*.�Qۀ$K2ꍭM���jG����_�Q5�@ w���ǂЃηTe����~�%�&0���έ1>���Ȱ?kB��%=q۔��*0�k#��K���l���ĵ-k*g�	���j�-4���Gr��?y%�|����X�~���,?�2�p:��a�K�v<��hU�`����X#T[zX��ҍ��
��{3_R~�	Iʹ����'z�I��/���L����tY] {���i�>AJ��zD�[���H��j�1[������x��c��j �'~�=oep�NAYVU�  ]|
�cL=�R�DH��vTh¤YO���g�Q��v�ǉl0��?,���'�&��nZ�`)%F���ę����C�p�}��[;n׶;��/�eP�����?~����`�Dt�,D?,Q"��7�2�ʎ���a���W0����l@�:B�� �h+=�H��)`�)�KR=*�cr��:�h�l.f6g�Ȥ�F����k�4dC���q<!�̷	���N��\����~�,t�a?q���&rSFH��;5P�
���>�Z�6�j��,Q c���J�	�c�|F�6Wz�C���`2;��6�I9Jz#a�F�v2c#�:L��\�+8�f?3���j~�}fɎV23�	0�c�-F���V����I�f�a��w��^
N�kC:r�=�i�݃��۳f���Qb�ݲ�Q�5n�KA���}ᖅ9�Wh���׬�H�9 ��m��˺�NN�����(�]���i�1I�kiA�<N}�2uX��q��/ d���OX'J�/��dk�4��tu/CI�R,�åY��fe41��Gk��=A��a������k����:�y��V���50�#�p���H�0*}ccB��ٿ�%��إ5߂��5��ӊՌF{��e�#A�+/V���W�X�=�kڏfC)�؝�J���	���y��4|��e���#8uN�.hb�U~�5�A�-�7d}�� jW��w��6T�ݞ2�pTO��c%|d'���U�p��~})�6���\�X������)-���v���U<yk����)=ϰUȷ�j����Igg��T�%j�V\4~Wz��2)~}�(��ڎȻL�||�ń�
��h�}����+�K�}��m���L�,d1�4;%8q�*�«Q||g����X�il.x.�H�n�U�I��xl�1���M�XRV�G�?xԡ�!k�e9�\9^+w���As�e���cRt�>���h����HSF"�K(Ծ_�#��da(
���U9�.�Q��\E���M2f5~Z���%�X���2��|�c#�RO��3���O.�V�F�/�+t��i�"���D�w��9�S���M蜷��v�ƫ���@� �%��#^�@����v�����+_X%_�Ff���USF��i�vg��8l����ރ[�=o�L�l���&7���m�!��E%B�Kk�OL�DD$YLQ��7��$�w=�f�d�2#h�r�S��,蒏:e^Ȧ�z	��1�x!��FX��~��}�Y�A@pc�Q8�l6��7&�Z����u+h�<����䖵�G�a�!���hB�tkԐ-C�'���;��~�9Rb�nгn�("Yp�)�9�-B.ʢ.���]R��;^����`��ۘ-Nq$E%�=c� 7�4���?xL@�̰[8�5�h��:�:С\>�Ȍpe��v�Ȣ����1��	�KW�<�] ���o�=wo�>h�!���:���<�ߕ���^Lq��.��T���`�ba6kǗ���n&�:��>$2ߔT�1ɾǟK��"y��g��u��,,�`�9P��<��wvIf�7����vmȯ&�@�MbaK*;�q^��׎���g0UZZ� ���� �C4���t�V��V�p�K�W&�`���Z	r"�s�N;S�D��`��t�[�3��G����3�P����D-?�S�ȴ�Z���d���*W��`;i��]�f���A��e&Ǆ��yd��V��K�Z�0r�����l��`�~Z �
J���%�y�MJ/\$u����V݊v���S�ϧ.���- �|�A4�`\V5{U�A|>�,�Ev�=.�ٛ��8#�1��1U:��_E{Q8�>f�q��v^���ҹwp���}���ۇ�t�킪�b�SAt�7���0�ŧ$����Ja|�v2KK��O��L�e���A���d����j������Y��:�s�~��s5X�j��P�fq�ݺ���7�<�!�w���e0뫬b���p�Z�"F퍧��m�C7[N��$w-	��)�T���*'X��G�5���$���'��Yo� �N�j�\�e�5K�7.Aޘw������-�	j_'ڒV��3R`�{ab�͉���N	<+���l��`�\�`�=ɭs>�ؤ,v\�ߦ�;I�
�[�B0>9�*8���f�U<��������;��q����!D���e���iș�3�B|��Gc���x����E%ųn����@��3|�o[!z�7�'zA偅
�ߗ�U���M�`�&�#��@<�B^��N������@��E�Y0mI�P����H��y��.�r����q�Uq�)�����tQ&l�"�S?����-�w��}bD�Ҙf���E�_ e��cV�#��6��̙���a'��C����;�+PP���9�ׇ��^��n��쾖���?v�dԟ"ӛmㄅCT���8N���
/ۯ��s�︡w�6�Uf�	�Dz	�9�D}0��뭀.W��5��q�<��'��U����f@����hD�)���~}'� �qC��� i3DlX	<L����,�'���K!�Ǿ�7V��]�*k���+����D,D��g�JB�n��-�m�$V��=% ��/�{i#K_=� ����gJ9[��=V�򕦯�#'d��1�$Y�"��<v;��D۪y���c�i�{�)Uf ��g�/��7q�p�	b�x���;[���W�!є3M��@��.��C��T�	t�I���e�A�%J��r���p(p^~_7�w�ۖ*�?;f�鄆bQ�3I����*8��`4b����P!d!~�g���̫y�̈́� �%G���,�n��(�L�7��"������I/�k�a��i��=�T���;I}
Һ��e���
';v�V�0��-��1rTX挋tЯ��in��7{����%�/U���i������r �g�.1�ZY�܎�V�f�|D��H����'�SP���U�2��J�|���K:T���ˋp5�w��'���$�vd2��tI����?܃���	�߹Sθ4����t�S�~C���G(Z���[�J���I����,�,.RYEw���R�+�\Ş����J��T`�K��<n�y���du�3�z-�#<�0�P�����d�<��s���+��:�$7���;���R+�v� ��K<8W(΃3�˲8l�z��M���V����bE�C ߻X�w��H«������'8��jӘ?�P(䢉�a�F���s�Ò뙜˿��՚�EN��l�'���?����=��f�u�!`g��8�D�X˽V�9�§��$#&o�!�=X|\ѳQ"P����l�t��'����/-�W����1�����wY77��?��r�f�N�^U뀞�����|aS�Σ�����wۺY���^lҷ�F�7��xh�����RL��y��ԝ��oʁ�:r*�n��$-P;��C��wM1^��IK�ˎ�Hnt�+���\��3�ȩ�=��b���ًמ�������[+z��w�¶EhJ��N���\�6y"�E�Z�1�d�2��@�"M�Wŗ����Uj5T^Qe��êт�K����ܽ☑���K~:�����-IwZ�.���py�^��A�Î�)1X����)�/1��b��bx�wU��$/� �S��I�=WT��9�)������gU��B�w���GC��^�9��lQ#X�MȏA�n�|4�5~m���Nf���o�A�n(�Q�,��,Gq�)��2��{���<��x�~�D��.�����X�+�g���ϹS���N�:�v4M�{�!��c>������?��ӽg���t8<z�0|�l �a���k8�z��Ta���������`L��F�Pt��|.�E؁z��Q�.��Z�i�5���D�6�����,f�}b$��^���'?\��1���(]{y/D�ճi3t��/Lˠ-W�GM��)�6�oK�jފ��25PU\9cV��'�t���Ʃʥ7�l�U�)jI��P@)���(A.Xm���"^�ⷒ��v�]EZ��_��C�oB���҅p�W�΂�D+��$�P�����������c-�뚽['x�P��|L��M�7T�mr��C�������ƺ�_Ue/^,����+���dǱR[�F+,�dG�Y�R�������R����I�0�F�FlG�+Sۉ�v|F�jS\i�X�3*�r�{�j�0hV]y:5��>F�JJW���6_�>c��Y>^� 0$w�Q�eF��^p(<]>c�����#�@�K�05iI;������$ 3 ��Kڑ��q����^��|쾩=������-�m4��~0؆X^S�@)�TR�M����6�@Q��r9�Y�M�vӾ��ۗ�������-(8�R�����@x��g#Vk[������"ZZ�Cy��e|����!fJ<T��e�[�/�Y�?�O���L��e5+�]��D�,&e�x5j0�xj���؝�Vi����߶�
�R~<^v��+�n#��w�3�f�&���A�z�����~b�\A?l�+>�o(v��<,� K�"%�H���o���X�(�
�v����8Q�7h������R�3r颭O��q�hk���Db���g�8�����-B��|e��lAO)5ÂD��.79��s��>"�Y쀔&��H�A�/M�C��U���p 
h-<}+�Y�n6�s�Wm3��/�+i��h:����'R���R�T*�����6��Mpw�bhÈ9�]w.^f�C�'\���.�V$ն��K9m�s�eX�0l��
Y�	ٜy2J��nA�l��š��Gh��N1��{��x�D4��8�P�;�? �˚'ݩ k�Td�7��{�}�<�,g^�h<���Cԍ�7��T8f��)�(����x3��z��2����~������;�.rj���V�g�*P#f����A�|�H�����}�+m�������%=�-ɺ���B���Y�72r��������%ｮu�5˩h����&�Y����+^/����C`\�s��/a��h6�V��W�u�)%rm숪7��d��ʐ8v�������[Z��y�l��'�`�o�Y&�|���9��i����7c�9R{��s-HPx��#���aq�Y	��z�k�X�HH��\�Y\b�Q��$)�K���~��0�"|.]{��kQ�_��r����K�� �v�f^Zl�H�7��;@������呖ew\1+]�.	]������IE����u�(������@��'�cf?���!�N�wֶ���$g*o�?h�� \;�ki���1X��J���h�p�k$�LZ=C&��P��p�쉸�-��ϖ�fCc�~s��~2�� *�G*�(?���s��מ*0j¡��,7�A=x��?�M��r�wL�ج��,��ҽ�谸K3\��ϵ��_�������˵�Z���OcK��Q"��洹]�+�^\�C� g���f�C=p[���R`�:���!�2%�w�qHˢȥཹD���� ��/]���&~�Yzf1E�MFw5��|3�2"7k��V��c\-󹏦���`��u��j�û�{F&�����5��r�wׯ\V��*�Q��ҽ�	1�S� �T�^b�I^�z�s��K�Bx�53����N���_	kL����'�׻���W0`�52�dUA��o�<���w���c1T�	��^A�f��]1'����5�����D�
k�Q���c�4ZFc���aQ��[�����"�f$Өu˒W��)8�����%Xk�jhE���IbN��O��zaܫ�Z)C�!���/�J�l}"�Az!�X���F�i�B흿��v�g�_�����\�Cϼ�K�w�Ր	���5��gJ�ա��¦3]�?73G>pAid����<��\�)��Z�z�Pe��ǿ�
i`��JJ�pn�[^x���/�KS>�ZL�K�%�Lg�4���.qM~ӎ4nI�y���Й�Ao˚p7���R�ja:�@��	2�&ɟ����7�1����+[�4��������'S��^�?�DdN��q	�nGk:�L���.q��P�O���l���TI����u��<�_�X�\	��؂/�����<�KG��լ�4iutH}}D�0���ˎ#�D	G��cf��� �>��/����t贀ȋ��Kj�Ἑ&���}��t���[����j�������F��'Qt̼'�@���Ttz�FЕ|�qDW��gX�` ���W���"�v ;�g(�5޽�.K�B���«DA`�)5=�s5���W]6k�ٸ�cGzޔO�/��y3iG�D#x��e�~���1�]tiIY��=�Fb�;Ƴ�Pn�Ԃ_���9�����K�X�]��F���r<��g2�LS2ji5�$��:���w�{p5zn/�i�߈�m=�Ҧ�t�_Y@XyIܧ� ���v�CU�f%�ZTtry{��&ˎ�W}��|o�囃�/�W�K�ˁl_�"�2�XÁ������;�Q����V�
=y����+��:�W�MK2G���b��sx���oT6��s�nw�DCvEΐ/���c��g�1�m����y���ĎS��T7J���ji7�lѺU��b��t�f�\*G�^��K `�t��j0��@�3h���ǟ"V_�(�������~/	�g���G��)��V�x�M��l�L��;v#�m��`�i���c9t2���"ͅk1��5fw�$�9/�B�ow��C����	L���p��8�h3�_��ƹh���Bd�uY̩
�F6f��埽w�!��r��O��۞?��,|���;8��T��'[K�>oB��kJK��T���6�����[ӾA�-فg כ +=e��V�/�*����[4�[�������X0���bL�ǋ�:]���cAe9���PO����X�^Wloc���B�TqU�#�K��D�w�� G�B�|������{s���l��.��.�����M�㾔�Bm��d���W�O����tO3t��r?x�r���-`6��U^��~�&�o��^_�+�L�Eyk#/�ą+`�d
i�3��!��6�%j�������5[�mHڑbHxB>z[ĉ�DS����%u�se���I&+���z,��l�ʣM���hrSī:�߸�$ۯ�'mŎ!��c��.Z���%�Q��.L�𿷣�&���u�8��l2-��S�NX�IU�[^��dK����uS��o���K}�p�ml��J�l疈��D�Rcp�W��4v�^��EX�Q�rZQIs�?�q�'<����a{�φ�$��~߃&�sH���9� n��F2;��e˄]�Тj��>c;u:�V,���a�ǝ����N�VӶ3�<nb����V�����nW�6.�����.�59T���dZ�
5���~JF� �4	cX����w��@��ϩ�/�'<{�~��q=��y�z��Q̗�u��m�o]�)GBX1�c��x�p�(�l�9K�l�	���5�8��H�E)d5���`>����S���o"��L{��,�Q;c[o�Y�] 89;�SH��Z�tAv�{��ֱ64�Ģ�^t�iӴ��I��\1�Zm*-<�`{�<���s����ʞ�f8�-H�����y^Ox;�Ф���R�R�v����sb��7�[�����+/�Ӭ3&H���P�9�qV��b�OX�2f���$)� �6��l_�P�����'��j7�K�K�<*F"�KY�lgj�㙫����`v>��9-�y5��9Ñ_�}E���B��7�9�� q�4��Q,��Vb�߬��z�>����-�I�Z;�>�q$�c��%����\�ԘB
��,2:g �n�m{���&J�6)j$���j��6��qd2�X�U���	�`Be�s�/����%���K��EkH3z�x��%�5m�sUD�s����~�	��ܷՉF�c�"�'�pXlT7� ����'Js��u��K�\�[y�J\�"aҥ�	b���6�1;��h�Y|e�����������z���pL���n&��y�	+a���������vU�^�20k�V�@?��[=	�Y)G����D!�����%f���֏J�/�58G��I4$R��~�Y�6��S�[K��+C0}5�����=Rӆ�G}�:���0I���qc|D���2�Gg"	����*$~H,nM;�Bx/�JXt��J�/���adyc�]���UZW�1�+�S<'��v|Z�i]�r.�_y��`w�T�"�XH�f���*��l¼�21�T12���:��'��+HTd>�>DS����q�c֤X���.�H·�zƽ��W����������'�i������7AlH'�}͂���Ҁ	"1P�����)�._�U�D�i���~���c�=[*����Y��P�h����jȧ2��x��<��'lPSu���xC��_:��$���v���*�>�_r�Ҏ���P����B�+E��� ��3cܱ;��/yEK���9��$��%��5b��K�M�0���6B�Jd�Q��є���b�*g��5{��xK��Ù��6�8�/o��v~�b�p%��XلI�1VD�^�,$l�_z�_R��b	h�ҕ^�ǁ�౗'�79��P���u�֍v�%g������o�s5_i�nkI�կ�; �A�G����ﹰtm�B�ƙ���E���j��o���hN�$���aw-�I$?L8�.�"���m�3}|,��ϣ���Ңp�r���t��n�/~�������tG�q��i�#��`��^_0SǏ�D��9�fQ�Py������>k2�-<�e�SثQ��!FK!�9�f�Q��*�aϢ�?Ŭ8��,���W��6sw�*��>R�z�Ӳ�v��wdA��h��'_�;�(&�1apwhbG_��D�W9��=q��>R�G�?���>�d�e��F�p�:9��Q0n�{��U���*�C�s�0�հ;��3�a�G��!gz���>�8cw|��)`�H@DG	�c��Gצ��adq�����K�v�c+��}BF�T����B��x��H�z�FH�71]6y"�� Ң�)��7�N�9@���� h&��gO��?IӥH����kmW��TzX�\����H�ߵEI���~�f�$���d�� ־{�ʇ-�2m������1�Mky�%(���<�������|�}�� ;W�ԥ�-��c]�e{�k��w&�
Q����Ѻrw)��v�B��q���Ic;pY�M�2j_�,e��WK�����FV��Ơ���5� G�:*{%�`#����ͣ33��0�6��*agA|�����Y���`m6X�feT�����b�&3�~���h]XJ;�6Z.cg�>�(�o�_V��ܽ�)b���B�4g���H�K��{P	�����Ƴ�dy��kw/�(iYe�3��ռ���;^�@K�-�5f���7�.�q6ت��)Y���[V��/��U�ؙ遉�����k�#ȒMrV��R�̍��Sn�G�Ǻ#���Qrr�{"��f�W�l�u��c5:�֛��&[6���]��^yx�#c���	��g��)���cX2<d��7T��H��dD�kLg��1����*�fx_]/�X7Zd�kr��A>	���?*�Lh���+�j��p�WA��/H�ϒ�����Ѿ�����w���?@xʄH��e]A/�t>��>��P,|*�5�"#�˧�Hw�a�Z�y+M�T���?�4`�9���;@�������ʓ�o���pYuFm`���a���*	�kBk�r���k��O�~���Wa~ŨY7�8��|��?Z�$1��4�	D6�7��&F�a��g�;^�
l���K����LR��e������gd^`k��M�<���0V�ob�}Ce��rk�&E���O!�lqZ'@R�p���_��\%�(ٵm����a�2� ߉b�̋>���d��<����t�R}҉r��cǝ��j�Y�U�����ѶY���v\ӕu�,l�w'���|����S+�t��DKK ���ȉ���7`z�FT��.lϝ�n�kf7���A
j��\o�� ܧ�E,,��
���C؛����l���KEaZ�M_�ƀ�R��D���l�r�o��͸��hC�A�ɍ�DF���ۿ��EVI���6�r?��FE<�}Z�:���.YA��CM-(&֐��m�zԵ���x���3��Ǩ&�!�(�;��Fbai }����$o)Ծ�J�L�A�7
�����C"��\����T���S�ة7c�mZ�=R�$�0�JU��V��&֥y/������>ݙ�����0� �B"�L;��������ϙ��k�G+��5�t7#!ۈ��K\�v��,��~�[��kN��:ʙk�#��eK5�~:0�?�OB^�DF�p�/��!�_q�τ,2�D4�}��%�I��ݙd}�O�=/��;hX"����>N�=�ħ�l�'='�
�TV���ZW2-��.�Zw���0��b��u�?�����Z��p5�� �i�=I5@��l��f
Ɵ�Z����A8�V�/"�[�F����](�'n��z^�/ �������d�����<Pq�MF�hi"�j<�;�Lp�1�*�Zn�T��]x[��뙞1��7�[m̌I�F��~���P��~�0Ϻ�bB3ć���*Gt�c-�le'V�H�0���g�2���Y���8��S��dȹr=u`�|�s����¨�w3dB�pl*��7��H����MaŦ��8|`��W�,&Z�:�?���b�n^u}��L_�ݙ�P�C�nݺx���@�[s�84��p҉�?iPܴF�6�%���t~�MQ*B^�� [��l�SX{��S�z������������ǝN���L��)<}�D��u�cID� ���M�:b,G���c�b��>�C�Sޅt��۸O`Y����P⠞��ո��Y�dƮg�e�����3
�$о*,!��'L�v&�A�r��B�60V����VN�ih�m�Q�P�����
U��Aeƹ�m[[��#�1��W5q�*�n�.a,��^������������a҂���T)h�`{����d#4c�)K=z�	G��⁪Sl�C����?��@D*6�b���h���&�rJ+�Ϸ��PE
|�ƨ,������3]O�9�VB?t��	��������	̏mх�k�1�E� �L�m9��7PKv��U��#��W����ʩ���æ���)Nnrq}��\��R�Y�'X���T���ܻ�-���Lm#-������q/H�Ǎ���zH%`p�a�˶��Tj��B����ðڋd�?�7��<��%p�*�܏|�+��4c�Est��˥��KR,jl�Ʋ��l?��XC��>�
�f4]u0N�Xk�d\��:��Ѕ�(���u����z	|ai[֒��M�Rq菧 �����%�ZA�s��zJV�łiG��X4s~-�>��YX�hy����1�'g���^zT�
ʀ�B�:2U���\�*��GvN��j%�J]���B[gbDv���,�?�a�a�3ȖK�zs�;��BjH0���u�Ml�?�^�LQZ�X���qB~���Ꮜwe�m�7���G�����F�8��m��O�8�����4�����^4KcH�e�o)L,�(���O���*�R�	�0����rCά�:o�	�te��/�������!i��!�q��R�|i��ڝ���%����`WV��]�����5\��t�A͉X�o����%��ez!����j~!��b��"l�)��1.�w��X���&#�����k�3�̒w_�&��(��7�/{���E���������>�qu�i��O+H���B�r��&��P&>��R+MR7�l
�z�&��� ?��|������ �Z-��с?��&q��Α�,�-�85`- �en�\���\ξb$=�S�Ԫ���w�}Kzj45(Г!T�+t�U/Rc��WGO����4�<��C�y��S�z�m�=AJY
����_!��8�6�i�����[�N����C6D"0xpᣯp��(Kym��v(�>nkmd�P���i��U�}���J"n�u�hL�~p\�-`:a-��f#e��!'IkZd��1�4���d�˨�?�`
�T��0Q�\��������]A�n��7u���S��Q7��߁F
{�O<���%�xe̶���v�'\�t��d�Jea- ML'�ho�jA�߅T�\4Psxn^I���g܈��f��[άS��dh�B�j�l����x�9/��B(��]���g۳�o�L�.�|�?y�oV�ũ��u�.�7u�!�Q����w����q�{F�>9A�~|Vf�A���u�z�Lw�������&l���Ӥ%�2k�vF�Ż!l��i�7��t���RH�v2��w�Y«��Q�( ���:�-_<`��>T�c�@�u���BGh�[S�����uyÔK��i˙_F���r�U��2�����4���̬� 7��$ч���*ߚ��<�7����E�fQ-kt�M����=�|Y�^)��ؠ�1��&`� }�5C
�nK�v��*ƞAj�ͤ�B�\�Q�����"d��T�8/U`q�ɟ �1�L��(�5��:, �k��A�cI�l��p�L��x���]Ġ+�Љ
��Y��v{T����D5��by|�U���ӣ���;�o�����u�����3=+���N�&���v�8�����Nee�N�>|-['D��^�>�B����Ȼ�Vm�.�ꅶ��/KL�����`g���敿*]���NL��4=���lzI���9�e��:�e�dd6~t��@������/�p��p=�*��|�!�~��m�W�Y>��
�=�=�?�OU$B3�.l��B�?��ݖI��}.�Z�ƌ)�/tX�7�A�p�����	�ld���^��ɝ	���&0�쭟��ht�FJߎ��}O�������|2�|�rHM���Z��f�1K��Hqp�k�	3Z6cK�|�@ǭ�*v�noW� ����A����_��m��NJ�`��%���V��Q�Al���W �F�=�u���EPIqG�r��
D�ߟ���芻�����+tz�H����m�cG��J�4oT��`���X��Ù׹��GL�$u��m�[eln�	��Ȼ�=9�{v�U[G���#-��T�2�|'��S ve=E�bq�tY>���s�;FS�Y/ڙS��ɩ��}*`K�4�Ql��r��U��\*�������]f"HSo��f�J�_2?`]���l���/aQ� �k4�h�w���8٭9�ˍx��G���1��k�2C�'��5Pp�.az3<�^��HҦ���kat��������yy(Y�	tS�����6��a�h\������7l�s �"�A�R�Us�9"�u��Qm�jaԶ����H��S.��aB���3�U�ǕT�� <4F���(K�/��F�sk���[�2��b�*P�T���!O��]?ָ�<U��!Z�`~9����;)������#Y�ߥ��Jbߠ���yd�0���_<���� ��� 
E� ��0[���p09Τ�Iа�<��{�L��V�Si�J3�s����^�*2Ma"9x,���s){��p+R/�i��V𥖾�'M���z���}��i�E��z����5���>YG�
��a��KR�m1~� nk��r�q';������h��m�x�a��B�/�i�����PJp�B9�Y70N��b��g�G�F�Y���c_Ea���-n�[�����t���I;�V������j�w��PT]n!�r�����Z4	�Fw�|�$[Z�(+1p���)a�22�B�č���D}Z�l<{flݭ"�&>0D�\l'�Ʉ�y� �f�R,6Q}��S3/�.�=eqw��ҌLrT��e�O������ �5Y����?���骵�ڢ������]vrS��N#�2��8_� �*��LIQ�ϴ�y�a���ݑ}�#����؆�t1��j�Nv�SE��Yv�?Zg&o�>0�w%�ml[E�A��X�A�*��-�]jo��C���m��2��T�q��2�J�T�� ���ƀg��J��
��|�� ��' "���#'>gkV�'�	�z��,?J���7Q6I��/L���i���_��6�3Glo|�
xCLB�զ4�:Cɓ"q;Y�	��7z�oŁۤX5���)�7Y% �d��B=
�4xĝ�ʣ�B�{m0����맮)KuZ[mJG�4p�۳�s~�1OJ�:�4�G��(�D	�jkL���<��@�^*�]��
Q]j�0�n��>BAS����F3�U��R=ѩ/:�zS��������f����m�h�{Ƴ*�Q�:����t+�x���=10�I����X<�f���d���ׇ�1xҷ�S5+�Mpf��rH]�GeŚS�gUZ������ɕz���~(�T@dԭ
��jZ"BØN��S���^w*ǌR>e�$�o�Y�8���'�}��Y5�#C����u�Fc��IuH�'fha����/&6���?J� ^�[e�L���ǟ��p���ؑ;uL~X�S8f�XIĊ�HR���l����!�Nt��c�FǂW>�*� ���^�wΥ<���o���"���}���q�'�z�J�n���Ҽ�Z]����Sa_�pT�,`�b+�"��ss�A�!ͫƒ�?��E��{���F!#�o�=�$2��I�=�Q=A)�3Z,H6��˰W��srޘܰ�PP,pXi�����0�ZS���s3<B�5�(�rr* �����}V-ۘ�od���E%�U�D���*�f�����tn$�i����Ȳ���s~�>)ug>P=�ȸ�Z�s���:d����[���_~v���+2S�w(�H<@��↊	(�L�ɖx�<G�I�ng������4�쇹�;x5'&����Gw%q�P����`����uU�DִR������j����ж.��6V�&^��kf5��e�r��M���v��x���;Nw.��4pa$�����ZO��U-�:�1��n��_'ztL)�t��z��g!MQt����w"�8�������0*|����v�u� '�����$�0��o��ox{ݶ�4p��|���IH9���i/�L�"'E򫴏�����������hjT2�2K5�Ԍڠ�[�e0��3	o�He�p�F�Ee��
�B�:آe��5��z�v�ܐ����=U�I�G!��T�n����g���B6F��eöu�eL�\��K�03˛)$d�Gr����S81�r$zfo��xw^߸�'�-��ݔx�v�g�~m��@�5G��ȂK,lD��S������K>X�D�hZQJ[��a�"��H�b��D��~����m�ʈ4����C��򾲛;5?���q���z_����F�Ӻ����I��v�/����,Ϊ�ES�=�q<X'�!��l���#��%t.[�C/���E�3�X�=:2��]'��"�ŷ�jh]p���_k��wU����#����O�~h@Lӏ��������u��s+��B��o_-��P�'�7,{C{M)��|��ϝv���^� ?����A+wE�[S�h��}	��2!M����*|��=$*H=GV��v���t������ʑ�[߇��~th�֐W�� �q�PR�U{�%c�@��Q~���aH�!Z'E��f�aJL¡�v������[%q�a
��<�EҨ^P�Y�b ����?�N͵	��ξ�*[�kPUZ�,��_��܏��?�k���HSx�E�"�a�!iV4c4��-Wy ^���S��0��;�.Tס�%��+�p��Y�T���v�|�§��#�v�c��7�?�6��2�J�1AU^b�e�_���c�Ya*��q@��P^G�Soo��!�劃̸�^Yݯw�fB���҅5�TG��2�t��.�̿Q���eϬl0��U&�KT�{2g�������g3�rw�8���_0ˆ��~�1ձx,��5���tjs{a���T���s���H��Ֆ�K d�n8%B��=Ż�^N��g���O�M]�
' )e�-��%n$�"�wMs ��C��+���U����}����P̪�G��@����jZ�(%x`��GM,���<��E���x�R�c���"L`�8���4g\x���˃����:���(��������?̮�������7�Q|Nݒ��Fi���r��#�ld�����&���k��qA�+�T�qoR����^�� 3�.#ެ�ٹ���zP���.�7�i9-[2�(��K}]S����I�0l�I]Y�"h����ד(~�����۠ɦ�`���qi-���¼`�\Y5�3[�X�11<t��t�*�RA{��,b'^:�B!I��Ģp-l�`�w�ì[f�Zao����>�ԁ�G�/VkT��-}���f9[�JQ3��7��z���PP�-"�u�}v���f˖S��q�"���f.{�tA���bt���=���������)��^��k���*���1Q�3;��$�:���D���L�8AL;y
����w�D�L ���z�;$'" ��(���a�=��>��M�d���-h�Fp�!~^��;�)�����c��PT�߳�e,+d!��--��:3���d�:��2��g���T&;.���f�s�<��&�O������A�+�����93Yv�R���I�M�j�e��=WS�K#�ٌ�����3�w�����|�4���q�fSPV&5 b8o�ǰuSh��J��d��AVy�t�����́*PIϞ�l�����W{��x��W��͟F�6�+A��H�Qh�?�8�ہT�B�;{GX�3<҄��18�(qR5oB9�P����jm��PX��H����K�R3(�vŜ�-�4����)1zmvNB��y�q�H[q�/�h�8Ms����ڒ*r�i�����y��N��#�i��1���� S�j@L���y�"�y�V��4�X��ϼ��A1�3g"menԶwo������"��=�탨v\v�<`w�-�!�ʈ%�e�-۩%���Ŷݵ5��sH�S����g��@f��I��������+�a���ꗪ�"�\��%�]�ɂ#U���Z�<z���5Ծ����~D�.��:��o 
AX���2�T*I��k��l옖�_�YZ�w h�3�u�o�����i�����;+��l  ���g�D�,���C	�ϣ�.���#�w�9�����q�{�w��{d9��2
H�[� |u������g��zA3mh����ԋ.�7�� R��s������s��B0U�6�c.09��Q9��n�Y��Έ��5��8�r:����0(�E5��fcj��@�*���<[Gw�����-E��dt��d�)T1�1�]+@���f&a:�>��x�=��2\,~���l���5Y��t�b�pu4+����-�^�׫&�>ݍX6a��2�%l��M�qKЬ���@�r��-��l~*!��Y�.�a)���密�{)M�L����]��A��';���b����' �ҔZ])1�4�=9�VA���9H�8FRk<]��x��ݷ�������|����J����̈́s�&�4M��_��(�/��RV���M~�I}J\"��%�M��"K��;Ye�h[|�ϒ�K��ISȩ${n���~�yǮ3'�l.���Q���^Z���:3�� Ƙjœ��q7��DcX(���s��Db�o��iE������f	lyŰq)yp�G�'r����F�	ǝ	�~l��4Z�$'�H+ U�} X�O��ψ"�	G���� ���*����_{��`l��
,�0���Ŝ��|�eߍg~�aT3�1�,��/��&kj<��OW���9��6��J�a�v�I�X�����ݱ�=-�Q�dX�(�/+@�&�dCz�p�h/��%=tӿ��fr�K.���O���h�~L.��	ߴ,5|u���\�4�)*��[���[݄�������*�'B�Y�7M��R��ǅy33�Տ-��j��H����<�XϷ�]�5�H��Zd$��}�Q��E��־ښl���̥�b��=4�N�1�)�u��y�EeWUPB�?�,�0x~��8����j���)\i�
igB_�+�!�g�����5�e�iSO�a����f�ۉj2�n?�Qx�Qi��-���;�E�އ��+$Gv˓�4�1xQ�0M�tو�Y`o=HH�1��/ò�O��94W��4�X&%�x�$V�M��p�}�����	���@.��Yo����ŉ郔� ��V�}��G!B��������P��͊z��o䢁���Y�`d�ۜj�i��a~����p��=��s�_	0���_�u[.�|<��>twЗ�E�w��:z�g(j����1X�nQ�I�����@!�����6��gF���߂|VX�qn�g���`��A�4W����ݞ.C�d����MF4]��0C�e��z�}��®�l��N)�m1~���Bu�&NR�w��6��j>�H��+;��몣�5���l"
W���1˩t����1�u��Kq���V�.O��0��B���v�33aq��#��F�=f�����'�P��~tq�6L�1B��"C#���M�Y;$q�5�Q�X����<F潥A��R^g���h<9�p�;�_��~G�0W�H��W�-f�B�nKÁ���]��j��ަC�Q�G��#-Vk �D~^�)(_ry����{���e��B��
Ց���V��4��cuW������(оys+�����$�F�*z=n(y����yp�����LBM�r�N���U ��%�֜nEF�(ݧ8�6���@j!$T��p1��[�:��W{�����@��Uy�Ě|W�YNО��=�&6Ɯ��x��aЕ�p��k��~�LY+��o�;�˄�E.��Ȳ�qWVZ�J9���š�Am������Q(b
`�����D�m$J��ad��&Rn���Qp@+��I��^�����LA��琩�"q0�Ň���l�F��[A���I�V��^uˣ��6Q u�e���pi�%��M?g�/g���K4\� �Y����?[������u��{S���4Z(��͇y�	DЏvi4��e�qBfEG)[�g[��a��X����T������!�3�3��eإX<��z�Y�[o��U�ì����*8�Υ��O c�e��v?H���:Q�TQ-�����rM���Y*v:��Np��cR�+Zh5V�`��#�ss���p���ĝΟw"�%(�,UQ�[�L`�����m�y��G�A~��P���|2ѽ<,k�7��xO'�H�P���$�G�Y��	B?��0yї��XBI� ���z�����F����?j�҅�Cm����?%�^P�؀����0+�	��`t����U�|����}�;�����5��/n-&<Dp*?�D�=˃���Gj>�^��/�+75�H���0�DN��l*v+W_���v���K9{�>*\V�Ж�<u}^W�),�U��H'��)�aL����
�1<<����K7����I��O��� n���o�>��m8�e�isVh�`�	����y	��@c-���M�X8���cv��H[ٮe��9:k�N"�$��.@X�j0�|�Tοmg�����唤�K�l
�BT�g�Щ�7yt̚���|��'�'���أ�W&��D�����7��l��u0xT��u����C�T�#�lZy�T����G��{�Y����M�.kFi]�d7B˯������*��jxĜ��)$��@i��ҫO2WbC/��ov��i�Ц��l?)˽��BM���(d�v^�~h���T}S��s�	����u��t��Gx� з^�z:�����#���ڗM"^.:� H�ɤ7�ł����YΫW���Z�F�@�>��Ugh� c���9甴���՘��v�<UYR�А>L��ޞ�,�f�Ӏ�m�$6�_���N��C�q���kd�[}"�#L �?P^���\z�`��{�p��6MU��dX���'�)3����mPbS�5�@���h������p�,���LK��<���"�O.b�<=Z�3�~xl��l2�/�P���V�$�m| � �$U2wj�i�����2}25�����i�7A���
�q'������Y_�w��p�gt,�����*��*SO�_"m�@�}�����p�"8F_ BC��KA&G(���I�Db�T�D%�b���f�k�DY��������_�LW�uK�7�-.q?�KN�tși�3���K{_�]2���
���k<���t���Յ�1,�N3������q�U����-����`'�$7��J�\���3�E@K�S!�[�%&	Tı,��Eϻ��X�FA�i�V��%��~��%�Zo�8���l�@��
q�)�R30�>�h��[�?�o����LZ�tIզv�ˑRD!,��ٺ�-fzwE����+ ������H��T���L��ȶ ^�s`�T�����kȃ��im�x�B�d���Rٰt�W�yװQ�l�Ee��"q��N�L)�đD2�间o~�#�"��Z��S�K��v�[}���x�3�Y�kbA�6�$-�u� ����r;p�6t�����K�8�$Y���; ��di�g]����ޫ��W�>�|���?!��>%��5���-^<�9�iyf�b��i�3��r���(�t����(�C�M��G�~{-i/21�Xl��yO$�k�r\5���At�	���B���E��KR��)
��}�&��$*"��l��.������F����>2c�Lz��%z���2"��ٸo1ؼ�Aa��ѫ�)��n�8�_���j��O	���V˚*o�1��-=�j��Q�L47[ĺ{bu��&EE��V�5��J�n��|�{V�Y��i>e��ݴ����#i�A�C�0��9����\TP{Z�Ot�Z�n��V��@2���2St� ���v��N�J���.�y6?��K�=s��d��V�t��3�!�wPjqPDV�����r�;O�G��H�ݶ��7�ta��0�3x�ZOe���� zFMk�� }��B��2�hb(J t�I ���X�'q'��t̴��߬�ޘ�����<	�2U/��Ԕ�r
�:>i-��N�A��h�A��x̙�
P9�bkK:
T�/积�����B�F\�J�VG��cD�C���M��j	q��c�w��f��E��a�ƖY��VM[��?1��(�L�ۇ>VL�
b�pt=����d�n�"%p��;�R��ǜF�7��<;��}��>�ƚ�e��Y5R�ǵ�=�;�v�*��X(��;����K������ �l� �VQ��8�&�V�Z��L� �y� ���A���fa��,���E������D�2�gAu��b�h�S�\ӳ����Qd(��]�i۩����A
d���`x�E������>u=˓|��t!mQ�l���\]sz��p�vvǢ��w%�W�S���`M�V�vc�����(}o�ǎA�qV� �׃�ͩ�}ch%Z��t5-��]�Z-�Z���A5Hcc��~�����t1�*B]Xs��$�$2$Q�e������^���h;&���X��9[mWؙ����
+ɵ���ʀx��.�WE�g��̸�B��v���l������E,��A�p}Z��!G�M����� �r��vy���p[&e�/�8#W�;$/��YL���Y?MqZ��l��'(6��]�H������^5e��~����A�?.v�R�_�%���}�nϟ<����:>0����坝����y�F�]��3f~$f_���aQ6����G�_�0?	�BSJ(p����( |l V,7�����[<z
D�?��$,��}�#h������=Z�Ad�Z���D�~|��m7~��G�h ��� ��]�鍗x`?rҌ�P��Ԟ{��n����>�|�+!ߵ�����{��h�p8N��E�-oXM(Ar� �/%TVs�4��%Y�r���s��b��KL?Ý�B@�$�\L09���Dv��	d�&E|�"��	��6�푛uyGvsz�h�q>Q��O���hH}�I�o�W�W)�a��خD)�g����8��B���̜q�t/g=ǻ��&/I�P>��l�(!_j�Y��:�/}�yZ��4C[�_>�	�7n�*WM	7��ʖR��_
�>u+�e���=����w��ԩ�T�\��7S���� �+�22.g�޽��Q8��
�m�Y�K�i��e�X����@�;�|���̢�p�};��j��X/+ݒ�u��ݿ)3��hӍ�;�'?�ry�X�eX!$y��/���j?�>g�5�9��۶�0|/�Z�!��a�K������!l��Gf_��9+q�"R�:aa̟�un�4?J��O�"�/E6(�����s8��o�����I���� ���Y���Gu/��D͍=�w/�&v8[h�.��o����xÙ��a��v�H�x��5vtŖzbA�k�P�D����c���/��	�N>�+!F����l����`[M�X( (��4�r�|�����қ��~�~�^�{����'txFYWVIA��	DZ�:U�_b`�  x]c^��$��8�ҙ�&&|��/?G�"F|���p��A��Lß������0WmL޶��Vn��r��vWG�Y6W��������PC�%C��,^1s"�0C��
���	s�AF�M�Tb���"��d� n��êhpߟU}��]aꄍ�K�F�*$&[&�,ܣ�70>���j�&���5�\�roa�yE���K�E@u��+<�Tj�K��Ĵ��M�ﰧrc���JUp�("�?<X*i=wy#5�5�c�ŌN;8Of��9��|�/-$���ʁ�Z��O�ه�ߡE��o���{2����������.b	ɭ����{�J*[��E.q�p@����&�
�e?䈢��cP�FvpP�r��
%�9���N[�PQ B�`V��/Ne��(��>	��)bg���0�l�N���#��5U�J�q��3�fH����epi��a3q��<���0�~Ѻ�U��C����4�����0�gœ���aYa��+��	� gS-d_��!�'��}r��:kTv��o��ݹ2\6�@?�\/9����rJ�<t�i�N����ݯ�
�z�)�.̺��e���hϸ�%'M���Yj��~��1��k6�UONL�;��zR����oNi�L>���/]����k�ЋG�ȶ��c��� �}: ��
�TZ������;Ю?�ku�Um����0jM�s��R>LD-GG"��������и��K8��M�z\eM���V���8bM��l����bʖQ7Z퀜����S���sU�;�r��%;
l�G_�@���_�92@��_n;|q�K�֛���^�����C�?�&fR%/�`�tq��P��G�i���BP�
��#�� kd7� �e�לΜV%�π�Hrϋ��aH��|�x(r�$�
�[��������np/�a�2I̎�W�z�[�R��EҚ?�
I�;V�ɭG�*%Z���3;_�e�Q����N��$5
M������������Q�dĳ���A��Q�Z�n�9�O��r�pؑ�p8FH=�$:Q6�!(R��SFxe܊܉��/z5#���ɠ�۪��Jm�^0�����84q9}b�^G �=�ZG������9;���W���z�K���#��C�8g:r^8b�������['	�$]oa�T���7��S�>���`�^t$Wjm���:1r�C�V[o�9n7׎�Q>����?}��Z?ts�0ʓ������P��O'͑�*�����Z0�B�w�,��{D�`|鑴e�j��P�D!���YϾ1W��_��Ff��7���C��h霯9/���j�r�
��{&����|=�e��D��zI�'�pʇ�$Qu��ӌ�f�JH	����k�Ǌ� �R���aDC��e����k��D�ޞm_�v�5�~���T��v�<�s�Q=�|�ݺ���h���Vb������BZQؗ�_�;�e7��v�tj$+7*��z���ɓ�� �ň��!�r�?��h��GjA���>jmq`�uLm��1���� ��Ư*#�@��]��1kq+��O��	����k�0��ZqA�ґ�l�c�Ǽ�t�$B��H3�e��836���j�Q�oޞ
(@����?�6R�.�0�R�U[�� �]5 �#f0����(�Z�v�t�9w�9����b�4䰁&Z�;��Z&�`����(Bhu{�4���t'�)�B�l�z�uFA�7�Xk :�3r�Lʌ�r�D6IC~�V+/�N���/)a����JP�z���̠�h�&���=nW	J
�ю`d>�c��x�bo��E���tw (��ų{���懐61�;W�d/���K]��m�������:�����Rj;�0 �M}m��v�X�kǸ�alY��P��1:M����
pK�7z#f�v��4��b�N.��Y�sw?e��xψ&)|Ti�b�����_�Y(7��Y��snwv�k��!\����J�<|�-�Q���u��)ĪSfD�Tn��əY�g��뾌�	�����,v�W�t|�p��-ϬL�R��*��od�B�p�����%�-Т����=�_aQ����X��u�F�i����h��N ���}F���,�}�Vb�؟�C��7������Qf%�MW$��T"%�2m�����ø�c�\
崐�Dމ��?O�p_%���)�a�훒K:�gB�&1
�s��(�5�y�i�k���g�f�!F��J����٩�����X�S��c#�����[9��踢�c&�NC� x(K���ZL=�����r���9��<n�N�>�!��x���C���[ 龲��e����tl�7ٛ*�	3�!�+6�[Qc.��4�cB�/d��1��F2c7w1���i5uk2&<{I��f��#�9�s#2��^��`�H�G�����F��b6��2��eث��6J��H� .)'�^8n,O=�y[����|/��Wf����f��br�LZ�\qP��|�"��乪:;ճ�NE ŗ��"��g�o�������v���VK�M�3>�ʍ*v�b�kJ �Ś4�W<����V�((��@�]V!_ig,bZh���l =��)n�O	���[t����iFU��㌺�	"�(�Fŧ���zqmq���Nm`3Xx�DD�Ĩ �UeD������wSD.��(4�A��\�Ґuw2���s�`?�=�Z� �>?�Q��2;Pp�����yч2B#�"�>���,*m�M���Q+9���.z��\͟���5m��.��|�P0��o��I�r��G�䨹5���a5^���c'2}`�J٬Q��k��?��d�D,bm�By�<�ӣ���L_�_eٜƿ��u���$Ƨ����>hdQ����VxD�f/#u��q�����dblEq+��1�UO�qfH̢�/�	"y�c@����3��$��z���8����G�k��+��Zy�����nb+u52F�Wc1�V(����1X�~Wf@d�N�%��C&R�q�p\&y�_ot�	}�%>밈���U�@i��b�ϣ+��B����
Q�'�<K��H�����t}�bpn,�-��x0;K�쏸�x�i�O�O寂�XN���+V���ɝ
Za��(���<nԪ6rՇ�z
[��x��s���d�o�=-��hKn0��
�3.��!a�L��msN�Ó��puJ���"�'��!&��
�&����#�]eU�&�����?��N��P�=���~��`Yp����nP)~���H�����^��m׫�
3e��0�3?0V�1���6̓�͊�{-��i9K���3�]�U�ГX�Wҙ�y?üK���J�)5��ٰ@�1-{�Pq!���w�A�"�R5cҟX�P��grC�&(n_�V�6�r9{&Y��YG216�(�T����o��|/�s ��{.>����Zi�\7A�4<���X*���6k��ן��(�=�{�w/֦w�݋��6�L!�~bp�g��WF�(��vNG�I�s�H�?��	$���O�|ƽԳ_�p� KS����'����z��wHO�[�������NN,A���x��O�J��y�@��t�#�v�O��I�&_P��rpd�S����@T�<PY9��\�F��.+Ot�J��C~?4��^
Q �E�&���^��ȶ?,_`�=@�M��}�$���ʂV�@��sě�J�?#�9�"+�2=^Md��q9��^'����U���{s�S���&������˥4jy"�����Q%��_}�y� ��|���z����$�)����t�a��k��	l��+ej���]�^=~���X�TF��vgn$�4w�8�%vg��y�,>vZgO>���_�G@��9b��.�?\߅�4�'c�Q��Y%m�{�h��O���&���&[]Ük���9Qz؍I_%- ˌ��8ɑ�֙��F��$�x�|��*M=	��$�m�Tb��`�تg��A�}�,*�,�w-m������ZM�<�G>�����̬�'	���ˋFBq���o��~(�ER�R� d�W
*�p� /��}?�F֓N�.�A�a ���#E�ۚ�:���r�7}���9+��%�o 3װnE��Q��kd�!0҇�+���,�_�*|��8�\kh�31�]��/��s7"��{r�qi�ذ7_��������vo�fT�%E�?߿0J�X$���Zǎ/Gl�'�w�8/j�q�7�6�UP]5���堋+��b�&�&��̅����%'���$�<� ����BDP�����[�X��'��K$�r��
; c�Xs6�e�>�/����˿)i�Z�v��~�r��~�R�@aW���Td5y��ٛ�s#�d�,�0�I�}?�i��[���<��΁+�QC�Z��UDܝ��a��*j�9A��$�,�b$��p��2ps��a�?P�;u1z�
s����㰐�|��}�nZ|K��'g�Ǡ�:��ơ���F�^n�k��w��Ѝ3dw�ƞg��s��Ⱥ�ϓ����dN,}f%�Ч2�{�}�0;�<�1`(%�M��mkͱk��A}?�����Ƙv��"l�NJ��XV	�E���$:������/��H�85h��G�~�XYK(P�@DӞqM��՚
�nAhc�Ô����p�c��kP��fh+j�P�,�����Z��a�=�����k%ܩAE��i�}RE�S0�U��i^�?1�џ�^HP��#�9���H�;�W���;������΅vz�Q��Q.�h�V��\"ke��	H��;d�I�x����P�';ɪ
)@�� 3О������n"W# ����?�ǒA�-`�~F|{I��h�W�b9�@N���y&��W�=�>F�p ��g���~��[���yoy���7������ð~�m�%p��p#�9��C�"EGص�ځ�:w���j���d�h�A�X�;�Ɯ/��'tM ��cҰ���4�6�)jʚ�:Nt
��լ��e6ߣ6-��B�h�.����8��B��p=��$��9���/��YL9�m�`�J�X�)"һ��1�'�f��%7��5���d������;�KDu�~��7�cM+&�BZ<+���U��/�������.p �t6�I@�-��kB���	�'�䁔%v��;���O �K��E��l��FjQ�EZ�
�����O�W����s��k��:6o����C��X�������]`�e�"�j�9{6�ɳ��	�"�}I╶����L�É
��LRŎK�y���n�"'R�9���:q���2/��n��!�c.����3-�_~��;9$�����(�g�e�c��(:
�Qڒ�gO�ߑ�,[<��ٿ/\o�|�����yLX��R-ļ�ad9	�F��h��C�NS���F���"f!�a?:���J[��h�W����46w��KqLV�K�)�����c�JMv�>'e����{Ђ$��1�'�1��υsX�}�V����ÿ�-�	��U�&�b!��!`P��EL|��h��./b�u��7{����"%�J/�֬
���mң���8,Ɵ�����H�;	��R5.Q���
Z���JL�SG�w�Iy�NT���g|�2����D��~RB���e�RB�8:s���A�^�C���Xr�@`�z��xɓ��u�@��0��>d�h�fԅ���xx`14�6~)�W3�����7b��	E�|�"Tq� ]�%�:o��"� .��E�_a'X�O����5*Lؠ��%�s;�	��^z���K]�,�q�������YY���S�K&V��VM��+���t3t�[2�!�vg#Qs��p몜Q@o��zuZ>���b�!�}�^��bDE�3Zhf��+Ut!�t������OeV���$RL��O��43~���s�}BΑRKfL�
l]����F�hN��V4DV<�O,�֥ �o��z	��r7QG�PeZ?��YKI�D�ٍ��8����^op�H;���`��M��`f�ZI��y�K�Y��k�%��&6рڰ��G��Y��x�#�h�#��3#���n	�m��?��|ir����Ώ�R�H4�[�_cՐ�;,I�,�;��/�<[�<kO<idȾ�μ�s@.��x�5,]�MQ�!�����v����2�4>�g���M�U�5�ٿ.@��n;�9�~!l*�(PY=���%"|g�9�M�s'f�ᶺY9^l���q�w��ܳ��� �|��/dǇ�)�;��{�'�Y��Ē��4��ă4����@*�
�[1�2U�V�����ӁY��Fo4��
�;Jt��ܔ^�ڠcH��L �Jg�su���i%F�T���\00s���]vj���h�9�?��T%��3*���ѕ�g@EVh ��3sJsI�&���?�A
Ԡ�����7-[MK��}��g�g�ɯ��\3�v��ɹ��� B&2���)N��{W�`蠠鈛�Q��[su�H��G{��v��$D�0b�4���.�K��y8���2����:g�ƯC(\'H�5��R�㓓}�������g�*���4���ڵL�la>c)y���W��Z<A���X��>��誇�����r��ny)O��~?��`"$Ἢ��{ �T1��x������C� 3��k��vP���Μa��x��k���Q��z���.��l�{���1����ҟo�L?$��S���9���~����뮖&���<�#͋�_��9�M�f�E�؊�z����*�c)Ŗ2n��Z�+ϴm1GWZ��ه�6\J�ڧ����SP�@��h�z��Ȯg>O��g���p0��h��d�h��QB�0���^\�w�@k��b�vè�`�rL�C3<�d�������/:O��Ǣ-<d|N�0^(ʕ�@��mU[)-�X��=��!dl��� ��SXg��Ύv�I<�ě�˴��VT�`7�ϼ��ƀ,��˦���T`�{t	�Ϝ]�B�ߪ9��z�j^]/6����~c��U�Ā���h_�I�iW.����@��*B2�������bC.W��������T'��<��x�����<d�3��O絺z��
w�=��\�x�b
e����˞� ���3X��z��y&�|�%�rI*ҋ��%{��8v��7	0��HH}�C��fCz�;'�j���@� /�����;S"�}��e�F[(~���Ĩ�;��To��\�S�v<�78c�)
�C���{v���
��`p���0�>L��Y�JL��ZnR6�ή����H^@��w���onT�M�,�b\Hڂ���0��ŸZ��/C�PLhA7��(g%-��&���4����H�k���m�}l�m��EɌ�CL&R=S������cr��֤`lL�GLY�b>�����R48�@���4��/���ڋFY�_C�j��S5�k��I��b4�U�Dݶ�Q�rV�T�b�GΘ����/��E�	{%AG���2Q��*N���\��A�X/�6�g�
G�+�nA�!��%��p����"{L���'��\�F@ٌwR�ѫ�ǃk�~����u�9{�X7r��W���Z˻�C�,�3��f�o'%m3���9U�3�{tݼj���q��%����'�O����9F(Sݕ�M"I�"�0���Nxy��w���'Q�S'�����R[����A	=�r�R4�r0M�T�����K�w�oI�}�T��IYY�@�T��R�fS�������W��A<E�� ��K�I�w�O^%*L_Y��[��7p���+!���п�@��{���-T���5�ٷ��R���S|)�[��|!�q�I��WB:�
�A�	ҫtQ�4e��m_2u1!pN��/��?�?lU����=`��_��Z+2	�tӰ�a̩%��/&�6Gq��M��1�cFk,�_"~� M����"���±7�4�S-J�w��䯄�h��ݙ�8I�.�X�BqjGP5F�>�
Q�<�|lb g�N���Is&�-��~��r��܏�������3�R����a;T*H���V�VQD�^��g옡|wgᔺP[dD�7�TI	��,ײe~3�� �v.LF�a|q^�	�J/OL��l'��x��EY���_�і/D�c*Qm�D�8�l���_��ƌ�J#�:��@�Z�4�0,��+7@�:�b��6EZx�V���[��64�1�>��2�#AO�b}�[�b��L!�d��ShC�oC�CS7�7���yw!�	��.�p,�ȗU-�d����Ywc	�S: 1�ö�rY���1A�rDֳ  7x�+���轣J]�bQ��$��O�"���^N��P��^x�(5T�@��h����Yڰ8�=6�n���RآFeh���jk��ԣʴ�E��:hX�t�(�WT�Pc�f��nTB�B(�}�i6��ub=���E��@u�����p���m����Խ#YG������1���$�1!�Ȟ�:���ח6�ǏY�G��r�U�=W{!b��&�yچ�-�n�{��d�4)�ds�n�tI�~7������<i:�]������󹩅�r� 1s���6o��=E��>���71��_���{v���J:���LQ������n�j*ϊ�?=�~�@�E��LDR��!/�/����~�]A��C�7_�!gL��o�N곆�0��4H��~6��#1� �oDw%��h�S��o}%�>&G��_@ EE� � �5gJ|nW�W��z������+ۋ3����Qz��na^e��˽o/��G�D�#�@�Z�f����6���c�6�O0g��R��}�9h���V�s�����dY(�s#z���e%R���/c0֊����'`�C��"�Z�a�C�<��eL��&t}�(�-_��ƂE���ucd�8~�J���vLH��/���e�g�4|Ёa��D�*%�QS�'�Ì�W��\_}�8D֞/�P�������*�.�R������?
$�U�m<��6�z�4Eq��ˮ�ݾT?e(��`7�Jӣ��h��مK��8"B|��I��x;jN�����4f/���s7SA7^?��~��"�J���w�^Ls��F]8Y�n�5��mE��b��b����|Nā#A@�X��A�J?,w���w���C��n7��$�B��ᨡvš�a<��[��N�6�?ּ���e���s��#ٟ��5�����FS����i��C�
����m�l��jN�-��I�� @WyԨ��c������=��st���Fh�-�?�$���p\�k�y�i��8������\�^��U�3M&��l+}3��Q�4�!�S��P��f@�
)���}'k�����cNҜ�GR!�@kcP1��̔���a��]�|��y��h�OĽ������R/�f�M�¹�`�͈��\�K�(ያ���;c/�|m,�-�)ÏQ��L��II�j&�dX����l/�Ǫ��צ�(�Yčgߨ����
~vW�(� ���m3��r���[�U62��\�C>���g�����8M���k�2�����+F�:e�?�dx�ʝ�}O�Y1��z�����L�������Km���୑]H�B�ӧ�7�c���Wv�F?tl�����lӕR#���������r��E/���Q7�/�WZG�l�;PO�m��[������%a��Q06�l��ܱ�_����YJ��1s�F}���1C�5�"��z�OD�_@|��^��b�PD��/@ X_�o��D��Mޥl	[28�GXˉ�p��f^�F<���	46~�;5OG���_k!��v�M%(�J�`��Z��?\��J	��C���D�׿<y<�x�\���<��?�������Jl�%o�~�ho�Ju�V��/^�+���b#
�Z��z�rv��F��N>�X_?�\�{>UG�j�2Tc��߯c�;�� ��٤_�-Y�H�k+�&݇vDņ�81
��1�W�U乊����@�^�����������x%[�U~)a�Bٟj���l�Z��x��Ě&��i�C�Fp�Pu��B���zN�����y^�����.x_T�M?˄�\#��o��C�t��,����D�w~·���[�ڮ�čTDH�{��u��o�����m��$��W�v�*]Bl�6ꈻ���ҕ)��7˗(�d���+��	i�6��?��ʈ�i��,�7����Dg�Qyߖ0���#<���>
Vz;׌�Grgpc���{ɶb/�Nc;�X�r�i(%`�}��Z�3u��{{C�o�����_5{y�2H536p�vW��[��.ůl�	C��aWϠ��(����A���A/xDtj��'��-b���I�c�����o�}���>M��J+$U��og��/�ѥR�(���=-�IXr}J+��k��~��z�f�C0��'��*�"�
o�7U�
���>�Rs����n;$n.ZąYqbKƁ�/��KS\��=`
�`gh�*::9R��	��}6��L��^yu���O�=(����w���Ȱ�9���d��Ʀf#��R>s!s���he�/���Ⱦ/�x����G����G���WjY�����<����9�9X��ٍ=�pZ[�#3sp��(��{�gx��ϣ1�ܲv��:����pC=6�D)S�u��nV#I������|.�+|��_-Œ��$jP����j@h�+~�~�Q',X@�	�;��]�0��+;N�<c4ؐT�fE(�[D���'�ۛI�^�,�0�3/�zθZ=6p\G��^���~�a�(#{��&�ۊkD�������F��*�/QIQ/�BF�ȿo�G�~�k�rr7�&�dh+A��s:�DC�d�;��Ϻ�:�+I�}w��l2/p���_=@T3����!l��"9X��M"@cڷ;VE�H�d�a�������B�*�܃��L�]|�*ufz�N��V!� W!{��0��T��0 �1��$���c��7ۆ+1kw��&��jZ��`\`j���&6X��ڃ���_�k`��9�����"�q)erC�U.@�r����Ck��~_� ��:`�����b��{C���Ha�w5�Ϩ�!����3�4�������y�
��:֮I�a��S"T�����"b�I�ov7B�D�D��Pc*��gj�?0�_0GJ;��?�)O�iV���0V�_��x�CeK ��
4{��B/���gg?��#����ՈʽA������e�.����M���M�i/<c�lU�ð��m����d�$|��61���1��j�kH���(j(l[V(}l�{��w���˟����#:+s���op� �'K�+%��I_�-�sW��:��=0c���S4��x�xj�N0��b^J�A������C��n�W��w[�o���$Ҹ���g�|/̼=��B��,I�-ZT���'��ϔ�ӝ����Yxh��FZ�2L��IȐ)��x}�^�� R��4ǷЧt�ϛ�gqB���������L]-Y$�������j�I��h@��]k����O���0�.JU�E�悯�|�|r^�>)��B��H<�<�a�6�t-N��F�9_V+1�Ms��Ȩ93�MYlE�m!`���m���1=�b����x����WF �t~q,;��e�A�_�3�$]�����"@(�[^M������l�K�z��&%��bZ��݊u�����ڑ���6�:�C�rl��S�yɒ��0ӝ��Eav)��l�/xQ���u���"�%��h�o�q�JU+3��!m��Q��?���%ř1�|�&d����?�4�����TF��Pn�:87o�e�=A8Ń�%�>=t�ǹQ��OןZ '�*~���l橆��VHՀ�p�7���{t�On|�m� 4�e)�۬��q{�fW�Pմ�;��Gު[k�z�pfX�姛��lWP`x�A���R���h-j/���bw�/s�0Xa)⾒g�Lӛڐ��M�I���]0�0R%2����Y��a�:q4�iA�~W��P��͍'����Ya�륍P5%�KJ�#��'cY|@�<�,�l��"$�tY�X�G�2�a�V'�)6'?�����w	�*�L�Zw������G ��)M�&�6��x�r�|�$sd�~|�8��S� p#)"��Oi���J�D&���~��Z�;���/Αq,�.}/}�f�#�E:��}�%#~Q�L�GX�_�����
�x����C^k,1ȆWH߫F�/P�+����.:�!t*'��(R���^��g���f���N��ɏ�.Of����-a���B��s+-B]��<�R!I_��Oz�!���=��p&Y��tU}���ѡ�$�fY8Qԃ��&s�ak��DJ�:?�j��1Ѡ6Y�j��֞�?T��*x`�SK�$��a ��d�ڏ��gdz���<dXN"��Tl����ӓ�����sј��>�NE;.yd�Err��� ������:y�(��l�\��M��*Q;v���'�$�m��x�����~�!��I�/h��@�-Ȣ�ʂ�z��1c �͉��q�!_��%u"Ib���O9V̱)�E?]2���.��94�0�����#^�*�q��T��/ ��ў�.���Fh���Cv�v�3�wC�!�D��d��b�����BA-��UWP�2�m�
��'��q�lb�O������q��ֿ��ޞq]��,pD��+��~�VM�֫a�����G�`ۋQ�;_�
���2Ɯ�cg&����("P`O�"�H�ZK�}ASa�n��_?�&�!��M��2��a�Y����G�Un߮�l��-���O�X�ǊZ���y�l�$!�����4�֒�]���ZxW�v�	4M��u*���
���0N�ez��*�qNNP;�ޞ����Ճx�qz����2�݇��' ����Vj��\���C4"��}�x�U�&�b�(�~��VE����4l2~��i��jn8���ץ�����i�+�`�xXO%gs�߶)j�Ԭ�,X1ej�(6�%��|���	�n���;��>RľN��1gX��Ȝ�%"m�Z�:XY����YyY�������d�!�ڞb��@�]�Z<?��\!\�H��(��:�0�Sʪ^ w�����{�q�<,����inEa[)5x8�Z��>ɥ�,<�Oިe�{��Ц֍�«KW���?��*G��{2�L�.r#b��m��b�s�H�ޯ�$���A�Hڤ�*�>�w��4��i�*�
D����"|E�q�����bs"�<k=��Ռ-W�w01����B�`���LM�H�9��}��+�;�4�h��P�n��j)�ټn��?�ZvZ�����Y"~�>�J��_��!v�3MF^��:;\~��U�OC�l�
Az�0]���WD��Xó�AI�RFY�d%�U��Z]���
a�x� +C�����3F}5Q:m\���ھ�5�M�C,�X*���x�L�K�ï���^޻淀w4���	�^�a����+�bi�!`e�w �r<UQ?��f����D��͂"��q���tL�6�!��x�LP���1���Jӥ�*��@1W���&�-����+��%�F`��KVH���K*2��->.�˾�y�j�0FgF�*�JU=�Gݩέ��Z!�wH��M$��t�<n)��f��*�*�X0�c{�%�)J���jv%��{g���5�6����b�(dzu�&_'q�Qc�����.M'n�t���h�r�ʕ*(i��ǲ�t%����6�XԤ�k睄�y!|I�Y��pAP���G�}������RM��|����v�5�Ի�e�O]��L@k��/�|��b��1 �9dגǥ3|~됗+TW���N��S-��?�XU	���"�E��&���G\Ի*��zH���v��Xۉ@~sKfk
��H2�ΰQ�m�KSq�\cMu���c �9�3�t��DI�zΪj����tx��{	�([͞��zN��_隑���c���5�_'#&���
c1cۮ�7۲t�w�Յۑ���M��v�N�(]%ݏ����S��)�
��q/ q�O8��2�Ə���Qj�<�{tȋ�F��kZ}ޯ�S#�U���"��A�����Ȓ��6"_�a�����:̇7Gy�n(Aٴ_�ህ��B^�z]F K9 �$Z�(I:u�+�E,��9��[���K9�2p�Hiu�җ���>[U#U�y��l�ϼ Q"������Mzs�2c��4���T���cSr"�G�au&N0�Fe����"�[�c*��X k��sD�[��oT�,%��N���ǳh��F�E��u�5w�r���O�۽�A��M�E�d�5s ��:�E)���Y�V�N�Ogj�X�Z�l��~�f�Yٖ�|ؙi�1^���Y���.����n({>b����L8�6��n�l@�R*g�IA�����|�
p��
��j��_f���#��7�_���	c{�S�~IO==`�,뛋6��h
Oǣ�'�)�w�,(<��a�ro,W}�am	���%+G��C2���q��1jgwY��G[�*�Km$^מ����v�3��pRR�<��	Kf8hN�~l!Ҹ<r�e:a�|���K=ض�=Qg��-AQ�󞾘��eJ���_�~����Z7�Ebn�U�߷�2[ꎇDq6bam�G	0�Y�PU70�qIN�U� jS��*�	_s��{�$���s���p��c6�x��>���M�:�L�^��
x�aI�˂��G<T�Pܛ5�?@����̨m�U��)0x?�a�����M�}�@�kpY�PU�_��,)h�Yr�"f�����zy�
` ��qA��p?ǂ�Ɖ٧a��+�y�`q�E��:�U�Q�Dm�@z�L�rGD�X�6�r��Z���*�;��]�{W���9{r�;�u�OB�N�&�X��[4�φn�˯u��l&}���;���1�w�f��5�ɂ:�㖙8ī�Fdד�e�$O����2yeW'��OТླ������7��mc"�W;j8qv�Q,Yl4k#	H��d�L��6\<���W�27[��ve���i(�f.���4�oML��y,^��)M��"�D�x:A��{jU�����}ٲ0��R����&$��moʨ����j [$��G��1��2I�ba��Om�E�|�!t8['��8v7oG��v���GA�`�d��[fu�Q����)�s�m�b�K �_)��_)8Z�/���!�Icdz�(0)=q��3�8�m1��[��qVuB���-~x��dpՍ�M��׬ź�I�[�[X�1^qҨ,m�m4c��ώT2�>z�����y�Aa�W6I�ͻ��M�fܽr#��L�`P�r��wӡ���@�?{�!�����A���<�q-s>�Һ��e�P����w�7bE�q�H�1��.�9|��x�����?��3��w�̡����J_�,��|;�bUԜU����>��%w�� ���Q	v��c���S�$�a�wV��� 5�H�E(/�b"���P�]f8J"P�x&�1]m$|;N��i�`���4T}Z�9�a^�3xﲊ#�9D�-*��L=������ˡ�٣h
�c͚σ��]�nօ��i�������S Ep:P�ɍ��*�"��"�<$҂��Ӎٚ�	�*��V_���iXsV�s(���GQh�HЎ�#��.ݸ�N7�Īdt�XV"C�.�����D�/��U�"�yKh=�E�sZi�\��(��6��U�JO��h����|>�K�\�/�������ͤ[b���҉�/X��>��E����z�R���W섭W�������N�p�n\x2q��&mh1J��OA��[�X��W���r����B��l~��[VɎ�e/O�(F����dɿ�u7\�]��N�U, �w ��ƒ͎����XTحb�O�A����|�|Nǃح����u�WK�aW>��K�~[h�8i.J8
͝�Fܹ�_�N�ot��)�9$�
,���У�������S�e�َ�i��'�����|�C����Vc>�0�����K32�Mw"�/́����6G~���}�B�Q��)5�C���f�`����ї��W��B�����Ur�W6�!�m"��\���ȖMWh:i�i{u���^����i�$ ?Ǐ�Id_��I�o 8�@�T	�J����$an�=��Zl��+�_2�y�1[Sk-kPX���m�N#���4��5-�S����zVkX��Y���G��8�T�.��)҈��.�-��t. Ɏ�2J��+��� �i�����%�����1䬳;��J���K���Y�$���v�Y��s��f�pM章喙�2%�$H35