��/  !5ц��Fc=���F�jgg�.!l=l%!�uN��S^�6�)�Kgn���H8�`�BH��RXMTl#�4N�3����;p�)o���;�Xu^�V"΍I%���V���G��!��g� ����A=������4��Ó;
����6F{į��0Ѵu�;o�Yxy��t��Q�;��J���0��VkLA��I��v&����+�U�"�X��h9�*�S�R�0s'|��RL��M���î�̙��1k���*h?�e���\p�����g����?�z���*h�_ӫ�ME�Fuօ��&��W���;�yJ�{�b�,�e���M�<�2jBR����Y���w�G��'�V��p�K*k���Z���\�����@>��t�&��T���78�Gy)kE��M��M�ŜM�ź�Sz�&�i�8e��x�k�?F�)[:Kf��7��Lh��U��m׫3��Tt��WG���k������}�G���g�+<�1v� �}YN �*�<����-\��[����2�� k-C��6����v�!i���7�L�%�I���� GG�GU:q�i��]�p��{o�^�F���W��gr��q>�oE��'Ug��0�2��	7������2]o[< �����8q) ؛>+�N��\��Cd���DCJ�!i?�M�H`��Ȯ�(���\u:_���s۶\�]F�٩��2�)V�Ȥ����N���=�ې�Vn��遑U���5'|�)QnN,��艓�|�{�pӭ[j���-��7��@Kґ��Zz�m���7���S~?����s�r����_��yN�eh���E��؊T(���'�A�%~����l��j��T	6�
_p5���4gm0O�hs��Qӱd�hA��ٳAV�R7Xv�):ԮB$�f��ktPN ��zִ�,K��R����qH#��,3���p����螝O³�6�kƓ(�N�h��Aq����Re	xn��v�,˩�/�U"��.y�ֆ�����Ii�sNC644P��Rg��w��G��^W����E����1�i�a����>���6������߬����ƭg�y\�v��D���>֧^��-�,ԵbɇLO]7�H�:���u�U���o5�仸kOڟO���C�������Qa�2 l���'���x�:"�z a���>��c0d-�:�K���˵����s�0�0i�OTf�%��kN
��f�r3yG�y���P�֒��7�z(n��L8�<�:b��ݼ},�yY�_R�$��������0mo��!5,�����!nq����| Y����JV�~���_��*L�~L�+�鈴��d���t�dVq
Q����h7D]5�5�����V_b��Qfr��jzi�΁k��XW�v{�I�Xf�	wD��~k��)A�q�ՌK�L;�D�˓է����9U�ןP:��w�!j0
1	�?���O �Lz�����tI'�*V"��=)hęF�G�E���
���=6���z�7�o�S}�f���ɏP����y�R?�S�V�s�ռ֏�|6��"��R$� �J�Z��pѡ��l}a+��|�Y^��L_w���JN�7��顮m�0Ͻ�������;ſ�)WW���u�=�X��d�xQ��;�40rL�>ł= �_��.Q��+�!f79�%ڣS��wh�	wV��W)�,�S���v�&�(
�h_O��U�<� �v3{����6<�m����kp:%A���A�1���,�c6H�8<W��
�"*�*��(B׾-�uec�m'�k�K�dԪ�J���D.T�3���:l��%���'�����I�.���h�ٹ�����N/>��,�ˮ�?ctu�b�ԧҕ9���(��=IA<�����[)��'q�Y?Ȯ�~��8�#�ɳ�����<�"`8d��\ꨒ��ڦp��!:͟	Ĥ���Y�R@�#�?��Q}_!&11����Dp~$���/:4aT7�h�l�Kq!h��%9�q.K��{�*��q��$�
�H}\2*<H�0G7�[�������ȸ.���)��.n�lp_�﹛I7o�&-�1�q�:�ݨ�N[b����
0�A�Eؗ��������j�ad<�6���@Y�D"��,�����#�X3����[<�!6�,
ǅ�;�
�	����`��J0)��!O�t�O�����j�ϼ3��J����kp��;�~7�T��X��M�Hۯ��-vg0�9��4G�N��a�^rq�>���o�����_^�{D�܂#�����3�y1�BI
)����y����9��H�3r���`ᵁ�ɦU��(~�O���K0O8V�~��x~�c����h����3��^���:�h��l�Zg�[�G��яՕ?PA��3=��d�uog��8Φ^�6ZP;�q���3s5Y���L���I�&�ʥoΡ.pw�i֪ů�����+(h�4Yo�B�޻�����<.�[�ɝ>�/���nEs��(�[ΏP;�h\
3��;z"�R08���yp�s�}�$�\����#b}'{�"5��B�R~�`��mƬ��ő���7�S �����i�!wN�����W�j������+%Q*�l~�:��A?��Q� ���T�a����Y�[H�~�!�\�-�6B�Q�.�q���iX˃��R�A1v�C�I3^�
�#�DX`*�J�aS^���kV�N.��r� o ����q6��(���U��-�x�~Ϊ7��s��E����]�gX���i��j�&1�����~�̰����S�w[o+�e8�}@�q����Z��𢨺W��G]�w&?s9A�Nhh(�!u@�����\��΅*�.��]N�t����*	75�&����2fO"[@�/ ��O��R��|B�L���e�B\o�;!A��rh;*�����f|\�v�ږ�����Ux�5��+�?ٳ{eS�4�l�R���G��L��IWL�-�Q��}vq�/
�M�	�X�(O^$��h��a���0�
N+�2�W���E�n�FĪ�0+�ջ��0a���C��~CjA����~��n� &�U�"N��Xj,���D��x��d�h�6�%��˫�%�����SzKyu�74������ʯ.b�#�F����*�Q>`T�rEn��%#c�((Ț�
�������Q��5D:C�.19K����U�7f(��`顁2��<��Y��Nv/���$����C�S�X܋%� g�AYE�U,�d�Of*�x����1�ʰ%7��Iik^?	�sp��I�|��Ѩ˨�������kE�Ư�@�3d�0`h'	dr�@CeԻ��	��tIq,}��+�Z�`�ɒ���2]J���%r�D���� ����vp+rsd��R���Q_TU�~��L�S���V� �(
���SM굚M�K!Bc�X������Ȣ#+p)������V�%�z�u�.�i��-r#Z[�W4"}D�  0v�ք����z��yR_Gv�`����C6 P���6XA)�s7��U�/�[����\$������0�����B�ɶ���o+�. ��u���⹐I磮N�st\�Z��R�ivwBi���I������g4��08
;>���u�F����o^��tWp�ڄ�\{���I���s��c����f��B$:0\�Z=TJ�('�6�{��3��I�'��]Gu�"R��� @�	G��۫68Îw��Db�rx����E�K�2�w�_X 	BLq�/�帡3:x:�o�.v~�(rkS!��z��:���y�rg=(��A���]�~[���wNܧ�;O>v �ZC!~��4���4�Yt=�b���^��?�~h|Ŵ���_�|`%�u/�P�`�,m`��a�]v���ޛdERh�{�=�����E=C��_����ܲi�� �h��\vN:���9.������n;!_�<dzw���7L�ă��ךX��'�����WdF	�\:.�ȟx�6�Z�m � ��\���Lvr(P��9��5km:RCvK�k�;Z�E�="9����!|�<�����6�I�
rܗLK�̾�:_�@	�7�����f8  c��Tk�_ �R�A�CP�l��C^0�  ^�ۚ����	�)7��;�;F�s��hX֗5�^�o@ݍ���EF��D���5�9��;\*��:ۃ��'��#��h��8[���Z��b�K!]�KLKX����LW��7�.13�!?Xr��]I;��a���%�ץ��ɧk��vU�C)0+�������mZ����fi Ѽp4���tD�y�,���i?Q��'����aAc��-���>��D��<r���I�p�a�Yt�ݮ�jS��(4c�����dt��� r�#���L5�Y��q�$��r)��P{���C
�r O���+�s�@����+,��0�p�2ԗny�b�B�k���˹S=�0K��r��|7,T�$�L�:��BDIR�`���Q29��	j����	�*+֙%�=����Wy���s;0:���׼q��z���[�z�n��S����'��=��Dҭ�G!0�#陰��q�&����@9�"y��{�d0@9��ѩO�z5�!���ql����W!�O�͟:1�_�~��(�^gO�p�"�·���P<E!� �iC�W�V�6�
�Y^綻I2uͿD�Z���KT*���������bڑ�����{o%���.�$���e�\�m�EQU��Ldv:�ε9�Aq��K�6�s���.��9��ǟ�v���^�i���ѿ�(y�t�T��ѯ�~זQP'"�PQ=����L�hnW�~�i� ��W}_K��/�-�˄,H2�;c�9;�j�7'zb��ɳ�.�p�֖�jMS�b���F1%}�n/8�(�CN����A\�%�����eU(��{헹�IM�pK��������A_=P��uP�m{��3%=Tc�B�E��AwS����ڇ�7CO��Uנ
�J菘$�'s_��K�i]���_�U��uY{���o�]�;	����H
�eA774��zR���w�>��
-4��CL��D�8�z�B��Ɍղi��j(��F��#dc-��y�\��s�t����1C���A6Ph���o�(��>�;���o��Z�!%/>�V� �.?mڄiٚV�s��@��| ��4vw/�����)�KON ����fg�1��t�⤼"�<�V���7�L�8�z�q������&3~N�>3O����4:�<4p�(v"]�vށ��F$X�{��Hv�2���j�!�_�5�J��z`[����i\H�U��g�p�=k�T����b<Bd���s����y~p��
3���t^��s���'�`Z��b�EA�0�>��s �w˿y��}N�,l[48(O�nU�W�V���%a�oZV�u(\FwK8�0�nM�x'�~��i��m2��W�Z����.�����D�lx��ۈش���so�(FjGBBk�x����)hl਱B�ָ+�â<k��������̗x@�� Ѫ#f�O�����4�k7�m�;��
�g�[�
�<��+ƚr��F�u*���`j%f��ʪ����Z�"���h�J։_������Eǫ�	�G���(��I��w��$�vW/����_V|-���m�%�P8�5KO��P|JT���8�O������`jzo� rMk�� <�eRdr�\>	lsA���=�Y�|F��J�}����x<��,j���[�hc�ʚ�sR�	����/��2,�|�Iΰ�ߊ#tq��QsqܛC~	s�9��N�h@�#}�(%o�B74��u�����1��q��'M=d��}�dvղ��&��YQ�*��/7�[4EU��@n<~�b���@�6��=�l��R�V���L�E����/[C�;6>HR��f=K�9ri�.`����xYij�(��U���?om�X^v���a�pb#aO�3��v���oO���{ǔ�0���,C&&m���B�?Eh���j2149�'�����>2w9q"�U1f�D�I�e��(ǎ��Cw�<���t̴?`���g��`�t �� �����%�p�t����ZU��u��u�-/��4S*B8*��ɶ����� L�E���9��;�J lT%8�4*'��8#�-d�G�����+��W�i]������KA�p�J>�_D�������Pɔ	�a;Ïx�̧�\	X�H��$,	S��e��[I�BY�{]�w�.���t����%�_��\0�
�����ﶪʅ��&}�@Ę�C���1�����Q�>�3�Ju-Z�N���?-ři㷓��ҕ�BAVm#,/@+�a�&/���aZ\;�j ��0#�޶H[�����������s��'�d9����D�I�F��:��q�Qa��T��Y%v���m�ؾS���.R_g�J�1�{X0$*�z�����חMavƑ[��F��|6��r�yE�-=X���d�gF�B��eモ7�F�ǣ�Ld�;�7P*rw� ���Ȇ�KS}����̄[��	D��e��:m�yR@F3�,�齦�$��1�pE��@<��|��ԡ֟�w`x>.w*ʬ�Çӻܐfd�lʺ�5�Js�[1�8 -��p����c�ݼi.J���w�:̗�'�f��+m� ���_�A��E��U<pf�.j�7rױ�Pa̙�y��JM�������lYT�'�[��-t��+�Э���aE����?D��f/u`*���g������4��M�ܨs��JK�4���0�at>)�6C
��P�<Q��4pS<����z{�����t�
��P�/��H �i��D�SH�x�j��J ���
_^�VT�R���d�"�02�ws`]�kW�V($����ح�t]k�|��܌	R��F֍PQ��k���=+��O$�����`X���6� q��T�ϟ�d&=�N`�t7�5L�R���-]����jF��2�.%��PV��׻X��P��`P�X�0<��E6���n�i+��#x'r���C�,�������[�iԟ�u�m�_SL)�d�gԫ:�W�JF����b��,��VF%e2O8`�0�$�$�|.������{ӝr��^���}���D����v�Vx] m@��֝����0����B#�M
���Io��X{b���LM Io�4�
Wn��:껈 �\j!���󁏥����3�yd��(C��%�
��@���j�Z?�b79 �v�F��\o��� ̡uɢٮ$�lb%���f�*��N��Y=OI�8��欽f��S�#q��[+���K�Hq}koaj�ʀ�SEǇ"\S园����uw�w ��"�u+�#����'8�;�b�#s%�_�*��
0v�8���Rө�_�����B)	`�n"|;�$R-�4�D��Ʉ��J��54��i�����`�Y������a��*�̫,u�c��-�f�{��Ev��X�� ³?�܇�,��Uz�r�xSI���5����1(õ�6S��釸��#����A#>�]{��L�2I�܈��׍d$+�\#9�^�-~U�Q7��"â�ɫڪ�g��Ų@c^����ɾ��u��y\US*�0��C��=[�r�ɨ�������mF��#�mθ�2H�;��V+���ƈ��:o����4Ll�e������%AN�'�b?g��G��5`�l�B�F�Q�|�o���)~OsE��t���,��5$5�.n/r�W1$CZ6f��C^'��(��j�k�v���S��m  ������.���a5�aH�zo��7#ׂ��k�<i�Ro�c��6kmBB3:�^|Qa���D|P�,�:�D�*�b��5��\���%3��l�b:�*~�,���Y�E��u��n�ٿ�TaY�3��\C>u�w�ȑ>A���'GR{�YkL��ꥭ��d��`{���},���Ee�>��Yig����f
�&-4Б΋��o�&���0j'p���pQ�u��R���]��c�<8h��iS����jH�	g	�mX���	@�:��|^pi�!���d3�v����F��nkno��W�4R�~�;�oEE�/9=K��Թ��ϽR�"X��K�����9�� ���z���V��R+K=|��a�
{�0V�pq1	?�:w�dx�n�A��&h�EZ�o�\~��������=��1���� ���6nqL�ڒ��ڱՙA^'k�=43�S��H���.�:�U�br��u���.n��"pf�A&�@�*��N�����s�����b�Z��3di���߹t����o�AM���D�c ^~i�h����*kĳV\Ii��!��G^;O�T�MJ���BUToMuţ���^����-X���Ch�_F��GW
�I�=d{i�y�TT�O@)`��[Y5�Ӆ:X�g*s�<N̜A�	���E)G�Mݜ�Z�Pj
���=f�x����Q=�`ݭS�h�]�5G��m��?�M�	������6����qix�S�7�@ky��Om7��F��m!qWK��O2"tzW �u�t�-|�U]LYKk&�M�
���?�d�N�4�&\���%k����O)�]<Rz���s�΍;+*$��o�9s�y�@���1(��Ѱ�&���_���K�1�����W�Y��4`��^��9w`�`1�)��ۊ�µY����Ue �Q	���!+�w:ݜzY\���v�{��JT7���4�X�pA!������U�-�����!b����+�Y6�����]-���Ƨ�jj
ǜL��I̵�
�G�Z=6�w3��uQ��~�� v	�F�#dP��Fw����`@�����F Ӷ�8�b��)x<�������cұ��YW��j�t��C �x�9\���0E,m��c�/&�pS��"�W�M�ְ
��Dx�l�C�>��z�bP�J�D���M��4XkDU�9�c iW(TL��9��v��7��Ly,rpiV���g	50?��Bh5_��1�Z����^]0�����F�� 0���?_R����6����B�rGn� p	���`��x��@efZ�|�-}�[0+��B��OU���C#�9��`�|X����:�u��bb�t7�e�\� �9VCv\q�����3������\�<3-�Y�S�T��w\�:Rg��]Aұ�8�����9:8Ja�Zw8ٵKIL%0��Pʱ_��a����o~���ۼK$��P_�A^'�<�Г8��+�EP���<Š+҈a8vY�%��ꀠ��~#D�1����R� k��,s�9S�=���AB�ALr��e��ގq/rc��U2���yw����_�d�X�ۚ"�#���?�\(6*:�0Q�z\�[qB�Ѵa�e��Ly׫e�e=gRqT��H-.�̍Y��'���T#�A��o�CT�m�Su�����3K�<,jat�~�Fi�ۂ6b�3�{���/���̑�<`[и�2��0�%fqgڤ�l��97��ٍ�Xo�G�k�d��5�{<�\=D�Q�t@�L9/��j�/�Te[c��g-(�T���0�����^�
�l�9����ҧtTdb��o`P��W]���ť7�:���߅���Fz\V��! 5Ȳz��edoD�q��ia����R�S�.�>��f\6�s̷PY1��l��,r��U��_�W��k�� �f�[h@L�͑r�?�K��(�`˽��=д�U��"��?G��a(٨�0B�Q�s�����]�/��ێ\}��+�s�T�/��]�=�$�m8�y��i��7��K��+���/�/x��P�ȱ�bGӨ5�5��<YB�����(��U�4�r����7V$����sc��W���0i���̈9j�����;�G1xp�	[�+$$J_�6S�g�Db�NA}��Ky(�ƅ�A4��3����y��������^�	Ĳn�+-fTig̻?È�'7�m}����DN�c�L�Ǥ�Q:tj�!�!�'�<�=^~�Q���m�\����ڻ��L	G��P��"�h㳕�),�CUr[�m�w�l����ϵ����n�a3D� 3�F��+Z�����93Ts�-1R^6g������pD�=����=��mkl��4��2sE�@U(�&6K�1��żw�������4�U�;���ǅ���}�N�]��h�Q��zl��k�c����.�R��	��gŦ��\~�6}"��^�z�]F�%�A^�*C��U�ص��j>�0�#���	���֑��e�2�+D#�z���'04$�
����,�6��![x�G;�M��T�]��mti�C ųMB�b�l�C�VJv�2PB�0y�-`�Q�VS�_�f�yG=�ۦ��l��io�"N��������+��8�3��y��-�؅7��	1��zYmLg0='�wzȹc?Wi#���e_vF䳒Ok<֧B<"M�<��'�o/�y{��{�&�X�%3���Z"�V��lm6�UkLcM:��<%�]��1MN���wk绅PY��I�\�޸��\Y�<H��(����%gwM%�}�C�m��'t�T���툮�f��jk������l����%,����J��zb����n�ƱW<�u�/=k�|U4�\<�4*�K��8A�qi"p��1�%�i���'�i�*߯�UfHx�kr��F�L��Ik�aۜg�������Y�s�DYX���i������g�ͫ'[
���+�4�Hdc_ n���O�fcOmc�>�K�=������H��f�UpbT���sh��#�غ��]X������=����W��O9��~ ��ׁ7��b]���é�Z
_�����@Iu��i��I�C+S�+0������̚/"YY�Y� �&i�R�'����86�ۄ��v%���yW�?��͔�"hm��5����]�w�**WD4J%�<.`����@���1���x�� �0
o�?��K���`�]�>K�~^�E�4�����Xi�-�8qE_iDg� �=.wz0!��M:8��e�o����p��7�.�s�B���8�*���(��.�?��T_I���⇝G��k����QE�-1��I*��,94(�(w��
��`���l@8�A�(~�Y?�(S��S�D�+�D����Ӏ]$�$!�4�r����y�����NZ,���{�"ǒ<���V�u�8#��K���z���Lgs=��y4�1lXH��lB4�Q}�7:?���B��Փ���t_�!�o�N�*pDJ�󃊰�3}߻P���`���\B2v�eO
�x_{����O�Yq��AP�9�?�F2IV|�bj;+υ����E�u�%dg�-��xST�`�<�9L�&��5�
�jk֚~��Rɖ|�_uQ��jm7�(C���?Mp��\qw�<��A�r%�)�)ѝ��wh;�J��$��EB��C�Z�U`�H��<c?�%��N��q؊���u��_:�[�J^O����Z}w/�FL��F��BMh���$S��dP��!0�tr���}W�'�$Mj�7J�J[�/j	�x1v������$� �UHF_��%�� b�� �nDQ�Ms�~����>	"������ykX�⾨�@�F�`3�N���@�K^�d�ֹI7+-Ă �m�d�X����j��w��z�;�A��1�`'�OaE�?���x�Gn�7�T,�c2�"N���t�����	���(�dZι'�%Lv�"2�	����,{ĭR4�9.���'k�E�7	��ȂO���@"��t�x�q����^ ���ct[hY"vu3����v���%d���'s����X�㵳USP�(:���$�B�#�:a"�;|�Q��(]L��]ε~�_�Z��k�A˧栤2�0�����G��&N��T�-��۹�u��3����{th�k����>�\ɐ��E�#�D^�`�0)K�;߭h�.>���&�2o��@�pi,�!��F¢���Ȅ�����^�r3N|4�uf��X�0�k�S(�=?�Ȁ�K>e��QIO��eƸ0�u�TW$O���2PN*!�Z@���<N��j���?�[�����-��j��Kbxi��G��L���ٖ~�FM��Uq��~fJ�����o���[D��Ds���$�w3ЃO ��OE=_Qê�+��YǃC�~�n����[&7/�A��,��cp��{�(Sٛ1\�c�C+hޯ0�#mLUa|�������Um\�J�>�`�3�;�=f��V"!�qX�c/3w��6��I�a�/�R�4�F�%��^����+�F�f��U?n�H����Lki>�����u�+���0k����I�B��4jԬ�m�$��v�{W�R�R2��_�Z���A��tz��>#�~r=H�� ?�]���.n���_�ʸ2X4�'�Ӄ�C��6�����/�Qy<<�$.ڸ�&����P
�G�-�����E�6=iSN���$�G(y�1
ɻEk2�D3�*�;����rН����s���H��&Shu5�Pټ�݊�$�0���b�����)E]]iǟA�=%�!���|�m��Э�(gց�-�mJ��5���a�)܄�~��M�"4Zg������|w�x9��P�5h^��\���� �&��~�'�M��tA���ڎxoF�mH,@C�����G~��M��.ܙ�v��{�����@bZ�#��c+S��F���xm�A%�,���F�����9ԻpN��/��~�����5+=�D�q��8������طr�Ju��{��ɘ���Gy��.-"� Y����~�e^�a�z�R�)�?��Rx�8%�"�����pE�\G���e�sU����ش���F(��~?�	P��2�ڞoIT� R ��mu�	j�^�H�Ͱ��k���Wjv��f�L�z6�K�I�"f�+�}a���j>���Ѓ�I�#lT�?%�x�w)�+Y/0F�$�Z�ܟ����po	�4���<����'���U:�tȾt���Q���˘���\���8����Pb�Y�8���g������J�C��:c9d�hu�l+!S0����R*�VAEkxs�ҶI=��H��[���l�ۆ<;���qx���A�W�}Hߪ�x�+�w���MP��1����m��?��
�C�@<����=�(�L!�W�/�Q����,��8v�� 3G��ŏ������"���2���}�HG�x�t5����nX	X��ey�M��$�Nhd;���Y��:�a�vW���Bs�7k!_2j�G��Y!~��9���z�`���:�u/��D�n�R>���� �$�E�m*�9�Lh	�D�<��ElJ9����vþdlr�yEtU���_ָ���O!��+Jӗ&Nu C��T�]$���@��(�D	k)V�����N�D�.�n�Miץ�Un��?K�d]��
�^]痜I���w�����4�h��ܺ�� C���U�Q+�ڏS>�P@��KQ����H�X��ݩ�������-���557��gֽ½�.�dm�
�j	�3�,[@K�HWL���ۢ��io��TYj��3�%��2`�ZY��tǸ4���l��bճTh-�8��*��I� ���z}������0��� �n`#�p��ƟtӨH������/�D짏7�h��8�@�+��Qf�_�Ky��WG��О]8����HLvf���%�������ʥ�Ө(si��z���O����V�oÍQ�o����
���DW4�+�0]Md��狣D%�
ф���&�ZD��P.�	 F-V�O�� �vZ ��{ N�-5�� �ٮkW:�>CٗN�*���dS8F�;7���vb��#��O��-�=@f,W~���(c-��e�+�F�8
�}���������a�;�ppO��SdF���ƞ�P��N;�c'	�z�j��Z��c���\�j�N0�nC݌<��.�}'�R�3�ɉ!�h���1��x��%A���Ú-��I���=��_��}����	�+�bD��(l#|�� �9yJx���|Jx�s���Le��1G����MT#�5�e���͒�F��iU6����u�ڎs9������fS�+���Aq��8)��`+c�,nw��x �jӀ�Eu�?mRہ-jdk��f���Q��B��d@I<����0��H*s@���9F�j.<��h�M7�����~߭��y�1\����^U���x�,�����2����T�`�����3k���%T��$H�: [��:���$$�'�t�;xW��ԬIwz��ϳO�����TR�IjM��z)=�� �0���b�,b����h���;�*���EY>k�,���f��ZF�ܸ�������)nn������~���`S��D5v�t�����TƪWX��m��F��j�E�&�Y�]L��>)�h�'*u;��Di����.�~���Z�I��{'߄�!�[�����Z�?IH�����,�T���p?�3������Oͭ�M�nQ�\��`���d@�j�)qB�;|s�ق�[2�hd�;�ԃs>^�H�4�ѫ(�tR��k�٘�7ٕ�nƚi����ws�M!�bD��)S���x��F�~(pѺ5�7�G$���I�Ok�.W�"�raȻŔ�d0r�D꫆a�n�I�� �W���61����F@p,��Tw������4O̕PR�{x�[H�>����U8f�C�%�;薟�@ .�~���R��s{֯��K+�ME�#M ��s@�2��܏�ǳ{���9��(�@�!)O������� �m��g��S���b�Z�SCȥ����`�)��ŋ�ǲ�_�&�0<�ԗ1��]��!�Z���v�y� \�ѡp�O�q����p������L�~���ʰ�8ݱl?�9�	��ą�0yʲ��4hk�_�	�&�"!� �덳�X�����lfv�_E�ƶ��i[�^�&ϛ�&\G�N��$�3�����7z@v�K���k^�$�W�U�AX��F�#ہ�wJ��`��ҷ�|W�7RՂ �΄ڦ<���ת��ܒ�<g%$T<�ˋ ^���W�'�] �a�캙u�z}���O��8��M�]��l�>oOZFm̺;dc�]:Zd4`r�S�)jB���g?�̻I����O�5'
2��\e+�fd@^\�Z�Q{)F�3�m��<!���6TD��Cq�p�T��p͵֡�@�c#-҅ai�`J���Y���͞�3$�C����"J�AL��-��%��"���3���ɋ���y��δ��F���s��ǋ�� �6r:����[m}Y#��V�DːOݐ��&�;���H�}��m����+��X�ʹ��D�u�9U��`��3J۬{��BT�?�6�:�Oꆴz�/nM��>�׻!\�}��Ƀ�b�Dc'l��S�VJ����o����MB�,_֝�/M%n���uY.8�mt�<F�ƀ�}	��������_�Ҫ�;��(�NR@����$�&��/��E�	���3,�&&V^�>]t ߍ�^��y����R3�ŬJm`���nW2�^�(?[dk��9C���ЍBv^ʄH%���q�۩��@E����P6n��~彤k��k�m|̫�����}W�oR���u-���[pH4���;�9��J1�J����qs�音" �W60_�x| �8[���_Ĭ�#?�TBʆ{_�MD����֐�s��m<f��l���e��<&���+_�D?�v�v��E���5G�9�ꌰٱХ�������L���݀0����ԺM��⽛O�.sW޾!���A��f
�0)蟆8Ŋ��n��j5�Ì����a�5��=X��k0	�ښ��!�D�h���ܕ��`�!ۻ9�=:
�M��>����84��M{o%;���x��Dz��M_3`��c�%�M3���RG����˲`��h5d:�����������B�u9Wn�(��Z�� ����8�OX2�QA���0�תq��1��7��\�o�`��������]HZ��,G�u�}���bM�Ddw0�e,MF�X5�t�ع�6<��~.���7PA7���8�e^n9����%�?,v,(ԏ"Q2��O��q0K�s2�P$��SԺ�nl��Ia6�Ҿ�f�������f�	q�s�����C�bT׼n���6�SS�s��>%�K����
u��AEMX�ї���������+buӫF����Y%��m��bf��>O����V���Ax�p~A ���D�ⶓ�u��p�kh�"1���hχ�m;�*��j}G\;1��g���p�v_��X:���{��c��{j�Y�ha���^w���l�	H����M�Qо���%	=��@WV�;�������{�h��P�(��M<t�SM�U�^F-��Ҥ^�hxpL�����o��MkE�m�W� �m�U�.��/�'��7Sk*zF��I54M�J�p�hp���@�^�M�7m �Sm{�����UK�9�X,�Q�D�'*��@pP�W~U�C��~I!�J��d;���w�!��&� ʅMϛ�*��B����%3{\�%N�뵲{��e����Ξ��:.��-��&DX�yG`A�A=���6�*L�!����_�B⍠ʦ�UZ!��ߦ~|�\ei|W��UO� �r�lC:�K5�=п�U+-R�Z�������'d%�=��rD��7�O�<�E�q������\A(����gp����ST
� p�m�E��7K@/���$|s3����,�1]z/KYB;#�at����-%,o:�7��;��wأ�{
��'��1S!�;��h)"� ��Z�t�]8��?ኽ�j����!ؐ�s<<��@��&�fU�N��4bgW�!8my��HlX��>�x�e8��
4���������ێ�v0H�V�HoJ�j[�<?'��0t�7qR��d2���~0���C�;|���M�=��Po��ڶ$z�8�.�"�T��R	}��?g���F��en��&��@�|��D88�]ؚ;lV� ;�[1�JX@���D�j#�����L�j��3J�9�x1=}B�� H_y������K`^�RqY;7��\g�ӖdL��{��me���n-!�E�Q�����F��X���uߺV:�������6�A �7�Mۈ�7vG=�Ȟo����hI4�C>�/��pKIƈ�S5V�A�R���YFK�O�'�5╙BaHɼq�ED��5�	޿����E�%��)mu�!�r~�cZ�Z�!F�yo������]����᪱�u�o�9soojQ[��x�%w�%��o��uG�BB5o����:M|�r"���4���fk/:�F�bsFE����v��Ls�9�W���ґ�e���0�B1$�:Q���x"�w�Zq>�]��)�ގH�E�S�ؔ��L���N1c_	��\c���Yy� �	;,��ftDg�c���<"�@[�!N����,>�����1w�N��Z�N�*�WI�PƩ�Ǜ�܏��킓����ci��u�J��R��66��f���DѠ��U^�ʨ��!$�㴽ZFH���D���ꆎ�)���ۃ]�Ci�IV
�)�"f6��o>�ըd��b�f��}����.��L�θgϯ�?i��%fgJ �\k$��b^����ݞ	�u�vJ�PK
5!��[!��h|��W�z]������z�bgzхwƈ�f	��=� I��I��aYӊ�B�~)�o�����!m��U7�xs����Q���,D�̬x��Q�X��k���=��:p�>v�]#��:��g��7�r�l�1��2�>����A��̤�2�uǆ�ɦ��t��W�q��bޤ<�&����U0�i5��wh���\��{��AG��Cs��Y&Xl���Lw�\�f�J�?j�-q�7�b��E��#ș��%�9���1��n��H:i�+6rb���3�2��S�%yס�Orr��m�Dg��aҐ�"�ր�� 5~sp����fq3���'-3D��H��9KVu�I��`ys�-��	Α���Pu�H۲����h�<���Kյi�/^A<������M��;~����i�Bڇ�:}���+e��;U8%��o �\�,,]Q����e0n�"�T�r*��G�E�1`grZ;N�ж�#,�mr��z&yw�yO��Bm�NZ�w[�A?k��E�$�:_2|-!����x��8�#B7v��Dvb6i�]�r���v����j��ϒ��� �&u(܆պ����Z���(H�W�(�q>h?Ȝ�����(�9�ѹ�3��A��XY���vP��&ܨ��A
Q.�k�ڋ������*_�	ir�V�}V?�**4+�$�¸�Z�ʓ�5�F�%�l��bZ����ݏhGs24��ÖOŎ�=#�=�]Xǭ���m���y7G���y|�:$<1"�ʳL����y*��z[{%����r�<h߶$�Ǽ^�KZ�S��ϔ�Y���|D�"/�y���2�?��2����W{ɥ���E���t�"8,��A�Ϲv�0;��ap[�}3�1�mƩc����W�$�%X�y	x�����bdI�{L׷�M,�&�?|5�E(�d�?��]���^�&�9E?_4�LͅLB�8�9;��둼���%$PT���Z|���L\u��RRz���)7�e���+�J���T�'��{]�j�Ƣ+��PF���5�Y�k$I�jY� �vʸ[�����'��c�%�BP*���7Pm��n���(��@��j���J�?�9�4��lyK����H�r�MO2*��
"���*>ޞ
�&B��Ѿ,)�Ƞ��54�>�q�n�g��:7a���� ��Kpʮq���(��+����0��y��͹�|E�$z�V����lB�����6�v'���O ��LAd%4�p̿��<�N�B��jQ!M�[A�w���"��	c#k��c�&:j/W� :��u������?I�x`��@2�Xe��;d4!#`�o�O�+'5��c��9�v�?�4�$�j���'U��8L�\�<���Ot-�Me)�pe��?#NV�O��Ŗ��&�L&F�n�t�(	��ۯl3����C�|�O�4a-bU�(\�1�luAr�W�#`� �Fr]�VwZw��ȥ��ܧ�;�̧X�/̒@���v�p��C"/G
x����w�Y�D�脼t��^Y�B{�����VmLx�(#���-P���05��y�AS�!%x0��X~�u,�z��2�r2Y�Z�7鷎�D`_�7sp�#Ι�Xn�G[̴��9���GA�uG
�eK��N�b����ԩD���_�6vy����=_O����[�kOR7����q{Ǉ�=�!�@oK��"$�YĎg}O������f��:�$J�a+Hù�!��h|<��?���T=��kd�2ϩ���$o��зW���ۺ��`�m�����t��9�'�x|"�`�wO�=r k��|jT@s�JEv���d��l�&?]��`j����!��U��ۣE�C|0K���Y��o7-�Ea��Z*�e�'a����-P u��AoP8�bN�l���a�e���P-�l�a`����G7-g��������YC9����$�S<&�J��.Pѽ\,��l۝U-�/q�=T�u��w�*T��2R��h�+(��O;S�p�h�Wz��'p$�l����?�~mM��-�p�	Q?��ɳ���HP)�+�UzS� ˉ=x+�ϙ�/����6c�*�zQ|�$'���ɗH89>�#�ܧǵ�I�]]�NN��A��D�1���;V	~f(�����7"%B\�+&1(�e�˶3��vH��]�3��SLL�#���[�;�v� S9}�gA�����/�f`�rz��V�CV:�1�0O��B����T_��FG��Z�@Z�2E�g1R�B�E!14�Lf^(�����ɔ�G(��5��F�Fy3�k0�]�U:���
�)�TG ,�.��>�]?6q�1���z��$���B��#Y�c��&^Q��c��V�����%�y��u�L��U�z(�9,�4K[a���o�5ģ*��F�1�^�(�ќҵK�q J��t���%�U;ʮ��P?�,�9$Xq���5�ȝE*�	z˾�+�
���b�W�'���W�WB��̓P�!�b㛲�)�ϛ4BQ��I�E�)���,����%8CF/���,ʲMC_�����?-<��'��~VI��)ֈb��r"NI�u\M���;i%�R �:G���z^����n�`D�)p�|�����j�K՝FP��^�߯�v����-�=�(�&�hU��Zp�	>#� olud���Zl�'^���OP��4�'t�%t��T��&Mk<���3L�ɵGHϡ�;�uF�ɇ�a�Q�����dN-Xo��K*6�^��n�o����ڭ�y���a!M������F����]F1���)��Z��_9W3b�z%O�9W��h�X�<�|B���7�
��}��W��·�˜�r���޳rY����{�V	K�o{칧��K�J�4�p�e�����HOqqZ�:�,?/��L�~4�I���d J��c��Y�6���i1&��^�k�c+R������=��;?|�Ig� ~俸E+2��/��8)/�Be��������*�DV�j��j�A���̥���;�ו0 ��v_n��Vw�p�<tC����4_�������|�*�:��Sw�z������YH&�c�����r��x�9���D�.���e��k��1�����G�p����,��8+����LIu7:ݛg:�s� )�����[rXrSQ�+�#y�/{��6�� �qw���?�>P OO�����Ө�|�p����s	�,�\��Β'$PZ~ܞD��f�^�Gȷ���ˈ���2�."�	5?�X��H�c�4������L��b� /w0�Dop��.b�
@��+I2^��"�x��Ѵ�8N�_m�3���*c�Y�ˤ�3�z��$tS�>�
k��-�&0�l��#.�&����竀��Jڒ��v���\���2[�Yn���WF:h��V0d.��9y��ՌҼz����b�`��}��`n���з�lh9Jȷ��]G��W,a����-�Cj�N�O�Ի�3��D3�͊kP���]��qp�8���o���7�����@�)bОq�s�e�E^o�^�3q�e�%��˾�Egp��>�=� $-���d�㧈�_��W�40�!j�Ŷ���QE�0����"���W'�
���ߒ�*vvP��ă���i��0a�e�w�$7A(&Wk�Ly�g��}-�K#&�U�F��<l���]�{�U`�8�x5�~��.��v�|�v�A.��cS$��R�3BP[��RqŁR��ezޯV���������p���Bז�8�\gS�4/!ք�5Eh)��F��%e�������%�M�a��ǉIA�@b�����~O��L�m�	ZI�dq��eZ���zџ�!c|��#!̫��(l[��HT-黨Z6��'�tdz��uo����������*͢�S��	e`VU��\�^rC��?h>�5�ʖ#�H��U����p�����0k�5��Bqc���۶f�����'��c���%\���䥆w*J���9���0÷�w�ӷ���� ���	�-l3��� C��+���-(�^���@C�q���"��[C�9o%��~�-�ס�[�Gt�"������eA`�Ux���ޔRӉa{c�x��g���^Kw����=���z�k&�r�/d^s*�4l�W��(�1�b�����3ͅA��!�h�Dj�"���mv�
ٴ��@�wt
�bh_�����2��їlS��u�kzk�ZՀv��D2��w��9g1�@:��O"�o���Ny�S���[��:j��f�Ģ�yf'����VL��$�T:Wf�[N����cW��+����JB�3_t�d�CC�r���֭�� �s��.h�o��mZzc�B)s�Z�mG��u�hb�Wm���o���o����$���c���z�)sų��k).@W�ۤ�����qm�XO�{S6���[�0�&�����5��b�7�'J��D��5+R��Չu1K��t3_Nx(�$H��r�T�A
B�I3/h���)� ��11'YsO��'���
GXS��K��F�?n��d���I�k)�I��aZ�����y -��&�.L�pN����֒,��U[��_`���]oґ�P�*Y�o��鳺�+��Q���pg�St�ʑ��Ԫ��J6����U;/g�$<|�.���Nxóɸ![A|~�g�lW�wz<���a���o9�����^�DDL$|m���z+eT�sq*�-T�okl��ܹ^-�,kG*�����gia(j�u(g3�!Q_�[��i�����u�����aC��G��x�{xO��#���C	�����6< "��I��������v����o�z�~J|GF>� I�pQ�	��~��*��m�Ӹ����љ��y�mER��4����������[-�=@�������CB:KM��_P ��'Y�L�r�h+�� j�d�u���ٓ�Q����,_O@���(��C�a�WP߸d��C��~C�����?�Any���7K��P�<
ڨ_[�Z0����v�։�;B���m®�P]�{������� ��?~�l�ykT%=�F2���ł�	筞6�H��ڟ��=֐En�W\Œ�L����J�3_��y&Y��՛� >��<0b��Y��#l�eL������'���M����y�5zv�/�qbMk�,݇��[�k�����n�!t3�B9�n�m3����g�
O	��(��qv�G���,]}��r���G'�n���DUh�R�W&Kwv�;P��X��n,�� ���"�G��c5��35������/���u彤	x�ա�-��f-;筼��M��E�%K�x�3\<�0m��7�c�1�u.-]'87+�L�#��?S$zk`�ϙ�	̆$���&�E'�� :\�Y���ݙx���P��H�S��t��T���:wٞ�$�r�xBى�Ɨ�WJZ���
��\2`��F�lS�;��~��R�3�g6�i��w�Z�����e�#@���8�'~0�8��[�N�n!�E_[�.��x��ۊ�j�#�p �	��hxZ�[�c =��t�3/�w�������=O)%h�Zu���q8���
u|�1ëSkă��f�������{Y9�K�hh�_��qk��yU��;�M�h4=:��B$%�;���G ;`EvYD�]���ؠh�e�i�1�1�sC��?��©�7 �g��Xx6�>�Z���F%
�K�#R��BH�����+rMi��p�'f�Q�<zQ��J^h���Bm:�A�Ɏw2z�:���͏���X�[�I���+I�.���}Jl� )/�˿��O����F��H+����=�3?���Sm����'N7�,E�%f��g�(�j�3LB{v���ꬍ��%�� 2�`D��j���7��R����́��kYF�p޷C4�n�o��z��+�yLb�^6�N���cr���6 �r۝"���U�^B��J���D$վ�w3*3�������Dt%� ��Q��3����lƬ6~���t����Q��%�u��Z���\��SqL��S4���$�Mny���炄n�hރr����Rc(�ԃ]����*�l�:��w?:v�%�ޱ�n�����r�+��&΀͒^�}����}���"fr�m��0פ�\G�v�������Z-�JlepiՁ	輸�
�4Z��S�I8�vH"9R����i�¡�yZ]�G$;DȖ���Ǵ�\��ӾS�ʆy����s�S��cW5eRs?�{99'�h�l^m���j������5��):��Bq����H@��.N��A4�v��i�E]�2�0�$��kp�XIx�ɺ'�ݽv�����'����6Ѹ�5�N�.��K�vY !�U��t�i)Sz����V�ܭ�к4���L,ZtFՙ��*�k
�B��	G�Ɯ���\Cc���@�R������u>�D̜6�!����Ø`x�r6�71b.�"��/szv!�4��y�J^@r�a����S�L��#Ι_�K� �_�5j�Lbp��k�j�+���O0. ��oEA�z�t@.A~>���R��+������M�ܰ�����t9���
�����^n�8n#g�)e-y����8���.>�E숼ǌL����k).���`m�63<�q��gsu/����$l8��D˦v<��I�p����3|S۪M�,��0f �_Ck22#:�@���%Hv���oǸ���,J;�P�XEU�R(��]3��R�����$y��G�tK|�B�Q`�%>^>�0&�׌�C��K���H�t��z(���m�N�v��q�)���~����xOJ�T-����
�k4�;"��"������al�>��vP�� �B-C>CM��}��S��Ӊ���u,U/e�3��~�7X�m&�G\��y�.�U*,E������a�~$��aa��2*�w��+������ }�e����<I�2u��{df��G΃΄H�&���@��M��ѻ1�є��4���@Gz^YA8�9N�g{��"rؙ}$�vd�(n�~��6 湱��	�0���^��NxE�q��\*�����mǺ��G|�"4�;������g #�<��hk~��l0[�HL�L��Lz��j1�0�z�#<p����3��M��9�d���U<-F�%U��v
d�5"�+�@��m6�l��F/��"+��I�R<��f��>�^�xX�O5t}�M.]�6`�[9�Sm`	��.�|����a
SWl��!�Փ\��o����I��;�a��¥�W�����?}���GH��!k$�?��ܺV�L�B)����O;��<oH��
��\����r�ԭ?�5^�|�Ԣ��� ��l�D�Rhw��T��b�n��O�Z�G��|��z+	�V��'��3M@��2���ÀKu�i��a�OH�5m�י"8�#h���� �iY�4P/�vnn�r�l	5[���`��E7(\(k�H�x�S�+q*/�U]�JK���QZ[�x�y�w��Xe8GL�����#� ( �W,_#�0Z7�����]��q���3[�!dCf@@��E�a� r4�A*9VM�.�&��C^��S��(��e��j5q�F>`\a�S��f8�[`<t��4���Y��w����f���A�=��ʸ�VW�OJ`\��&�H�f=��Dcd6f&�\:�b��>��\;>�w��K�4���j�C�]R��'���h��t�-����"�J�>���,P�ÁA��i�jF.�|&������^Yv1O�&��̾�I��%i�GN��j�ט��;�1һs)�[��	ah��TC�|0���mX�v�L`9��I��:���7Nb����@a]I��s2"���\��AI>���[~EmU�M� ���L��΍�[��^�|���
����c��W���T�j�ȝ�Be�KfnF�5�7���˟"�X�ƚcf�H��)�K;��n(�m!2�=q�5�ڊ5G�B����d].
݈6.�����g�s�8�1[��F
jp��D]\��ڱ��`��W1��vA�u	�Mpj�1�R@:\ԃ޲Sm�&3r,u��q�M���v���:Z�tM��`}q�����x�F����}��9��C}�ac�6:�6��­;c��@so{�_�:@�ɽ��Ou
�
J�4��ԟ.��/.bTC�	Ifqzg�1�5*�D��K~�H~���Vl�WʂFNi��o����ӵ��{��p̆b*�%F�2s���BZY�<��0�9��U|\��ܲ@�iG�����O�����I�4=�-��a)�1�S�`��pI��NN�Y��	;�d�'�9^+o�eg�)���3k )3<�׉���zt �1�x��HZ���k:/����Ջ
j�9�\Gk������sDu�+Hz�,���ާ�/�1�P�H��xQ|���>��lD�oȵ��O �Ao�������	�"�좵�3[_G��	
��>u	�^���[M��W�s�@�"$A��m����!�U$p�.�����&��pA�Ll���,e��e?�h�������M�@	�ap�r�\~��M��͓�d�WR��g�����	e��Q�B
���Q5��L�(�ӓD��`(>��Z{�����`*�? 5P��ypn
�>��(����>1�������R�\�
�*b�6TA������D�?IQ�aEO��|�]�&�\qAZ[�.���׾�[�)0V[��W��F$Ȫ�a+�� 2t��pO�]qǐ ��~s�@^��a��"�Laöx?��R=��|-PT������Z��e�Nn�2冶F�",r�e�&�n��+�fW��t�Q��v��d�cN@���q=s����!�L4�%���s�󶛲s= ��/ܻ\�s9��9-��w6��O��i��E6;[���6�c�n?2-$$4��Mb@$ě�a �]��:PAd����oi��#�=�Ƥڜu�sT��*,�)K��\��C!1y�>�im�~R��X�G5$.E:�j���)D8f��#���4��������ޘ�
s��t��{B� I(
���۩;̺a-R��|FE���j����7*����׌�g�ߣkhyw�6��n��m���Ò�:ҭH�V.jŖ�V�7���t�#:n�g1�UR��;o���'Rcl�����[����&g�d��-�*39��'��:ΰ6B+b՜<�����!�ˡ�֕[����DnY�?.��s�F�Yùu��,���Vy�ힱ!Gҥ/E.���*;�?�G��K�<i�L�hl_��yj�0�f�$wn�G�)u��r�h���]&�����M�ZHE�7:	�Ժ^o-G�M#&IoD���_� ��O�qh�h+Q�ioZ�0.�y�h඘)P�
�C�g����l
�u(m���H���ZYHm�Ys�`��00�{�JjĒ�x�H@[���"��`�N�Q���z?.1�~����)��0<�-7�%@S;ޙ΀ʛ|A\���>k���r� �+��!�u�[��#"F��L��:S�qk�L�✽���o⮇y/�nL`��t�g�������
k��:>�dSN�I��������d ��sJ~�We�'�:@9A������u`u�5|��M��q���iw���c�֡?�j�J�;�08Ჽ>�l��7�x��!&k͟�X_����K,$�!���&�#����:ƺ�_�f�	�;�;���ߛLy3Î����b+H�&�x�Jyy��$J��?�A�S���������G�3�1���O��ޠ�FO}��i���oȈ<��dJ�7$i�дˠ9L�ͫ P�Pn!Neq7$i��6���xcl�	���׏|�����8|���M�~d�v��|��/�ѱ����n��������I>Wܺ[����^D:?�5�B|fL�-@��th�]���@�v��H*`p����������: �A������b����@@��\� ,�m�f��.�s���t�8��b��3���x9�h��]��#+6%S�ml`�娙�+�TZ*�'��9 ��lv"�t���O�on��zg��W���-���ղ�YFtuƴ��S�X/	1A�1���m�W>�)ļX*��J�آlo0�����@�3A�Ԟ��Ů����[�nο8��g���W@O~ ����/�Wr#���ۉ�v�.���-��7u$sE����� ��e�����Z�H�&Ԇ�UN���V��er���/�7����l-&2���%�c�3.��<�A�`R��!�/�ק�`��r������Q���W8E�h���ΑS�|2�n�,�����W7����'6�W^Ug�_�J�K�p���b^�;%�眳��xO��tk�fu�l޽�љ�|
r�MJ߇՛#i���n�
��2����	j F�$��SV&��&-"n�M�5?ܺd�G/�RLǘ_'�,�f	�싖����e)ݞtm7?{
l.�D�[��0o"����J���K˖�B�)�B�����{�� R���a���Q)ʼ�����4X�2��
ˋu�a����L�(���T��aK,��� ���k:k��Xj��,�Iӧ�5���\9ɢr����*����?�|>GvN̜nHQ���}�@�\�c�Z��;�"��D̍���q��5����vB�-m������Ro�="�3�Tݔ���&���Mb�IE����S�qmd�#�o�����X����i>�d�SV)3n�},����7Q���_��'�JW�r)x[��=�Q��F�C��7=JE�w��WŅ`3�!� �\"��/T��g�ˁ1\�h�"�2pҘ����2���,���f���ⲪY�=�� �v�;��]��O�c�D~�K�O�����$	���d��$���٫��G��BQT�}�-���n�U7�Md�y���K�ʯ/Wä��<�̄��|��򴁐`�O3��D����F0�4�z�Fn�yC=�-`x���tpUR;��T�߅Tb&��a�� �2,�,�N�8�;zU�!��.���m��vw��'��5���۾@�)��96��dȣ��_�i��X%��|%�hE�;�B�R����:����t<�����������4-���A	��ݐc�;�=pҦ���}��ʵ띴�!��A0;H�0O��ލS8�2��F=S��F�wNt�q�5�h�5�;��RG�7?J�ȱ�`�^sᩎ=�G�c[̓N=N^o����e���F���z=)u��<��	�Pȓ��@�+��o��
l@r'?��"�jG�dG!]�]b��
?��p�������Τ����)I/���e�| x��϶$\� �!�ظ�H���cK�m:9,q֤ƊlTc����g�@й��д:�eøii��+�w��e�ƙ���|l����D�L�M���{�mOU�`���^T�a�I�)��������M��jW?��Dr���)q���Ć��G���P�_�>p����VU�e��/�8�V0|�Fvhu�5��h�z���<y,�G�V����7Kت��g�fz(��o��4:g]�̳&ZI�}}���b�A��)$��rA��@i�1�ml��"X�YU�\Ǹ�m�E��	nVRM��
�J>)�6-�$�0a)y|Ca8t�� ���aMO�t%�ؼ�g8�t�����c6���I4�B���-6�{"��0E��R���5�o��B�؈}����
'-�����*{�7�4�}��$aq ������ڤr�g��X�)�Ό]��~H�F�-�	Ba ��<O�A��u5k ���9�����i��õ�<j�>�(y�𧃝�&�Do��D\�T7"�M�E�ZsGl�H��&�<P���R������3/�vb-m�rCJ�Ŧ�COi��w�F
�H�����-�4�C�"W<5�O���^��N���.�����ta��oM^7��t]�P���T ��G���s�
�q�KnbU�U�g��']��ۊ(��Y�L��B�{k�m�`��muS���d0n�p����g�����w��>��N�,ܬ�-sOZ�)�'6� ������d��!I��ސŔ�D3����S��3B�D����k['n���\Y���s]w릾qvJ��頕^z2�_>P���:��9�W��+���� �#��c�U��5#0?U15k��Ey����sl�5�`CR��؂#+툞Sħ�EV����#D��w��z�skJ >��Fܰc��|Tߺ��C�VY"�s��"���8b g�y�3mϽf�h[��I{�آ|(T��x1��T�	���*3��C&N.,[�H?q�G�X�:�8���SR)�$]B��Ne�Y�SO�	-�l��گ�8H�^�KZ�Dxǀ(�ȯV�	*l���3f�N��[��n��?�|;�Lwi�L�X����|�\�r.q�bA'��t��"5w��&T�`Ÿ��ԋ�q�6$�l`����~�wT���z�kݞvo.�Z���bV�c��{�Hh@+kc4��TZrOs'���lQ�)��G7���z���+���E�zQm�\>�T�/��<q����p��8�-��݅ʙ�KQ&B��O���*r��N[��B��R�� B�6S�Tw�)�y�ڙ-�'z��Kh�oxV���l�� ��.́��Up�8�ެWxf�3 ���0�./Җ��Bj��wy���tO)�2�Y��P����mi` b�F���ZJ�# �-�ؿ����inH6���# �ѸZ�T�:�)���a#�/t��m�V���4���&�H5��q'7�&��Z�4L��5P�x����8�L��@R2�v3a���2Ӓ%N}ōq�H�HT�K*nIЃJ���G�U�zg�3K;�5�߆+���ݠ�A�v&��]�Bd��.NMj�ƩP
�?A�()�~e��
h�T(`�"#~tp�C�b�	���)%��A=u9��3c�Y�q^�o$؟G���B�L�f�E�䈲�|�䮨���t����ɽv瀄�;��QexlZ�II�:2X.�c��7?�p�d(Q-m)���M/�cCg(:��d�~z?�$kvѭ��J����َP����@�#hN_}
�|O�'�b��D�%��!����f�г|H���d��F��u�#��0�m�i\0��A�W̃���E=^�y�O�2 �������'�m�zZ��i&H$ ��G[?�#���T9Q� ��sTn$!W�����'ܫOph�;���T�.Mo��šL�V7n�h�(f���!��bߠ��$X���Q�B��;�����6s���8���p��ٷ�o��xHv�!���m��%I�%�_%'
�ޘ@��{�0$�&'Eٍ�02y=W�Nl*2J�Md1J/���>��i�L���W/�6� ;�ƵG���i�5"�<�2�i��}lՎ�q���u���2�0/����.�e��M��:�yv$��B�#AT0��_�����k�AƗB��>38$�&��7]MQ�ָ~?rOג�O�d��>�(��|�Cs�VH��@����(�<���CxCl���0��[��������1� ��兂�<�j�s�h��9�d��i=u��b���/�=6i:^SA�������i��L��z���V�݄&L�9$Q$º��g��ʄl �0��k^"{v����b�(G
��4E*��$�1Y�Y���Cq3$w=ͪ�a�\�{�r�U�'����ƕ|&JO�t�]Z��l@��+�>�u�<(xn��W�G7/o�o(��	��y+���ke���T��"v:�V�8�g68�;�|��.+�`V�񐑼O���|��0��Z`��+V��J�R��ON�@���l��� 
x���,孔��
`�k���]}����Ƃ`�)���"}�2/j���sg�T�@����<� ܠ�8�"g�X{'���}��w)*,u��i+O����D=��~� n�!o�%�#����㠩��ޓC�b��F������>ׅVo�L(@4Ƣ~��6�HK�Ԯ ���������~:J�f� �"�evN|��qƮ��'~�N"y�����c~��l+����ߋL�nXPl<�Ւ�c����|��^ih��e���dR8���M_F�� Gə{H�r�0����`�iH`*d����oց�ܔxϲ�$��v�{����'��KE��.<g4h����	P�(2:��q��¼�A�*isq��h��>I����e���Or��l&�$��l��,�ύxt������^z$�~h��a�r��A�9�;J�s-P
0-w�'-cWd�C��,��Z��M������q#Նd�8��@L5E64<�i����*:��糨+R��.m�U���z�x����X��S�V�P� F�� 4O��5��<*4U�r�ϲL�!��q����<ε�_étB��p=]�}jl�Ev~�z�	a��uؽ�Kt㈊�dD�z �Sp��t n��B`<vO��8Ԙ�M�,]6��yc��O����W��������Bl�H%c>dꗁ-%�F�FO��\b�O)H�*<��_�� E���Ku1�<X�H7y[B�-�(��v��h��iY�.����+��!]|XQ
{��eo�H-D�(�����["G�a��ճЍ��x��2�Jr��P��@z)�!�¥\z�����x�-�F�}Z�]w�⒪xJ��1v�i�j %�SZ������f<��뚋��a��~�*�:�Fa��M�5���Z�����[/ö�j:uj��>����E -}�5���u�����ܢ�,+25U��0R��ixX�:��s�C ������=���ȧAmIC�/v}vA���7��xi@Q�i,_e ����a��V�H�=�w�_� f����w����44?߄�-��e���y?{�Lv�S]iGߜ\��=�zg�D���CNף�k!"s���~��A���[5����F�}��
S(&D5jK�92�=�Bs�a�қk�(fV��Ŵ��q�=�o��t59RGn�ԧ\~��Ϲ�p\�������~�� ��d�ث�Sl��ba�+)r�IB�����VC�-*�HT��я�VWP�i�mڎ���AD� ����R'��w'��AC�S��=id�d������C��2�ِ��	��_,�Ź��
!���}�H�5�V�'�թ^Y�ߓ�=-�^��*����N7�>7�H�.ᔿ2���o�Z���=��|#��E���nnq`�(lo�-ˍW�.�3�9��"��E��r���:o��c E7��9*� �C�o'����0GJ(��݄@�c��7�҂��LTv�	�Y���@�8 ��dŏ|��҅�\	�J_iHm�t]��r�"a�,�Z:Rj^����溂��¹cq#�Fp�x?5[#���;
�RA\˺�+�ʼ����;lgxZ�Ic%����X ��dVC�!Cj�u�&8]B��JV�	�\0�.\�:��
,�d�~{*F�h�%t#̈́��Wm��VJ@SMmR�S�����GfF
�:F���B	]���Nж��d�x�\(����!�a���{��pc��u�� �DЈ`y�S���3G4ŇNN��TY�tӤM�
W��1'�z��t!�HmN=��s���A���F�/'5
�aI|���}WSǭ�%�F�7M� �7į:�s$�@�sߣ�k�r�$�~G�
�f�9@g���:f�����>�ֺ�B��F�吂els'��K�T� ��Q��ތi�;�3�Ĝ/Zkg5��~1���;��ԉ�5�ۋX4�}#��w����f��웕�3��`eP?,ښ�c�,�΢�X���]���;_aF`��&?�����/A�D"��E�¥~�O|�ً�Q���N$������ŜQ� =3=m�y<�g��X�aG��b��Hׅo����t�
���33(�ߵ5���|��L%�w���+,��y��mG&hc�?f#����y;��4�p���ʱ�SmW(�;i��͇����:ύd�x@╍�<�w�	)��)+.���<]�D;�=�̍,:��>9uV�X���ٚ_����\��C�;�y'�P2���K���0o0v݀�KZ�,cR�SK-m$k(���ϮX������wb~Q�'��.���nr"�RY�I]�YNJ7ھ�ï@/�p'N!�L8�c�?V-+�{����5`}4��,��m�ؤ�`|����~�q���ӻ��E�Ny�,k|.iG1���B2�mv�<�*���1f��tskۻ$0U�E�b	���$��9�;�(^��ڡ)��
T`��<Ȍ�3|�a� �����W��\��lj��a�
���[��(oY�?�uįR{���_p�?�)�-^L׊������
p�:����XM7�V�I���öx��B<��N]�X��Ií�$�ɩ����5�$f
r���R�7���@Ш�uf6���?	��e�:�K����\�s2�B�pdɗ,#��J�Z�&���	���<v��(U�����3 +L"��b��Ad'����upͧz^���_m$ĉNI&�2�I��{��Z22��n�x�����FX��"M���:^G�cv���� �X�P&�E��� o��H�@?r�jI��=@tC��P��a(�W��#3�`O���H��=s��,Y1xy���ڰe���8��}�hV��$��몎�)� �D�!%��u�®=��$�������z*��%E�VhG�8`�Dzq�3V�iH��*\!�K���n�䀝V�僇9��l�[��K{��6�'`��C���w2��PP�l�&��~�Z3t��H�1�5M�l8JJ#���R[�)8rH�^�������3�O �SX=�o]�nU� `���AF�yv����N���M�L�[N��o�V���s�Ҁa$�씥h~6�'#�&���f������<[!�/y��PHǗG��%�^�\�D~8�mja���S��\�M�`�[��#0$C N� ��o��#�b������%9����-m���B`̒6e��գP��&sm�����u�-mSZzi�SC���{���^r����|۵�,xm2�k�u=-2B�%^"t<z�<�ΰ���k�L�A�]B{�R*�p��1�E�lo�+q⨱�:6w-�	~��M.�}� �,.�a�:pT�c�fl��dOH��\�?
�LSB�	 �_�����:�nG�5jO�8t�P��0ҳs*��1E�e����e̴�éi[��I���&�� ����M��φ�P)��}�I���f���\��}�oJ�O|���B����-]Y�r�XFt
�u#@��Ȟ0g���ו=����B�:sIxп��F ���Gʋh�����1��~��2�EcV��|�)0�w!H}���{p��'�m׈>x�#L�SC!�E���'|�x����~���hu���4-(%��.�J�0-�����"bCг]C#k0	�GJA{�%<�I\��-oJ�,��Gn �YS���R���]��{[~���I�@�`;K�P���]��9�W��'u�	�\��|t&��?���x��|��OתAD, ��Z��md�=�E�j�Nk�=r�z�ZP�N8��}AԹ���G��O'�1d�W3'��]���d�-B����KMv=�a�+�AK�aL�M���둽�jt7� �ܮ��BQ�bo}�m����w�$1L:i�޻��!&����2@��wK^�O��U�����w�^�e��2^����v0g��ܒʈb*gc�>���!��U�o�2�N)w��9P�ыX���I�/X���;%X��&�Ph�[ۂ`Ʈ�)����K:�+�Vto�N z_���Y�d ��˴A�T����j��؁�,��]-�V�b����{�afߑ�!�q1����)�R���Sؐ\Td>��K���T]+�~�W؊e?ܸ�����uf�ķ��)sn	 R���1��=N�˂�O�)�'X	yA�q	HSȧ���w
�G���贽]�G��/�!��M�`�j�=��8C��g,��S�2IT)�a��LL��C4"Lm��6l=�xXA�́�2l25<t���v����C��d1`���R���S�%mFJ7�g��#-���p}M3ԍ �
�J>2����r<Ǌ��I{e�{b8I��C2�B����b1��5��-�=M8������)�5)m�Rd�ccd��,��á�9��� w���
f(�f��"�;j�C�e��'z5���_��mk��U������$�$tt��0<��v^�U�8w��*{�Or"�7�w@/ղ���(TT��5o[���:E�j\�߃f+�c�1�.�Y$��cO�m�E��X�{�ʭ@iG~N5iUE�-�5&�/�w��*d$/bC
�[�OAP.����X��	��DU
��a�_����U�6��[3��]�t��6Θ�l�۪:�F:�F��>�x�K��qE*��+��\������S��?����%�9�~v��I�ݴ׷��E=��l�N�KZ��wS��t�W���[�{E�C=�,�̰^K����޽�I�sP���V�9�,L<��~:��!py�U>��؀��9Y��E�(c/(ou"�VSVD�s�._;胝��,��9�͟�Z�U^m��B{�_e���e�\���ߎ�;�E<4t
o�7F�!�ݕ~�}DӓE(�×�>� M#�T.��^��,�'�MQ!��[P�A1�e��]��҃vB��PLA�D���G�,"��~va���%(��,�#�W�)8�	��ok$iŸ(S�2̘���S����pD[�:u�>����+^���YA�؟��t���v������Uz��r���RZ�]RIDI);����_�Mgt�ΪG.v������eg��y/Z���7^2rI�xռɃ����Y�	��:��_^4�̭H�+�A힮�l�tƹD���-L��E��E�I ̧��.�q2\�����OCo�x��Y��p�d2ķ��E�Y�Fv#�$2)Ǫ�V^�腼Ť�9>���qz	�Ef���%~D��M���Pb��d��_����=�� �J���Z�-�N���RO4V���Z�.�V.$����Et׸c���6��OS>)�`b�vr��z�s�a��[���v��Q����}g��!��`�Z�;��3��c^ �M�D�2�79�X���Z��Hn5]�ȝXDe�Qu_i}$ph
;+��`eZb��yM�~�A|�펹��O FT�?�U���Q/�jEs��:��E�<G����mS�&�J�U�����?�l����Z'���Rq?��S����D��c�e>��f*#)j�d�0$
U�S��ޛ�fD�sG�m0{�iV�n�H�P��R�X��r{��(�s����Zp �gLU�O�U��ˮj;�{5��X���ԇf��X������N@���,��i�w�h�I�1b�୍�o�'FHd�"A�������9��'�����_A��Mɤ�G�h�b�f�̲�z�G�zmIM������cRH?����K���h=��dz�yEjqO=i�R��[�ceW5��!�N�Hg�W-��DP<���a��Ѭ�co�y
����b��j�Sw��k,�7(8�:�ҋi�bg�	�z��d7��$�e��{�f��.̺�#p�l{��ȋ:ɟ��Ŭ���ga�F�7־?����Z/&�������K�`M�6����S�m��Ԣ	���xX������q�ف���Ȉ�l�����>��Y��A�[���0Έ�V�H����a�cn�wNė��/W��7[f�z��V�.Ņ��,|P,�i�F!��=J��cN����b�xP���j�m��E�i�ۣA���KXZ^�]��7�`��fs��������S"i��TO[7���[��o����]�$B�㨩��-r��U9��W2�,	Vr��ǵ�����2j�e<Z�^<z�=���1��<,x�6B^KB�况�=��K�D;��l��"��x���g��?�>(*�В��t�JA�:��L�̯��O��I8y��P����w���$� ���G���g�yz��偨:aBúh��6$i.a�\�{ƾ�q'W1n��=�ԣ�TX^c���'������t����%�Y�O�^I��y42�� *�ל�	<6�a���K�:9y4��E��A�1�)i��cGt���c�֣�]���B�5��{i%���t�KR�9}iy��ӛ�a�sM)�9,E��I��}�KU|�i��{!`����v,:�O���H��~$�|�㯤�z4��d��4*���G���%�/�>�������x�(?��O�-�� ]|�'�xMC�1܉Úm��/�w�4e5�.��ni<��uu����B�;��tP���U����JπO�( ��u�p�YW�|r��6��檬�\Gz2�R"����M����Z`Mk}�ʹV��mp�.��:�-@5�R\fg�5�hՐ&��T�	�,��1��o�7���A�E$�沏�����5��+��Ə�@%�=���cH�eD�]�-%��ϳ���z�����p��HR�v�9�P��S:|�c�f��������B����~fkJ�����l�.s	"��n�f0�~��{�ݠ�N3?�k�M5=��׫ɋ7u������r.P!,�v1�H���i�Y�T	����b�Z�/�)��qL�Ȭ::�%pZ�w�p�fr�%]����%n8����ʽHi����R�h�=�ەr�?݉#O)G���X�--6��D� ������'���-N}xȵ� C��/���i�@@����6�퍎+jb��Dx��hCT+��L�?ߪiFP>���N^��`S�I^ݣPX^�O�P�s�<ެjњ�B3��:'�\��Iq�Q�Ј	�0T��!ł){K���]�]G��{v*|,wT��еߩl��\�@�F@�(?����H
^��r�b:E8s��u��_#�_�n]8&�mkŬ�e��cj��q���ּ��xh:����3���(oR�m�d�Y'�K��Ь���2����llO�[W��"�u���D�K���^�U����PLNz�nɮ=)sm��	%����D��|�I��e��	�n�����Jz�N�.|�OkQ�����Rxh؁��r(��l�a���k��S��H����'��3-�=��f��P��g�<���:�ݧ�y�D���F��/� �x�uVy��vQ�ko�;R#���� ˁ:la������YXj5/	����xIʙ��PF=r	�?�S%Yh�q#Y}-_Z�� �ҫ�s���?@�8�M�#���k�m�cȡ�x|�;����H�C�d	�{�CN�Ax�}���7�Gqa�5�r�ӷ��H�A�@X��\Ob�M91_�i�2-�v�Q`B�a���kM"����������Wp��<��_��ZjNgg{���H䑆�+�q,(�o�F�� �d*�-�w�H�����(����\��_=<�Pt�P��&]�����m�H��Zr
�KIh��(�V�g��Sx�I�~E��ޗ�Kڎ����f�ӛR�B`@ϑ�R���^�Vf�ͮ�^$]y�-��#>��\'���?w�
+����NI��b�%gO�4���>�*C�~�"�=d���pf������IJ�
�7�Ry2ؾd<�l-�k�_�0"|�B��|�XP��j���?���ٶ��Yi"���ك75��v�b�|?d��4�B������m9]��S$�q����Q48�G|�*'�$�q����[�4�_��� ��&^s[�c�Y-x��6l�t�P��/���3jN�ZY(6	ڍ�V�L0?QN���,����P�ٞ;E/V�l��[�Zqk).�Ev�	�
:,�#'w#��r��/�-���{�^*��x���*���k�&�N�@�Rt�S�}�c}��F�a��rit|�OT[���[�N��������I�%������A"B5Te��+Ξ� ��ͨ�
��2���>zpN��3�❔�J�����p�{��x�a���W�K�ue�Ԩs�X؊����q`@�%t�6���I������?6��N�y�1�G+ =(&�R �k�ȌQ�B}R#,�\�G�����k
Ĕ��L�f`��>Z3Zf�WYm����v���$���z_u�)��{>�p�b���{���v�&�O��^�ȅ�S�v��P�� &v�f�m��� zScɺ���\�t���-e��	��;=�J�\N�B�Ј�i���C�V��j��ϖ�����x.�
+��5!fVE��?$�Ge#�ᇿ�$O_F�kYͼ �WzP����=����6�L(��5�G��`�N�W�۳4-���7tm�u�b��@�A,{.M���f�7�s�L��7�z,2�OFQj��G%��Fi�b]����1��#*~2�6�4�7�Jդ�����z�fv��^���p����Opn���Y� UN�=��~�8��7d-�	F�8Q%�m,��������h5�H��pNZ���]�aٓ<Tn7E��S��1��tu���~y��z�4��kᘯg�.�^5���q����K�����DM���W��#in�0���1��6�:"�n���1�-����!���,�Ct�Y���x������S��`�,�L�K<5+;�wM&5� �B.�����:�A��������P�;1y�D7O�5҈OG&>�v�k�^9<�$g�G�c��2n��y��g��lZq�	U��s�N�|�-&�E#�D$�e"����i{��YZ��莔Y
����h��LY�Z�Rd�2��a&ϑn��bT%��EW��4�|�
���� ��F�oZ�f��FyL����(���j����Lw��WQj�C!c��!c/q;v��V�w�Y[g���_��.��0��1��G���nc%y�45�R������{��/S�����y�È.����cI]L`c�ׁr2m�ȌԵ4wֺ������Gaza��M�?_]~�� �e%��-�F_�$K"۫��B��0���!����0xt���u2l�I���2�_5g��h�,^�~��y/Qc��}Y}g,<��H������u��'������}-36�/��B�]�F��@��
d#Ux\g.�tGB)��UМKoE�SM�)b��lY���x �H��@
<I����̉�/IE.�,�=��X�c�&��������aB��z�i��v##RZl�[Ua0ؔ�!��Iso��$���1Z�j�@G�k�Wie=̶}�����D�Ph�����,ŧ	8
7�%�����	��]��9d#TXks(m��1G>���ˀ��{�~A�4���M�X�D��P�]a2�Ƒ�qnk垽�3�5s�|�^GH�����,������GG+��B�B�f�s˼�I#���bOy�V�}�:_o�]Nk@�2���H����A�x�������'����!'�֜Y�hr��&'}ߒ���aӔ�d:�Wnmi�x~S��F��OT{wg|� �+�O�8����ɐ9���8���0"��(�c'T��FI�-}(�dt��)#,/1�A������s�W�n$�X���H%���߹�/e�F�QzR���N���n7����v�
s0�J��}�xG��Q+��ω�4�B�Fg�A u�ˋ2��N+F �~�R�R~_�*=zJ[*^��Yqs���y��s�U��i�Z1�(R�)ߝwVԡb��c��D�X�� $��G2%�TF3���5>����y��4�V��9�kl���qG��Z}�φX���IȔN��VB3�����ϐMƨ��Lޡ)�4�% F����n�[ۆ��T��@c5�+@6.���ƣf{�U.�2j�{�pOf�0�r�ۀ��;.���mHh�m�s�sY�ގ�~�)*x��L��4dr�n�~�r�K:C.F�Z�K�ܿ�	����}Z�T�/_"��^�
�Zh��ǉ'��JI\#H)�rs:��}����V L�i#�^�.w�vz�{,�[�J=>K���)���EL�n!�cU.������$-��bԠ�V�`�ͩ.�D��EN�v��˞8� �E�F	3/��V;��c�K��
�*<�G�]�C\.�� \��)��-���$&�����su�_[��/b�F9�~3��V!�L��]�,�g,듫�#J}U�[�j�?��G�G��Ic���N�\QG�vV�?Ü���n���	�%@Kz�xqs'��n���5�O.yC4���U�79Fi������W,�v����:{Wn�V����TB� �6(����˱ �N�!n��� L��ot�}]���n�;�����4Ȓ�t���� 3 �)��х��"��fe�N*���OOB�ev	R*�<�YN���/��"ۖ.-)��0�R�D@Ü��Lb>9r[An���������c#���Yŗ�S�/�����xm�*�g7���r��E
�5 -*�t�;ڍ��+ڴ:Z�j�H��N<JHo�������j��,m-�*��5)Y;�GrY� ��ց'�I�y:p~���Y�zX�i� �u����r���b��,��|�p��|��ĦV����~J���h	ءA��Lc��{�-S�O�@m;9ay�ʀP?�^��ZNi��|E,K���ŭ�,��I�D��� _o�[6O�:Bf�ߏ�tɆ�Fn&�\=���!t�ׯ.������.�y]H��u�&x��*�B��D)U�r�J����
|�(���F���h�U�"�9sS�\�0�4�l�42��k��3�@P�:��F/��#����k"�h��L��Ti��U�׍��G��_��$�Fq\�vd=kNX�m'��vu0�*��N�Ɋ�G;�zE{�w_���)--IBɼ�i�R�g}bĨ����XNc��#�0�Ƨ�ܰo+�N�Հw�5'ub��تU��O3?5Vg����4nz8sۭoP�Z�
�Uh�U�ִ����7�P�v$'L-���L��n�y'���Ix��	�tN����������ڬPA�����W��Y}c�4:������
k�8�_�}TvީWo";�/�<�P�|������:~\x���}�_�.��'�f�ܔb����#��W�M�~�޵�QZ�q^)	�ܳ	t`w��9�u�r*���	ω�d7S�ĊD�g7�}���j�����K+Y�Ƽ�{4��]�D�O鱭]b<�N�H@��	��������p�c�$#3�;8���o0cV���n����b��MT5���vQc��p�w���y�#�Ş��?��@w������2�KT���]_$J ���y>P+��~�c�o�D�~Ő,HV��|�"����b����}o�G�� !)�N譔~3�rk��:�;�u�eTw����>���5Ɉ�G�/���ZR��� ��Za�S���𮟶��2:��ӈ�����4�f�v̛B/F����*��t�;�� �	˨���fs����|�J�1���	�_���sǯ��#j(�t�ZF��,�:���NEz�lƛU��Y�'�-��e�-6�dՍ�M�C�d �y�R?�2�Q��,�7 �� @V�Q_%Օ�=���п ��0��w�-�A�WϊX�v2��@x��D��߁k��2ҁk#$}���$&F���q# �>`��m���7'���9��b>��W�C9Ý�=�)Y��°q��s��P���ì��I��A������c���o>��͞�5�l��Qݰg36lPE��gh��~S�ï:��4�h����#��{)�Ø���� x���'G�<$�b�����������8��Jn��KHbn*���B��r�f���G;p'Q{��aӇO���m�>i����h�����S���o>2,)������n�}\��M��+�U�	�	b쟒Fq��U�9���/�uB��?wrx�"u��_��S�hB�EE�7R�����b����f���?�;�/;���#6w��T�0�K�HE����7F�Y�}%��n^�5��]��Ta}:��h� ��Ev�]��Լ`�P���0s�.�ט��O�P! K�kOdV!b�=��_`�A>֦,s?y�_]��M&�e��ͬ���p�Q��s(*���]a�"��qԪ��>%���*���ER1@�
��P���*ҝ���Ϊ�E�8���;:�	��69	Ac�D�b�+�t?�q��"�ĩ���$4�)��Ѹ�t0�vZzfb{.>s+����\��VV��1���-���68��TB�۹E�@+!,�d�݋#�Zvø"���z��<�0�
�M���G0!2�yl��pm����������;�Zwm�d�s>�����-��)���l=lW\B�#�$	�/-���d����se&a���g�t��M(C�t�@�1ޓ}0�-[6�ط�$��H���>z{����ͺ�~��	8�=Hu�[����i��d` ���FQ���Ck�/�(4�k�Y��k%������C@*��P�O��!9A@�,�F!�ST��ٽ{?=����Ó�p�"ڍ��J�y[9�\\s߃�*Z�g�y ��Z:V�}�?�E1c]1�p�d��(���1%i�!A@1\9�^1C�v^�
YeRt���Rۜi�:0\Z�7��.��V�Uu;��h�e ٜ�i˼� sO�$?��Y������4v��=��$;� ���A��Y
�rc+�΍&���ȴ�S��˷�[[��V�d܋C�Y&�����y��n2Sd��Y����ۅ[��8����$�]�������#�oF�ig����ɚ���z$�b�d���5р�����>�Q����@2t��YnV$PV��-�o��v����%������~�:^�~�O/����%5��ᐪ��8���p�V!����3�lA_�~8����I���f�0��	I�ĖČ�(�"��㑘Y�ݡ�j����d[���#�X�Ռ�$�o����S�i���g�$����ɹY[A���I?vT�?��O`�����|�+�P_��^�ؑ~*��uX�����_T�7�e[�sQ�ˈA�Q��PZ�K��0�y�3L���e�s�����/%ϑ�1�/�1F�o ��f���'���[�qh����b�Ǿ^�uV�G'��3h�r}7G�XJ��1m��]H�A�]ctfjM-��6i(�e�-9�D��X�|�3��^0��5;&�i��"��������Yc#��i���)�]6��Mo�j7��&��&��b\Z�,� �9�9=>R�$p����e@��`������V�Jv|�D�z���OW�e��R�3|�y�P���l�+ �`b���knMF��h���n��$��>���A�O	&۽'߬w<Ʊ^���y��3�6����:�,�'�m��ik��X���p�Z9,B����%�Z�<�rNpS����@�浊�$�� y�eq{Q�j�ਫ਼,	��cl����<�Ą`ۄop4dA�j?����-��B:�Q����'F�A�%��sn�+�M*r.0l�$�'�O�hNFdEG>ŀ�޲Uvu�x�׀@(�dgΝ+�CG�������Mt���m�
m�ք2��P��
�cS0�ʥ���2��_Ӏ�`EdD�@UИ��N ��&�Sy���0BT?��)8��[��8����tz�ڸ޲_��(�"
�&��d���WR�3�� Q1t�Dv[�h6p�卭@��?w;�I4� ��*Ĩ{=�8�V��u�� H���u�CH�����,P�!{9�I�Lh<�[���@f���
�J�rn���&���C���`%U5���)t��z?p���/����fm�I����	RZ4(��0i&�-�߬�r[M��}�Z�(���G4����S�����#4z�<�<C����جN��%嫱�gI��oa�ɍ �&��*{f^��'?�HER%r��o>�)1�p�hZ�?����Xɟ~J"C[�v���"�ʛ���]sKM���.{����w[�%`4A+.Iڗ:�-7
P�)���Q�䨮	H��e��߄B��>He�UDnf�r�Ưm��n-�����϶�Is�o~r�>I�F���G��t
	��&ـ/<�*���{�ɗn�-'��ۉPNn�ʐK�ģ�D��G��y@M�b��m�5#yut`#t��4�ݾ���`�<���t8S��gǠá������b�:��1/�Y���O���(3��j�Z���yo:W&�(�|t��O�X����Y��x?����`&��S��#��)�M���5.���ܥ3@A����W���:�$��3ρx�j�R�������:Vb=ʗt�$&7o'p|�
|'M��`�$��(�($N(��P�^����z`5n;3�s�HK�1���/���WǉfH�H�$v9x�O�$Џ�L��W��q^$��i�6&
w�ϐ����B�;9q�_Bo�7/i���E�X�����q=�Ր�<Z��"ԷS�焼	LtbD���oDחݜ_�o����篦�Z:���Fli�HҊ����_�p��e)���3UZ��b�S��{%,��~�z��,,J�(K�r���ʓ�����Fɹf��!-6�.��\�g�V%B���N���`�R:�����$��2�{k	���$&�aٸ��\�ǉ��f ���9�w;� �_����5�k���̏��k�g9x/t]���ʥüi�T���z`=�D$�*7�Y��j?�9
I�D��A�)����,�MpB!K)��];Z��N�����Z9-�"���Jtr�׺��y�0x�b܍犺]�j���Dt�߮6WJ���*	a܄��[���ov-���	��
1��2�ȸ}���)0��_
��/��-n�e(: :.|w��%`��y��ҒQ�&ۀ��#l����v�Q�2�rX� �_ڍY�{5��?�QuN�I9wFc���_�J�6)��W��zr�L#NQ(���>��� �����\�����ވ΂b����>7ǧI���=��YxQ���}�/d�r�sm�1�Xp-�1�˃V�����b�'OY����`�j|��	���ݕ�-ߚ��v\��,�i/�#�G�,��:����CB�ց������/��1')���Bf��M�)�m�q",~l l�W_��n�]�p}5�[���������^ײA�S8���=Bf�@j�}�jW��i2�J�uA�G�:��H���Vxd	-Ḍ�ý�2[�\�s2W3�IC(��G�2tD��IF �L�U��������ȃ�q���T� pȚ�Ly��T����Tq4���4W,[�7y��劵�ĖZ��h�>�8a��D���I��b~SI�*����iUh:�3��S2��S�p���~vuo�2���伿Ȥ<9�3�}�";M����\���e?_�f�J��.G�y�ɔNm���	T�*���H�x|��)>Za���N�[$�(�=�g�cn��'��JR#��o�.�R�m�c^��B�/H��q��΃�Kx�+����Ǭ�������5I0&PU#���,	K����fӢ�14sW��5���frRfr���RR.4�3���b�ªr�<�Rm�qD|�>c�xp��<������9|�S1�Ѻ��W���!M>2]���@�〉j��Sm_�xm����`��\�5����<r�-ޘ��n�Q�eQ;�d�Y]�Q���^�-�
p�K��`-�Qی��NJ�S>>\�͑@*z+"!*r�h��;aVr��$��r���sX�L����O����?�ze���]~�3������N�8��,m�)�#ҽ�'��ޙ>�U��#rq+A矈!&��9��m��З@�sډ
ʧ	b�mV?�Q�?�|�q���r8m�����m٥��􀵁J?`L=" �?�$�wGN��=�UvU�^2ŗ&$*,�(NE���%B��g��Ib�FB(��%�,=�Q�����悩�����9�C(F�u���o��ۍ	�m�%a���}UJ!32k�F-��\W�+��v1��Z�o_u���`��[Ky8�n��͗%Q���'}M>g6[5��l1��i�<e� ֩8b}HВ�~��ŷ���,�T:��E���Ő�\
��~B���߰$R�:��k��=4w��Ud
lzm<R���5�ȼ�_ף�~,��k�׵uW�!T4FX�a�T��.����D����,�������V��=����4cP���I��v0ɦ��7����(�0����+��f*��RtJ��I6��o�W\!�dY4ʯO#/���2VT㲥�<����u��gc���Lyog���ק c�?�� e�`�l�=X�h����am����},�3�	�9��%�Oɥg�-�xu@�_؋�,?W��7��36��f=-7m�}nR���.�Z�Z�-(Pl|~'y���p�����l'L��g(����)��R��^�v����˶��u7�W#�\���"8^L��c%��r��R�p-kȐ��R���=��뒂��O��4e�����/ �eȍST���y>f�?@�s�m`�W�$�A:����a�����.'�m!`}]a��x���\�.�T\i*��Y��� `�(��gc�9������z�2D�C\�X>�=%����`$=��UP^�Ϯ�\K����e5r�(�H;��|����Ç�J�c���ԁ�u���gm�tʕqt�ኂ5!I�Jom	C�K����c�m�*��y���*�8�϶-`"nZpڏ��)�&Ѵ/tw�y���]#��+���;����P�x�/�>��B�E��Ip�%���Wukh���ɗ[<)�c&��C�F�]�5�i@�<��mL�ʵQ��tX��@>uQ��n���z�8�������Ѓ�֙9�OL��F��~z��
8����}�tѰ׶`D: PN|��0�À5���mws�9)�{���ɸ�3�I�2���#�|1m�&���G!@��~�#���:�C��/쮃��)y�pR��Д�3J��
�V�`�)�,�eׄ:�ޞ]B�晪����v��K����]�ע2� �Yь�M�4N��r 	��4o�V���8 $��I�ABy*�=��{'�4����M���ɔ j�//Hm����A��`,���L\�``ޭj?��0�g��"ɢ�DgY9:�l�OI�(a��������zyʫ��k�zo�"a�K�F��y�V��|���E)L'6kD�,��N�f��c��V�w$��r�;�˚�ci39��m��`���g�o�4F�(N�Y腙�A{R�Z��٨���{�y)CB�	���O�?_5������?��]��p�r�x����e�n�ؒ�pLf�Y[0�f�ؼ�0�bxuw�����x@�#���S�y�tC��-�+
�`3H�z�e�P,b�1�r��QT f�5�&t��7I%��o�Ac��S���{K��`�����[5'��^���I�m�İG]?W
�_"��5��P� ��\��ep{8���s˝���E[�V2;ϳ�Z�6�ڌ忨5#�������S���;:�p��|�*���5j�\* �{����=%�RCm����!����H��F�{��V��A2�B,'yB�ϡ_R=h���"|�ϛ=�)��#[B�V襻4�v�mLyt�CE�׼"��\4�/O���*��`�*����!~���Ņs�:5��=z&=���5�NMޛ�|]�sm�W���W����c淍nL��̢^���0�>���ѡ\������$xN�q�8ٓ�gZ�q%:�st��Εq]Ҁ7
=!����Z]s0eH�'�ǃ�L�W�py�
�-}�R��u\��&�c��?d��Ym~K��a3���e<+���<���o�Ɲ�,�]�?��(��;@��ܾ�f>kj���GC���	���K p@�ͅ�@'�[%�W������
���=���/��2�JK��T96�8�x��"��0��l[ጅ�L��q��|ڗ"�
��{�P������7yJⵐu�S�	Η�Tqe�sN�@d����%:c�Y��G����A��Aم��+�J�b'���S��/vI��, ]�h^����A�����z�&HR*54��=�H�;�ͯ��)�e�/U�?0DN����fb������7W,�m.����)i�>��(���6���'�M̶4� �,���&4�2���Ƃ��P�� |�wh�E�z��w���!)��ظ E�B=6�Heq,���)�c�m����S�b5.�k-���A��U$e�9G��A:�!v�i�S��y��8����-w� ��$m����̇d���?����d�3v锣��>��~WI$j���P(���0�xq^����N:_�}�����S(���Q�*����l�t}V�o�s��z���K�k�#�F��$[�؛漂����G��J�}{�[�B�;���SQ�|a��A�R�E�J����W�_����	����	!�����c(����QV�P�Fj�7t7~�.ҝ�e�Ne���^� �Q����e�>(�ݣ�/>	�:~>E����}�%`�}eg���n��kq%�՘�I�f��3������f�w���ۺ�*��j:p��+�,�U��Җ{�Q���Ց�����+͕����!��,��ܹrm6�ܘ������YY�������mİ�#�V��U�����^���9I��w���图$��I��ur�	^.t�d&�j}�cV��4�f�f��!)�wOS-�Q߃o��W����v��I���U[��5���I\��܎��j�o��N�f4.ҟ��Q(1M�&��a:wj}�cu��Y̞ {Y��:��'6��`I(fN�)n�EX��h��:���ൾ���-z.Kˊ.)��T꒖�RX��Fa�Ԝ��]��P;���)�������#�
�Ys�~�8��,"v+��(ݻ��].�ܸ9�x�l$������%L��v�	���Eo�0�+9"(1���򊾅	T뭢h�1a����M2�\UP�E��ζ�&���*�����|S�}� ��ɋ��}c�3&��l,��]�gE�׾���@9��=$���Y�֤M�MS�:%Ѕ5�Y��J������$<����t�g��X<����
2?��\���l�C��v@9�j���t������&H]nA%���b�籀d3օ�[�����#�HZBK���SI'zV�^|�Ŕ%�����_�pt��Ү��� p�/.V���%�DbL\V�h<O��B�t�2w���H��߁��K�9�CN�-^GE�2�;̓� Rv�%<$��a.'f]v�L�ڹ�'b]+�t�U�a���I21B����v�<�P���?XᲔa��@�r�I5�F���s4g��G�ZŠk�v�c�I0N��Ѵ�Ղkg8 ��^������m F�0)PI	Q&NW�~2�^	��-*i�![�_�g�h8���펞G!�Z���ǫ��	�&�������4����IZ��?�NUP���zL��g��AuK�����R�?U�6S��~�x�������0eU�ր���/_�qpmn��\E�i�,��NC��^���e���D��I}0;3��+��<�&�4��ğ~*ɴ�⍕�_�,�EՇt*�si�Qx{�蘎p������.�������j'�8 Z")�ǻ&��3�O����a�Y����)
�]C�����Cq��K`u*qؤ�&.�*R!#k����-'⑆�����2J�]����9��ѰV7	.t�&cԉ����t��~Ѱ�Y�bPG?P�s������8�,�z[x����*����M1C��1̔�]���̾�-f�#�E���3�� ��=0�QQ/\d���:�^�}� �lr��?; ��F��@�����T�B���:o��/WR��T�&���Sl와w`�:=�gsX:���n��)���TR÷0\c�餳:j,�Ӥl�DyL�$��m�aV���s����-���"�ʑ��a�š�9���z�cU�R�CD�b�p�־���5��lGQ�_n�hx�~_�SJ��7G��*�R�:*�V95>�h�_�8ƥ�8Arc+2�rk�
�3���>�w�Ѐ��n�J��H�$b	��N�(�=B2���}����D�qF`�%ھL�?�G9��8#�^^\:�L�o�a�,J�C��%��3��N%��:��Orn����2�/=�u�D����T�H��}c�]yr����W������QQ/������-�iKUK���߽�=/�)V��h`'�l� �rLΙWAޕ�� I��:�M��`�L�1�����n&�,�[
`���t�nk���l�LwN�{���YE�0�x��m��^���ٟ�\~�\�vA[$�����$
)�b��zy�8F ��M<v��U�N|?�����pt�yY�7������'��a(|�e���&:Bq\��k_g��S�aq�/�5�	ǎ� ���w��,��&O��E���O�Ԫ'���Jl�ui.����b�5��'�����DXqW@�؂㏬�N<�([�Ɗ]!cO\���?�ݖ���J�cF%�>ru����\�MM݃X�T���}���4�z�x槄��+�v:���e�<��x��I8g�ㅓp��Q0�s2�t�\��	��3H? ��)�G��Y=Ɠ�[�]W1��}�M�]a8_߱c�g��!�u���q��A���>���Vx��doԛU�7�E�*�V�b�·OOX�����5]�|�r��ί�5Ҧ=��T�g���N�<`K�&��˱Ì�IH��Y�����7HI�hx�GCR�
��rXD�(T����0�����R<H������Fk	�Nh"JO��Ύ��C�ـI��3��;��ۻ'βB�PC͘���WXLm1��]v�å��F%W������=�T�s��.��_R2-%�8�z�.�@Za�fO�>ٷ#gw�hI��h��S��7��t�w�L�I��%���\���K��5,�~VJ^�â@)���;�$Y|�D���D�ӝ6R~�6��cds��ă˶bVn�8����I��ش2.v���_S�)R����X��M%��ݤJ�"s�#�m!��iL7CSsw����t����L�vy4�x���~zA%Ġ�ǤF7��m������&��[r���D����^z}MxM���l�P�i�˔`�7e�Y�肉$�)�mz�6�-"�l�u�bbP
6b��}�z+��F����g1�H���[���t���r��i��[g׬�s�Ž��e`�q;��#���mT�~���PNu��Ԙ�ױ��knN;M�Q��\E�2NvF�ʚs���9����m��~�w�|��e�0����6��E�~?�}��6�FXE��U�^a�j�bC9�=q��)����Y&0�F/[�.J�?�)"`�
Q��������)a�>!�wU`�����P��p���~�`�5�z����5�y�dbXӐ�Y�j>2�=~��N%��X�=�+'�Η�l�N�;��ШI�)��C��h%�M">�6�h?�L�����]B���v��o����i��\l�Z�>�ߋ��1����Y��k5��h�]H�1	Я�o����*FEQ�a�Rϥ��L*�v���U��-/�HE��E�u��:�����a�>]&��h$ԱjTJ�x 7eV�ܿډ!5��v�޿�U[U��gHM��A̰��M���i��S#vmf��+`�M=?���@A�]mp��XЋJ�{>dx�k���߽�i��֘�Y�ҩ:��8��/��.OV�M����"�UF�)
/.q��~	�z�/�K�v��^n�J[���Evo:��$1���+sW�u�A�9X�G��ډ�M���e�D/W���	%����c��ʷ���b{F�"Aj|ͩ$�k�q=+=���O�����R��<#գi���$W�\�e����������<16�i�?�{��B�ҹ��u��@��� 7�S�����
=3�5�`��b�� 	ŪTz#�j:_��ㆇ��� .��.+9JQ�5xu���r�6��I�~ǉ�R�l��1{��\��)1nl���3�
dU}�vu�I�5�5�w�iI|t��j68����u98-�x���{�D)�p�?�kt�X�s߆�������f'����i�@����6��#�*����j��~��ЉI���28g���$I��[T`��"����2�*y3�J/��Sn�Z��6��7ڻ�K��pO/����<� ��v#��hPk4G'�Դ�2So��y{+��K�W�V�:y�UF�1��%�N�H�C��i��)ܖT�<�npDe�Á7?1�sW���V~���[�W�v�J�����'M��O��v��e��+B�2�Kk��D+�/9~�ʭ?�w/��b�p�,�޿�;�be��%Z������>���f�\�h ��F	e��=XT�d)Uu�Rx�mQ�	X�]�q���2�ũ�Y�C�x��,��:WIҁ�Y`a ����F��gAxe��XO�`�>�m�
�:7^f��r�6BE\L5	�/{^M�������D ��Hh.�������`;���$5�����wTa���O���E��z#��~�GY�
2n9B ��z%���K�^:�BZ�3�/U�ԾSԯy��b(��"A�>�@���n�%s�p�T��⦐���/��L+���$_9e5c���4���֑j����~F�q۰�I�:F�%<�7&�e�b~���	�W|�A�uc��U<�����V��+f������Y"w�T���߰����9V�����W$s���>d��D]D!*a�-f�v�gb��&G�3���8�����#����lf�e��DдH̎��,~W�[A4|R�toR	�ݖ�]��M�X�A����'���-�e����X�#��.�m��L��V����x��{��ӷ{F�6��zuc>���{�e|�@��� �M0M	�� }[8 k��u�<�'�����KYų-�a�:J��=qn{z�f�6 ![}��i�^�]��j� ��)����%�qA�Z��濓q������:���b�4$�T	��� .̥A��1Q�����8^���z����!L$.�?�^g�`1;L�я�`I����^����P�J�Y0����G��1a�q�H�l��,~1��] 4�!.o��qN�2��ﯻ��Z��Hhąz�%�]���xi+��t�I(FHF%c�����3���39��G��*�V�v�����%�!��NJ�	H��.��ƞ��I����Y���fY6A��؇pk�:\�/�25N��z̊���G!��Xǝ-���lN2�b��kp;mߝ���F��	������S&��a�Io��E��ʰ/��C<�'�����i3�+�E��a=�}��E%(�DM�)��
�2�d4 �db�ך5�j{�a��hot��&�\�#�x���;rx����^j�S��d�1۷֦So~m[,���KIg,�?q$��8v�ga� �Afg�U[��J(���IТ��	�g*z&����ж�*�o�7%.aǹy᝸Lֻ��<[�l�1p6����L��	_������U�\+��?]C��l���BM�cM��X�t�x>.ȭM��Q����\��.]?f��h@�S��@�i��Ry�w*�Kox�o�D6��&�S��,��+�����A�\MQ��E���w�PPʫ�P��n�[.�=�
�Y�Z�ғ+���!B�����q��"�b��cH�3\Ws�4�"o�K�9="CzOh�A�ziС����V���"�+ʹ��A'���5ߒ��1N-���/�T��Z�|��:�����z�Vh8q��F�)�-�R��#E�ˣ�>����ڢ���O+�����$�饆�b���th5��h4h#�H�A��."�j���R>�3W�ݭ�1P�F����R ���õsX�ьD�愲�ؕc��yC���}1 ��_���WAXж�|�=p��r�}7<�$�}�3#��0�3�'��b��]Qv2zC����e��1$ﹿp��^+Q��t�x��S�H��?����<9H��]��*�Mo�Z��IE�':|������lƵlI!f�bqՠ����
N$Q������Mv`������N)��,[�(o����a�Ȅ�Gn�wF�{�N�j4��4?����ѧˏg�y��h��o��'��V79g#���s��٘��d��u��6�	�s��u6~�r6L�C���&���_TQ(_Թ"�-��?��CK�.�}3x<�)]{�-��$ݥ��1��g��,$�=c����ŗl�@�d��r��cv0eՖlIʌ�V,��߬f�����]C�"B���..�!{�~*ɻ��21D�I�����b�ƍ�������,7�w��Z7⇚������f�W<�Af?�gVU:�.��ev�dF@����O
���\L��qܜ���ߑ8�%����������,�􃩹P�@'����fya`2��壱��Y}��T+�{��6�`������������y�$��$s�t���Xu�Ö�D����{�����K�jwI$�7�9)�
���J�f��Abj�4�5>#!}a�ۋ�t����^�� �8�3�������B�Uo!o���V]��Q��%���%�6T}����/���}s���9�ݔ�E�3shR=���7#��pa�(
6(�-�SɃ��W|�S*���L_;l��i�b�,Jz�����Q�����̋ۍ��V��
��܎%�_|<�����rM�b�2N/�T�R���X�*X�"~�H8��Z%P]D*!�a���^%���1�:����F�<X�[��4�*}{_��yT��'�4�/�%1�v���qFr ��[q�kp�^y�P0���6�C�F���T�rx͎�p:!��$栮��*,�W?X5�I�)�L"|���Hh�Ȃ3���\��Fy'�h�Ih`ɯT=&
�s\�fT��h��h�8�����V[ B�AB���۸@~Y�\U�2��(f�@�(�=)���s�#IsX�"^T���B��N<_E6D�m<1�UL��%M��Tc�{M��fS9�!e�����H�}�W�A��:�w1��n�7-;v�fB:~:�eXM��]���V�0����m{����iXRz!���@UKA"���AgN)s]���4o1���N� cg�L����db} T�j��)J�c��ob�ؙ�g0~�:zås6*u%��5��ܢ%�̋�s�K����0�ŷT�����L|wZ�~�4�N�����ﮨ�+�0� $!5�b��o<�˭�.���2��-j��e�����[� ���vo뀾t3X� Ok����:[���j�n�}"�l��cD���^�/�����`Z�|�L
9�ZB�M��}2!E��������TR��9_L^K[��2Cפ���!����C "D��O��Ȥ�����??��B!z�{��8�	i��G�jT�\+�<��H��A1[e���8yW3 4����&>�q�+�їD��=ՑD����Y�0�O'��~f�'��x��Α��/uLZ�lZ�yL��)��P��g��m)a�]Z�2<q�/���?%'s�O	..IX�y�笡�"
WX&�-�j�Y$�|�2t�$Y����Pm�t��F�O�(��	�~/`�����yߍ*-#�)
��$*�O8p�=��*/�]VG�5��l	��i)[����z�Y^&}Ve��uP6����(Y��e}�J��zT�Q�=���WG!����N�>Y�F#w��2v1Lj=�Z:�X_�Ā��QS$�x��,]e�+�1 �X���nKڮ�hq���su&���]����X�iG?�m2�Y�mə�Gc�?]��-F4�ӈ���r9�ߞ�(��]�G�B0��
?ɳM�6;�����-�#������rzG��Lgl;�/"�"1ΐC?��������Z�ϊ��V�-I\����)\^�7[���K26}����-qD�\��l42m!i����)�Wվ�,�����Y��E_�芿}��K0�C��ն��<�o�x,�O9���,D�� ��� �a�	[�X��7+�9}���qBQ�U�V�sՔ���\oɭ�F1\��ӆ>�_n��H&�5�`�y�c˲��9�}
�0�%{�v�*M�uw�M��_���� Ĝ�^�4�L�XEl�����ӬT�1/i|ç�W���q���8T���M`��:���KO�l;�3����[�@O�qYqn������K�X�eK���"Q�S�+x��m+�)b*�Zs��}Vhۀ"J�{�ݥ�=G1+�)����%j1�q7H�G��%�9'� ��"����n�0RR�.F�ֿ�ޛ&�P5��y�7��^�6�����m;	�t#@�I��f�����N)� ��̖�״����I�Nv��V\���	%�����-�Ί��.��H;��r6�+X�K�R�0;1���J�l��c]5�`k�YqP �y�
����&��Ϙ��ud��F���<��������"^�	��U�Z������U������+Ơ��F�9�4/;R����dҐ��So{,�}��]��/m�H���Y�_��,��E���M\�r��-���VQef�~�ج(��&]���=C^��,аk�{�������}a�j61�ϥ�	K��_�8N�d�59BK�,���@'?aθ���-@���р7��H�#I��?�Xa����<�����>�'�Cc�.^�gO_��NG��hff��9���,�3CS���hw�!�.M�C#�kS��k�?��Bt�����驸�`-��,z\g��y����~}� ����қ݁�c|w���D�dO�{���_�ӏ��ә�?KӑZO�rp���!R��Oy�,�
i%&�qE��#�wh� [����A�v�:���2�V� @�WO����gRd,(�!�۱(ہ��i _>iT���M�)p�~���魥/:��j���:�����P�e�)��Vl�dO*�nX��6s�-yG	�=�o�~#��t�����Y4s�����f�����
v���O1wQ��GƓ��d_�_�bG�ѫ�F�<�9!���H~9�(�ts�TШ1��]t���j�A����oG��ρ�A�����r0�{ � ��ᢑ�߯B)"����i�-6��]lB+�)w9�AI׍S��!���&�I����ޝŐ�eY2(���^����f� X)�\l) �7!�R�J�v�G�[;�1.9ּTW��s�E�>B���6��3-|� ��[nt��<���I��;އo�4l������&2t\?���R��/ρ�ޕ�{��qƢ�O=���k|�Dp����p������r�(+�F���2F��f"y��#�	w/�R�������6>d�<�*r$���ta\��E�N�TR/sff��@�]�^�l��x79�@����NA��̻����`�pL��I�3���,���r)�@
�՛e�lǍ#6J��8بl���*�����8�P	+#���|#����I�����Sr�`tro��;p5U�vh�2G멜 L��9\�PGr�� �,�e"0��3�HC�[�yUo{�-���v��N�Ub�����b��<f���I�Q�����������~�c�DR1��Q�.�g%�����d�>��m�^k������˧d`͆b�}�}ms"���C����C7��Z^PT�frC�|�xK�Y�ǳGO@���+�h�ev�Ͳ�O`��c�?r�6�+
�o5J;�dk֩(B9�*�
Y��!��Ds�h�9�n����.@�n���ꀛ��Y���md��s�U������66SկJES�����gd��ŉ4��T����U�n� ht�����rO�4�I�]2h?uk$��ȓZ��H��5���4�%rτ��Z�֧����� �� ' �T/��j���/K�N��^����1���뉣
@�)��@u��� ˁx������H ���� ��T����BN����g��?0�����0K�n�gM9�K�wb�;��ƿ���"p1\HNY�B��gEl����0���t]W���w�����oCM�0]�o��J��hy���!�
��G1�B�9|˧�&Vdp��l����`"��_���p�Α�ޱ@���#��=H�~au������ z��_�� o\Q�ݢaQ�F9I�!��L�E������nI�6.��K� Q��2�_?���q-����^B�C*��G���D���@�����w�O��V��|�f��CQ��ڜ�D�0�ŵ����M��F<r�'��gvg_O����t�R��6�K�'|�`(kzdeҏ�K�N�����!+݆�����~&�8���^2T��l����ޮ><��$��d�a�-�E3��]#�#�L&� 
��w �`�^��xM"�S_���N�9��G;��n�ʀz�!�o���yXpØ
��>��Xt���3�
�zP�e��</N�����/�?Rk�U�S���c�J�#/��Λ+�F*}*���/˥Π0���S�S��p%i����<� �k�k��#f�z��]8ۮ��f��f(�5_���e�2�V���N*:���4�Ӎ~+-E�p�)}o)�C^�=�@r�k@
�?'t6����I�ų�D��sH<�k`�>3�0|V�o���6��o�8���3���-+��X���&L��p��A�)[n�bq�F�hO�N?OA���8rRy�j#���J�i�d���P7{��R�4k��`#�O��ꏚ#
qAY��),4?p7��N�]SV
&b�	{~'�C?���ֿ��K�nb�tD�g��T������5���a���)E�'���" ��L�m�1f���0��B̽�Z��}���fV͗[ʥ�U5,�ʓ���t]Ǎ�[�l���*)�����lJ��oo�WO��;2����KsJ�֜�������V0�c»��Tz���"���6L��9��5tEB�������"�J.p�P7Ʈ��IaFj���wV"x[sR_�$�厍X%��y�A�jÝ���j�&�G<�^ezΣ� �����\N�%��p1�n��z�� 4�V/~x��Y�P6�]b�G��ܧ�P�<�#�i���A�`ձ�{�I�8z�I�b�ٸr��T�<��Nq��T��K�.�3b^�	As�v)1���BL0VZ�ni1,w�\0=���� O(�2���2$�s����/ւ��+�s�J-�K�`�jb���fXOs̾'-U�~��>h�1,�������ײ�7L�3��D��*�1%DH�D���{���:�P�՗��h�ȇ{�K~.�k����'��C;���&c>~=#��1��ߡ���t�T�Lo�����ϒlP{ﱊk�
)uQ����fR�t ��!����Y�|�:]E4v�������$Ќ7��š��Պ.?K�CLt^`��Å^lXMQ	[�0���bD>��
"0z2\��1�x�� ;1Fx#�	߯�m��Q�Ԓ٪���uJ��m����忛񁋽37���u*��������Ӆc�ƨ���we~���m�	��O�FҀh��"<ì�VsGgd]N�+�,��p*k@�8.X�_�yӿ�fCz�)m�Z}�G�բ�5�]n�DX�������b��]A02X 6fDXӰ�{�4���O�=]i$�z쀠1ɼ��C?@�S�����w��� n�B�i�	>��!�~*|�xͲ�1�{�B���Ĕ����/�F���a�NbʑV]�] k�*�r. bV\D�h!p�g�֋��_�P�58u�VH�<:>�9>T~�K�� ٲ����D�B���2CP#�����_�̒���=������8�z�s�PP<i�7�l�K#�(u�f=�J$T�q8=�+ʅS!���Ci.t��e#�%���[1���@��I�%.��.ix��� �/-VX�XA�W��#�eujo�&�� �Y�kv�Y��}e���C�7��\����Vɢϕ"@!X�-Q������yy�0�WDs��?���]�[��@0����}>�c�I�3�=��Ҡ�-�)|l��W�/8r�,Z��ܗX�k��*E}�������x
'p��=�L}��G�ݭ�'�m(&v�>x��P���%wӬ/��;�#Y����\{��[�1���S�����|�����mA	2�j�����Ο
5��~���׏H�6x��2�k� ��4�.jY7ú�AT6�N3Z�W)�f�V��?�N][��:E�����=�b�(��ބ�9=�Ω����o-~�� ��p�,���Q��wP?�F�@sR�+K��{ۀ��;�*��Ck.���Ȯ���>����Z[�f�-Y�y�����N�Ұ��yJ�����M�r6�d�8�Y^��ʇň��UkO��n�4#�~J�������hs�r+�lrY�����e�u+V�O�2��x%b���������j4�~/��/��v/�{Bx���+}ݙ��\�5���c<l�ej=��C �L�)�4��p��咘v.��h�j����$�gA��>��TA ��3�D�4Z@�y�폭~���j�9���� ������g�?#���4�r!	�_U4g@���۪ze$��f�{����Ŭ!b~;`�/8�hu�<ފ�7?�4W򣓕�+"�}!���%Z2�C�a��s�k��X��30 L�ݲ���T跞�z��G��r���Y
�hH8�;V��ESKЈ����Yu��'dԋ��nC[6�Xqq�~`����An�v>M	� ��d�GP��=z��k7���oz����8C�=��xD�����פ����7\gˉ��c��ؽ�I���(��H31�������\�&��9r�����!�b�9�UǕO�uPF��]�Y��8�ni�2��ɯ�:�d��r���6�ӓ�� R����с���Ve�Ǒ	�=koH�`��}=��S�Cq	K�yy��<��~��)�t����u�m}�pǏ�����>%o�ܦ��(^��2����W[1��>[���	$�$�:~ط�@ۊ ݴ����<��gEA�3��$ �.�k���.^7�'��,��&A]<Ĥ�Pu��Sش��&��&-^�m�ԕ��J/��x���|>9��h�F��^p�>3fàb��� .�"�� � 4�H�\
���.�榪����8I/��@c��������%�	X��[�֑�ĺ�s+Lٹ�4��A��N�	LK�N5^
h�h�A@�X������f�4��@_g �f~��A͡��F(�^�
��]}���Q�0(�L�[m�Z�s�;��9#j4�� X������TvY���z����4hՐ�
x��3��
�Y�:�f��ڳ�Swg=~��-(k;�d��_DBJ���[ߦ��*�u��1�B���e�M�'>X���$�-f�����_ǥ�~����vZ�g[:%�g�y\af
�3�=�S��*��Uv(���������n��E����0�hDJ\k(+�=ǁ�� �D ��~��|7ci�7����Q�d�P�y(_fg�]��h�Y���s-ݿ�IL�e.\|*[�V�aI9�m�b������-����_v�{�-t�'V��>kNA��<@0��*E*�$�/�c����n����y�µ?I�1��n����5���`����',݁�jL���<�ӥ����A:���mb���D���Mk[�7�.�V�Mq�y�n+4��S,;�w墯�>���}<;����.�b�1�GW�����1���D�]4�7f㌮>y��4��KiG4��b�' �]��-�{N��9����yz�z���� ��zf��XwsKؒ�ۺ) S��>5�Zq6�~?��e�]A�x�:P~DS��Al����s�}���"�"rF�PQq��G�f�ʆ�L�NjĽ�Ii�����
�j���H��EL	�$���L��1G��Y��4vG�d�ο����D�oL$��`dA���p;H��I�v��i��A�{���:�q�����<27LV�����Ow	CL��HE���AV�0���.�j3&�Q<��7��E��Y�JP�7�t~��Q���۩@�قӞ��K� �1�B����?���]��R[jΛ�-�����$;�om�j+J0j4i.E�����"V�-(�\l�*�eR��: �A���&}�	<����<Ԋ
��Fb����MzS��:@Б�4�2�3�u���ҟ�P��#W2���)��W�L��{��0.��V���4�܊��xYhH���7���&�T
��k�������d+�*���qXD!��9g1���PΖ��z-Ḯ"��;��e��$uڮ�1�0�k�EM��2�}��{X^��R�f�#._Mh�0_�x��la��(�t4/��>dK)�@��+d\8�-�kTp���F�/;��z�&��x�D��K[6ڽ��s���ά��^AF�<��W?J�5x���G'�������6k���ڼ�ԼH+]#����v�-��v�_�+�Gݍd֚���׬,��-+������@�.-M�Û";U�y�)Y�sy��
�M�<����mE���|���hUi��?�.m�i�=Gz���HXH|˦��j���a;Qj@%��~��x��&�䀔�m�`y�.�֌��w�.
��g�J�;��������Ɋ�.�v�YX:��d���g�2��[��h�~�Ո�8�B4��Q�����;�>��_1}ﲪ.$	ȑ����ț�1�2��ĉ�t\W��EJ6�d���ٟXܩ�ߍ����>@=Ԡ��t;d&ȋ��1���Ӟ�Sf�s�)�������d1Ϭ��jL
�co�siYz���5#�O��#c�����gX&4zCx�}��L���"������c}�+��v���M�أ�)�T��Q#�
o(ό&�/�\��ה8]}^�i�
У��a�bG���=�W5�{���iy�:��"H��@�z\g� ,ܰ�N�6���ēYt�q���8��~u�f���e!4�(�-ԧ�_� �y��0OgY�B��l�P�#���&���\�k_��G��SNl^1�Rn�(ť���n��<���?0)��X�F<K�6qj����2�����I�տOm�Hd��9��?�d3���c�Li�d�M�����[��`QX�at�4h�Ǹ2�2}.�?n����?�:y�����;���Kc���TaN飀�������W�1/($�(_��z <R!M���bOa������1��'s���+ֈGU�y.O̟:f����u74K!-=��g����7�wT��\o���o���N�*����-^�HlD�繷��:@>��归Y���R	}�����;$ˌG _	���i\�P�]I�)���1�(��1	�+hP��S�tz$$�s�}ZA��H	u6H[���x�y��f�Cs�5U|}�}o�����Ǳ����E�Hk΍/\��|�A7v�|��ͽXX*�Ӗ�YK�`�IF;yB�ҋ�� ���uin��B�H�V1�8P2��QQ����!OB��ߥi�pG�̈́�Vu23����o�)��6�fkh5�k"��H��s��ݝ��D�؋���QB|�E��������nD#�1�P3i2r׽���0u���8�M�n��ᴃƳy>ޤW�:�ʔY����ϡ߭=@��Y*eЦb*���.�0��3M$��%Y��<HN)�m��[R
��6$�.s�����%׋�ج��gq��+9�He��f��Y�c���-���B��h��rQ�f�P�S�7�}�&�ʧ����n�jY��9�#>��< >�S
�R��nu~����|Qt<{��G:AS�l2�b��:ؕ����W9�D}�a&I]
�� �Ã���Y��U�׹�!�Sv������U�%U��0E���Fe��}�ٺ��Qe!��)�9��AF9d�4�Km�?Y��4��=4�^Y <)�a�`/ξ�Fi�+��Ǭg�F��\^
��zj���(����ah`Ȥ��*L-�ظ��$�6S�F�@��:��j�Î�W�;��?Z�7b8���X����ʿn��{ c�ɻ�j�l=�� ����6R�T ����/��
ތM�k�r�46 ������ɠ��Lu�7ۉ��aƇ�K�������p��M60��ՠ��8ء����!�ʤC(^����i[P�r$V�ׯ�����������1l���ޮU�v��F5s����
�|����{��[�U�/,&�}�����8���K+�x����j�<�U���S��d���K��%�E��ޫ���0�$x���\)�|�g���}E�%�S�w5#�]�����#��aT�x� ��P&�cMo�$׹I�j�9����K(O���J�x�:+����kKlYH	�Eo
$��әZV2�h9D=��aB8i��o����I�mI懕����8Y��]��JX[�f�X�[��
�(�x�ѻ=S�e�v��Eo���@.<ť
��d�]��9�1k��vQ�����5-O���O�@�8�	� .Π�\T�v���h�/�J�n�и�r��{�y��`�ϕ�&Fc�k��I5�Q�cy|B�iS*�qɽZh���c�'�1�J��s�t/���O�#h�N��e������-��U$p3��E������PU4��} ��q��Ԟ殛M���m�հ<됣ԫ���m�P_��)K�+zB5��-�i��wv3Bx4�S��<�$p�C������H�7Z	����p�v��}�3�x�TV�{�L��L�7�[����N��	�e;!D�����~������W]�ԤaBX� �_�4��C?����ۍ��z�mE�cz1�}~B1��]%�TN��ƍ	�C���3��S�)���t�w�Y*��/��<�l���1�\��tLi�p�מfn���<����8�C���X��b�!��c���W���5VT:cK��]$Kyx��x���bD�L応��`f�M�����<F^�֤X2C	O�ށ����-�����_LYq�!d7ua���dY�m�6�iJ$��٥�F\É���,m�;]��$�ڃ���1V'�E(�bMVow��+��5�\��:?e`�f��G��M`Z�1�\�r�g����0�8Y��%�#�<���]�f�zaM�1�J���\��b?M�����N��*��<�|O� �n�� �JP�k����Vj)=������*[��6wE��*�0�����
�����u�6��t�p\�����,��h:iH��+:���)7,7���z��7��d�Qi^;Y����WP�SM�Q�K���F�~VF���0n�Z(��Wiٹ�6=֥�Q��?��1���������pT� �qHr����F�<p��V�OjD���h��b�2B��)��[-�����̹��n�Ӏ�ҁ�$�"\���Wp��+Da��f�p�P8E�'���+;1����=���O)�9�*�Y�8�m �:����Јެ�m�>�o�w��xcjb$.�B���V;#Ӫ���5�Ǒf��u ���P����$ۇ�v�?i�h֘�ؓ����QL�ޓ'��' �i4�啱�w����0x���׵��=O�E�H����%��+�qB o���;��S��M�}���!����r�ڹD�8�<c ����L�� ��P�����uM���^�I2�1��2�gs��'�e���q��,��}� S�S�v�U��$8�nC���Jnw���>\lkt8���0j�su�������'
 �9���n�kp���B�B�'���s	>���T?�� �M�a=@ڷ���.'�g6l*�k�b���G$��Y���RbA�"73�7a�X؟��#Ӈͤo_TE'�����|9��L��R�͜l�'��s�r��0 ��!g���F�{�	ߢj����Ϟ3D6Y����E�k܂�}��O ��q���C2��t*���U-Cu�e�8�ƪa��4�?�9�}�Z�����z}�5�TG���r�eG�M���	V��0�Mr0F��!G��j�P�Lk`ȅ(c��$5ܳ�"T���^A���A�r/MW5����P������?.��c��M���!����Щt��t�������� �~�l��4�J�mn�V�3����)����Ju����9��T�FK N��[VP+��W����W���d��.Qd���{������t}\��:lW�e�-Q�,��=X��ȹ�ן�f����K�Ȱ�S+QV�F{�g{���`7ܓ*�¡)�b���EZ��&��A;oNd�lY�ū����w5 ���֑VP���h�L��L�#��IV������ ����Jv�9U�s_�M
3���B�ܕ<�1=wH�Vю��̐�k��++�`z��II��=���(_�hu5�P_n�o�?���:<*�(l��`�53'�:� R:�K� ��ݱ	�&V㴀�>#ì듿��Ԋ^-B�V�\�
X����f,Ve��aG{�m�`d��9[~�bѤ83�ȇ��:���+��5c,.�ڥ#�ԑg����:��D���˥��q9�
X�ıV������_-R��̓Y�?Et"8p�r�"?�g�.�A�M��{*���!J��޷Ԣ�I�F���jA@�V��$_[ж�T`�Nڻ�o�NA
�ɒ� "�i��?�E:L��r��t�� s��Yc_}�YdHj�niGs�R�E�֪ȭEu��F��J��8��F��Dq��RשU�>�*V�#��6T0�]}W��s����t��������b��e��N.rJ��eY�d��Y���%��B�j�A�dah�:�D<��N��J#^/6�pp�>5u��t/|���4Kxt��f��]W�	��Yc�E!sO�� �\!���3�����3�^v}NZ\#瓱,���ӝ{�٭����꼑g��p�J�h�G�����9�F�Y����a��g]����%�䍃��w��  �?��er-;\�
�����7e	{�O��f�٬}L|��Ӥi[%�'�W���"%�:��c�z"j_k��1��E�F�S��^�_���-�A5��C*����X"�����1£d��{q�υl��4K���|�!�S��-�{�xPyn3��}�j�@V��u�\,<���� ���,0�"�B�u��~I����E����X�G�lW}{*��(;�>6J��C
��P��ͶB|��� ��L�fr��ڱd�[L�0���\��͡S��%*�&�X����eB��]�?�����������0p;�G+�p�pN�MRkMw]�lpKw�s3Z�K�N9m��s%��8PO�:1{l�F�^��q"���q�8�%r�9
�"��ÑQz߀\�cp��q,�otS�|��5�*���� �Rɯ����R+�X .��&��¨
߳�
J���ؼ���9�GA@&��W�S���zmu�����J�fp�	4���fzv�O���QQ�h�]擑^Xpc�D�r\6��2Ƕ��F�5w�����5��T��1NR��!�Y�$&���o{	w6`�4����a-Rn��munK�8bGU�y�uB ���b���2l�r;2[�L�����S�qs�}�yf]��Fܐ��=��Ù4ϓ{�� ̬��]� 
��6gc��ц�ׄʩh�=�(�#F�/׊��R<��5�rA� 2<J��K�MVE,��"��m�*pE���	o�t�:�	��R�!뫹����f��p��jx��K]�b�Hhq�IڗÊ}ݼ$"&;;�]�W���V։w�V݈x�Y�0�N���V��k�"��u�RG�0R�D�ˠZ�&|�h6�Ģ���p����	�h䠓>>$! م[��1��F���A�9��ocp|a���2:F%�_Nu�;[�dc��"�DS������1�Q��W���|�r��@�;8�#��S�D5���q����7�x-p4�]uφ<OY�.��ϫ.��9q��9�%�ln�	�V~%�M-Tt�O0�1au��&�/���*:c�L�p�9ę��@9[YK��r�#��y�q8�l�94t5�=X=l;���Q�f�g�/�3$�t�-'����E铸�x!�0eWJ4����P��r])�0����� �O��'�������c����ZN3�������Э�l�py��Dit?�U��uQ��_8�X��vQ�ێ�[O6�k��@Q��AO䐴��]��t.���a����
�? �BP��=� �}�ɌVB�2 �%�5 O�ZD��p�!=4ܮ_����l��.�w�#e�f.D�5e���1]%������4*�Z�M����5�����ǎ�7�c��:�F��xߩJKA�������ة��3���ؘ��X��im_�p�L���g�R�(]9p�]D�������ރN��|��%0G�7Xf��r�{h5�dl.�����7�Ig��� e�<�?ʅ�v�q��ms��5_Y �ۥ�|$Nf�uAq��Ŕ�8u�@�u4���~[��*��J��V7�F(�ѐ�t�%�lK�Ԥ\A��b�'�)������tE�K6�WP`�9iG�?�Q=���ܳǝk��i�޽u_%��k�Jv#��%��kk0��N�ý>p�M���4�w����t�P�K�V���(N??v����o&e�B�)��TR��4��!����fF��@$1$ni�q�i��P�����x�]�˃�t�+vUo�PU ���/Hd��!0��M%Qu�P~ݝ��F��g��x�y����*08D�e!�wh�h�mr~��k;Pl ��U�xF�!���G�f9�tt� ��C�0���g�%�b��l���P�!�i�����|��6&6�;�Qg2���8_�����δ`׷ۚ��Ф��c|`�6)78�@}�W�����8�V�oW;�CFO �>�Ǖ'����d5[�q|]�Hu�jx�>�Y%��$G�+�r�^w�.�ٿ����UL�Ur2&�����jO�ё�Eu�2U���͎ )��
�H&�\����to��z-����l/;��N�Vl���{�s�Z��[�g�BNXO$T<H��%�\��Q-�`|Nb�v�n���o0y�Ɨ��ެ=2a����K�zx1-*h/���r,p3 ^^1��^��r^Y#��ݒ����5��}W��+
���$x�H�
�~�]�p� �X@܌��y+5�òG�כ�&��Ǘ�`-6$�©ԇ����i��h���2\	�5�*b�uO���#������ܗ)-C�\��P$
�pZ	���y
��̼	�0��,l
P��p���s*����.y=��(�
�D�5z�#��@Y�M6�|YK8�Y��K׉��?���!h��i׳:�>N�T�s���U�U3�?}��4���J�rIǹ�zv�^_�S���:�}i��)*ࠍ%6\�pP�b�X��ꈕ���h'�!nO�?�� �Eef��0K'�w�	\�E��8�u�Z��rw�݊���ԗ��@�P���Jj?ӂj�$�)�lv�Ż����i>��2��peUMib����6����-��Bp�!_&�����#��r�Q���e#针8�������h'!(���s�૝6�v_´g�����q��.R���ə�M��*,����V6�r �X�`lX7���Į7�+��'�:(̆D)~>�H��UC=�e��ͽ�֤�%�%�	��c���JE�<�ی11�_��#`c�E���վ�H��y�:��T�3�n��a�虢`�����8�g�QS���!{5���gy+Slv���=�'�xf�.�Z�1#`�� B���5�1
g	F��y�|-i�<x��q�.6��;e�j�Ssy�G�vy;1�~�צp�:�,��42��מ:F�J�p�� �J�U�2�~�-�'w\[]�Z������z��e��,�EWI���M̞?�b�~<������ZHvL��^���l!h}3���W�b��eֲ4г�*�;x�������F	��q�	��V��3�79)��i��uD���<����$^G��r�Q��a�R�&NS���d��W0��L�A�H��M���
��'	R����k���t윧�YsA���U���^���`�q��me��� Ͷqw�U�F�U�������9�k�Hm�0�v���[3��4��Xs�B�Վ�9�k�	o|r�S�h�BPUm�E�ȵ��YBKb���11іf_���P�;�mx���/u3i����2?Y���{`�4�P4`�96���U�q����W�-eqDr�D�CiXMf � �3��۞�\O��G^}e�� ��$�0"�6��2���'�]4~<y�Q/J�����M���3�xH�����O0}��;�E/� �m0�(�r�+ҘY�
�o������#�w����<��lm-2��.��49��]$�I��4���ge����
lX�ۑ�s���A�+�|@�J�@��%��Q%e}�Ǵ¿�*q�n��N����e�>8$F�QG/��c���XR�E�5�糕^ ���Ō�������
��O�ZeIG�in�(�E��b�۬~_��u����D�d��A�r��q���xsCP�oKO&ݎ���V�3��)N���[��.�[��ݭ�P�y4kg}q��M�ү�'��@]-i�
s���K�Q
z�dY����-�S<'#�Ae���4F���g��m��Z�[����j�{*�a��'
�j� >g�ǻ�������}X��RR8JYy��^��͆�k�+�9�Xx�S�l�$:�U2:�JS��&�ߛ�dX+��<f���"���l���k�)sVo%���e��Y7��t3#���-:�xK����)���qu�|hw��Q=s
&7DW"�r�`��+
��+�䴗�ȝ�C�*?��;��gu�5
�R�1��j�g�+��1����}�U��A�2��$��U ���HÀ����\s��������5|��QŒY������G_�2E5j�|S�#�qΥ��Jj6�5�hCh=hƒ�j�	��k8�Z�3�ls��Z>)��	 }�o��W���-��yS��!r�$�����4/W8�L�މ�$����^A-�<�)L�r񲓘�f�:	7�ﶒ����}��/)۱F#©�Mӳ�j�:3mq�Hn�o��������BmX�6޲���� ��IO��Q������:4� ���(&dH~�BE���_
M�)]�S����ظ�KrF1D{Ɨ�ߡ�����CF�Q@Op�J �{��ğ��N��1����#��{�!�P�����Sy�	��"�=a6����B�f =S�_r����*գ�]722f#��� p'<5�P}~n�/���f�=�Θ�@��m|���k0�'��;d���'O��9�~�x�?�>Qjw�y^f'����tM��nG�t��<Z?��ɍ}�{�~�eQ]�Eݷ��:�얿��D�Z�<��o����u _M˺�c���I�
6l�w�rN���"��	�	�P�OL-p���7��; L���ODz���p��el��=u�y���sJ�:*��n����ƀ$��`V >���jhKK.Z#�,���{���d��o4�Y��gy�$}�ej�&#�����If������b�B�F�ׇ�N>�^���:���%淦�3P��������(f��iqI�0�tIr8���b'���N���V��5�V�si&��s���oKi8��dW����9��B06���=��ƽ��yd2r�[n� _��/qg��a�����9D��"/:���C(�rX��UR��~I�dC�(�
"%��~����q�ȭ�yؙ�Y�t��xY�^BG�D�eH��^��ӽ�fĆtW�@L��ԵyD;*�1�t���PG]rms�Ҙ�TQ�x�h�`� �?r�Ň����4��V��;�0c R����&��0:G��)œ朱nG�ޮѓ�m[w�͹,Q/2XX���J��VR�1���T�?1�K&g�KB��
�?R�y�i�� �-��D��_g�û��^-\�]���\Ь�u� M��c0���Ӗ����Ѻ�O�J��c��3��.		aD�pz2l�Gq�פ$'|vb�_���8[�P(��['H\~�;��'�a��ό���{[�3mǟQ����b��?�f�($��xq�]�DIxi��;Y(e���c�
1�'E�xέ_H�D`� �+h�B�K������p'ZŐVk�YrX����7򭁈�uI-�s��]�ٮ�:�!����Kb6���8�+U��-�Ƃ���â)-PO%okp���-|��j�7��E;f����������;e�+�	uylx�;8fvm��tZ܈�
�� ?@,���Q�H{�O6��z�SP����ѷ�E[��rn�΄�ZW#��p�&��{3���l~�� x���h[�r_�+6�z'B�8quR��TY���eN�00w@5]{q�֓G�5�i��Y�l��,��,�>[�y�s��v��ʌu3ztX�T��7�#y_˕B�R��FĐ�'{�BW�ʹQ�%�SA�8?���TQt�` ���װQ�7�(��J
���`�k	4-(��:W���HޘC�׮"{�%r�������k]Ī�]>n��$��.qn��\Q�"UQOMe��`�k�� �H��H�DD���~UY
I*����Z��=�&o���"����9�Y�a����ll�e.�.~3��O�����$p`�G���&��5���8�'�T��4��Jϥ��<��B�o�	�DU�J@��rm��QY2��N��|B�%��_l*�83WJ��������Ew4��;�M�r���g�&A��i�&1�Vft,� �_�h���Nr��Gn��%��ur%0�P:����b�F����Q7�WMЯ^'��s5(��mg�N�18�g5�qGѵn��
�T�M�h�bK�L_c�H�7��
[���@����d$�Wޙ�+QU�wh��[ls�/V84�ޥ�ɽ}y��x&A�9�'�%�F��_~��Q�l��|�`���D*d�[�^E���9�7�:^��������C)�y�q���T,�"Џ����>m�Qg�"Cȇ���⧕vQh,*BgJ��M���o��.�x�d�V���ú$=!����f�4��i�����B�]��gz����a|�8ם�݇]#�SR9/|P��X�
�foY�s�<�ӂ4i���}&K���K��P>`�Q&��m�Va�C�L8L�WբO�!r2M���=Բ=��J}ְ|p-MU��"`�1�'���������ݒF��kɂ��i�;����ht�L"��8�s���]�W�PM�IQ����;	�S�'@<��0M�)�~?�'8&����U0sXkE;��A�8Ӄ����/ܯL3rM���ȣ�w�UiĮ���W:��m��Z&�m���3��|r�)e=%W�UΧCխ�\��Y���׊zD�����)	���FR�������kDҩ>���A��pK�>�c�miL����Wa�	IK���-ZP�ke[��#�qԜP�e9v[��Z��&��ꤊ�5�p�2�`��趟��TM� �LgKj�e�_5�ڼ#�E�n����'c�;=ၺ~�c��f�RJ٣��6�Q�Js�W�W���,캐I銾X����`d��*E�!մ�Y.3e�6��v(��/q��+4Rv���`�Jn㲐�n$��+�J��V�6ڤt�T6l|��U�#e�6$]vN+gP��;$š����w�k)����Ajz�*<�0^��|����~��@���ow�)E6�A����RWiEv0z7G:\��
����T�cǍw1�ZR��ڢs��QGBc��1MU0�Y��_��ӝu�昉Nd�m��_�����Z
���b����+&�;�@����ԽvHY!�������c`Z�2>�����i�6T�}o�y*��c}��^u��A�XYN��tɷ��ҿ����7��Ʈ�	Y���5�U��m�ԑ�28VK��Ŀ�׮y��@Ѽ�[�ڛ���L �nLLETgQ�DM$kÔwc"F:�>��Kֹ"F �09J7�@ -"$�)��h��;�
f�U�~%�~�%�f����E�5�m��d5��r=��+�����z���/��#�V�X�j��~�n�;��)�L�g^췷ns\Fl�i>��,M�����=�2��L�&��>)͇�>�bֺq"ي	�a�KoD��@�3l��Tw�仕�n�Kl��1�:�E����d�U�B��M�1z��=׹2�Dv���(�D�rd��ŬO��E�V����s17��mOc�i���BK݇F�(徧���2]����4���b���}�����_��|@���#f�d���;�Ҩ�%�B�ATL$�TlF��s,��~ K+n�@��XSGG�e=^�ACyR��,��#�$���vh��«�,�Xf�+G_Fu��"}�y�,ȓ֜�k��(QLӵ���߶�����פ�Cs�5�����c��{-v��QdQ��)�$.�]��P/I��
�&
���4�+���3.	�����	�Q+k�jo���fL��[M�1S���dY-�U�l1�}vooDG=1>�4}7G6u!.���&�X���fm��Y%%�:�JIhkD�����R*�s^_���ϳ.�� q2�Q"�s�G.e3��I����tGV����V��E����H�����ٗ\lRt&0��߶�q���������&���P�����s^�l-(f��f���8�U�bi��t�Й9%�0�µQ7ڔ ���B5����&xFNY߁5�C��|fB�L�M���RP-�f}�>��=�Ǌ�2s
����������<��@iaĽT��j�t��=;>�Ȕ<���S϶d�����L䟩7�H�z!.�(��hf����˚���C�::5���T̈�,T#o�¼��q����YiC�ۨ�����D�;U%NL�L'K+�$48_h�B ���S��{z��`���0F�w0%MIҕ~��X�oH���i=�8����Q���ri��yp�-�l��<�c,φ��^���Dr�ݵ�9���G����W��ϛ��qO}��ʺp�T�������yM�|�������@��]���O�L)��sz�C�5���I$U�ytW��l9`���(��Z( EOuO�����-¼�M�z.kQt�M�ı����\�\�;���b;2[�P�����u��	�,d���~A�����e�P0l�@!n#A�ӳ��n%1^QnسA��2
F�sW��c���]4S�����O��_�VgY��ؕa/�Ǵ�u���V� ��O���|,�������Zg��yɏ2��`�iԷ�H�Z;�U���0��U��$�M ӑ���-��y��a���1��%;H�^�Va/��h�=�LEHH[?�>�E��mV1J.��B�$��zWʏ�:q=�=�˾t��b�����k����������bf�6"��<!!}�*!���)t�-��zȷ��X�8�L�	"7�ӅNw��{�M�X��"����	ˠ���
2�����n״�3�Q��p���L��.h�5��NA����H[m[�7��ާLjz7�=R%�e>�!��ͬ��0�z5��!*��<^��Ά�"��$8�qo�!�\e;fs��܊��'n�3+�/$����5`����*A���im���ж4�\Ug��Wʱ*"Q�pͷ!�7��ߡ�����W�0�!T��2},7�{t^���� �f���jOo<��.��":��_|39���֟,ᲈ���\��>�]Z�'���Dh�M�R��KRT�q9zuVn�%D^'�����G�W�6��(E_{��wW�0=�)���BI5ڱb������&
f�嬫X��I ^?�G�% t����rjy�x�
�UWg��Mmw�Q��k�8���J}x�YiP���3(���3�\S�l �S�'��K�h��GQ&�4|��A��8�	��Hh%xs'�:G�"�]��n���m�P=ĠO���Y�L�	��"@K�'���֥c�}���cG@�� u)oZ��`v@���@ǵ3оǳ��f`���k`ʱ � � '���O����(���⽃�D�3��ή<x��++k��ܓ$t���6kr0i�(5�l�	�&n'�~
��^3�5*�.^7Eɦ��#����$L�����yq��Ү�����֦B��^������Tru�����)5��ݾ�!�t1�!Y��Yr����t�BR��Xs_b�>2jUy�D�r��'������������K��Qv"e9[S���\���2J�"E�+��s�! b	J;mN�(��*�3Ӱh��_AO��A����G=r����i;�^�	 m?�d��@�k[,S�v{P��\l�|�l*�y~ UT4~��6T��D�8�,	�`q=��b���ٱ�*�s�DT�h����?�L���b�t&`S-�J4zu�u$�*^��R��s!�u̘D8~����3r .�Wܣu��M�]���ρ�{G�<�ho���G�OER{�}� )>��n8�$��P7���R<Q(>&w��e;��M�`��R;�1C����R
�6��R�!��]h�8uU5�,xopM�a�Z�BFϱ�y�� �)����歜�zCH��LІ!�/�݆�N%�*\9�54��	��Dy�$ �'6��h,�-*���a��ep�Tj��aS�?J���T6�f����~1Z����|���u3J���Η8c 0��;�1�5�qP�����-&~�!ä/`���"��;7�o{�5W{
�zr B�6"��R��y�V`���Ȧh�љ��ϔ��ԉ¿vj�@o����c�7F|�6���xq�h��.�WN��&`LA���v��rܚS������+��Q&y,�K�0���#���y;3n���ɛ����b��7�<*�F�3��r���Q	V@�J����}�/� ��:XB��L�|�AӐ�Hm���O�Ԇ��jxQg���xV�#F!|+\�"�u]U������U���4#	+<��W����R�p����O�ҡ�j�ç�U��蹱vV���,e�y��=^,� ����t�B#��!��X��#]���R��6leO��$y�h��;� S���4Ѣ���HVCa�R�z�h��M��%�T�phi�[Uy��V,�Y�f��.�~��~YMθ1��@�C�S#��J�V�ؘx�hJ^U�]/��a���S�0�#��=y�����$�v���)�j�
.D���N=�&$)ˬ(�O�k@lLL0wҭ�Z�ۈQJe
�����K}�8��c�,�KU�u�Js�3A���&����JW����0`2s�"= p6�R��r7����l㚏�R���Y$Jk��� �C�z��7���ń 1?h>�aa�Z0�K���6�s91j��Lnt�+���ir�Z�"�1OH�;%,۶�1���է��%Kw�j�u�:Uc{�@�{�o`Rpݹ�h|�F8*�BYLh��s��MYd�)M���`#)&��\OOC����D�,Ⱦ�����i��j� ��}F�\Fd��~!�$��)/Yc��������ǀ�e��?�j��b�(���6ɐ���ȩs(%j�bh��'�{`��B��m��KB�-5�P��'j��و6.b]/���N�b���{��_�X3��!�f������`o&U�T��8`(I~�	�2�����|<��&T�J`���N�/BA��I�eL�$BR(�g�^��J�������X�F�N������z<bX1t[���L�J��yE|�m�6�R��x9*ݺ���JY6��(�y��.E�Ӯ��m�"aYV���7��\���=�VKҡ}�Fᶹs��_�\�rN�@�>dG�h�!HdH��GBa��л�b��B�Z�H`,��ƙt��dK����?�8���Ѓ����kI_����:r�:ܔ$>x�����N�L�7q�5W�{�IVz�nv�&�����[��v�i��=6c���>+��H�0$�`Ae7�����d\Q������_�'ըӀ'�%���z�pn�Wm�T������c)
;��R���S��K�0��waW���h8eK6�'T1c&�p���|y��ZH��)Yuֶ�oL7Ap���w������6��
P��P"y!}�2;��߆ק>�+g]]� f +q���uD��5�˗\�!�v�TݺW�
�_�p�*��1�0�]Qj�aD�ni�Fh��X�9E�h����m�qAR�r���	���aj!J�}[�o#8���FG�K��Sf7N8ѠA���3���D�����f�|�v@=��(�dsV;�RV���k2���ۨ���F��[���ߴ�R��a�+��&�KKZ��q��iS*>�ex9�k/�����Ŷ��f�_���jo[�����ɮ�sd�I�Zp��r��$M��Ŵ��]Y����Z4IU�nM$��Lg����[��9���E�W{Bbmh�9aޕ1��B7��V���̫������F�#�Ǥ&!Cs�&W���X4J_��|�Q��b�}��
O.��T��V��t-]7`�.�x�2�3�m�hpp�HdY�&��J��z=�v��5�X����+w?5�Gߨ��&$X`�k��U�Dh{|�`��v	
%��V�4�� -W�g�X�<8z�Ã΅3�8�x�xQذ-V3��g�o�/EҮE��6m_��T����g:�=_�T�9�T��Ζ��<֎�%�s�X#���fQ�Lzm��!���Wp۔����ކG+U�]Y�m�;��d�C 3:�� ?����n�2�
��x+����7����u��M��n�l�1���a]U$�CJZE��f�$�F�_�#H"��)�"��=�:�R*����.�������.}���:�i�M>U�.�wA�{v3��#ӵ�n�ک��j"��뀌to��Ī-���7�1���ۂ�â��5�w����8���v����b;2�4���j�e��'�?(R�/V��	ڵk9�o��g�E�%*r�4���:�#���`����b�l�Ԅ��A��l� K�l��d:�A��N�v���f���
�ds��Yv��V{(�@E��nopt�Y�ɿ�˔�1�5Ԡy63�I�{�e����槵���w*�}��C';�i��[����aw$�_fv���\�����Ͽ�{�rЪ�ػ�Z��I��<�9��%�d��m���,�}��.O��7Q�

�
:WA��1R���A54��B:jP��-�z�Vޜ��w�AK�{�����°���|N����5NU�pG��`�r���/�{�*�]���=Z��_���|�KOS��«���g�g�-��p�j:\���� ����yQ�D�2�k�d31no?ત�W��uP_B����;�  I�=V�~[}vLæ���WnC&�V��H	��Ǽq���Q�t���k&]�G�w��IlF�$��W��9�c.m�i�G��Cq>zFB�Q��{>X�"�b�")��P]�rM�#���:�̿�������z�[�u���.�Pap%�>X%ٓ!�����?׮(����m����ͬ�{�	>�aM:�ڸAKW��k��p�ާ袷�D��o>So��I����>\��08F~er5�5�W�,9*T�H������i�5�e����q��(�>3K	��,�`p�(:�#��e`✪)Ӌ1mD��tw���`������	�ۭ���� �6 ��JH:���A�p�� ��/��e���ҶƉ��/���l�un�I/q���n 4?�먚���InK'�V�q���D��@���k�-��+���B��:�#����gi^�����Nn���p�n�2@1�8�����L�0N�u2�D��;�±t�����9�:�,a�5��E�w���$]0P|���T�	�e�X�DU3�P����ad��m�&����`��A��u�1������I%��CV�<�T��S��U����/+	/�k�sW+��:��팲�����J?����}-x��FN��u_�|�bK�M��穦�-eh6Nw>���u�Xz��e�`�ް�R�{�E �6M��AU����2qEG�N����m"�#\J�=�!l)m�á��j9���ۋ�[ǜ�7�}�j(*6�Ԣ�|6���P0a8?6,�g�93�8-��d�3�}���WW��]�M������H��E�c]B� �(�#�*�.��g%��lj.e:���'=Rf��U
qq*��d�sɮ�<2V#�:zg)7Nd�J�\���ֆ��:��I���4f���	@����1)�R�{V�D�`*��[ʁgLlh��9ѣɓ�Pr!�E�����n�yP	�����[��G�$Ҫ��KM�����=[~��t���u_1Eh��H���S1V��<�	�l��KrB [�M(0��cN������@��H��f;|.�hC��C�m�A�\��6�y�_�2�F	��8 hx�7�ό��,tc����U��0�#���ށ֖�-��F ���>���E�1F+&�CJ��-�҉p�O�K��X��H>�O�[��u��$ǭ�bs�nOLV��[19zS�%�/��y��Ț&d��y��	��K^���w����e3�2��9�M��k�1��(4j�U?�f��E��y3����@�aX��v����,^hQjM���2
�;�!�p�+� aӐ[�=bf\�u�a6]�<��N�^��T�t�oa{%ߙ��+[�H*�����ă4���`�V��6R��6m/�Z��{'��o��6���G�dw����i{݇��2B�f��Ʒ�����f��e����Gme�tR\�Z�nѿ-@���n�v�49�>�d��ģ�B���;N�y�-�$g:iJ��g�>�"���ն"/i<����y���:k���X'�Jm�9�`,����7"ٓ�%��y��r۴m*q�:�P��>���ul�T����(ŷk0�s�y6-QV��M#'��C�S��Jx����Z�I/+-@��p�ՋlN3����_H*B�l�[A2!d���>���(U�)h�`%'�}'��s'] J�QLu�l]�-8J1�xp��~s�CD�H��#9�sMO2�M!}��LPu�^�96c�A���S�PF���*�3$�o�綵MR���.�}Sh�Z�%��d\��qt��;��;70j%J��կ�"9!��Ħ��t�s��s��U�?"�Mqp�(1����������j>��:M�@Z��q�:�#]����Gxp���KVf�&���,(�I��M��~Ť��m���bɊS��#e�H��%7~ ���U��x�
��yZR4�a�\|	Rf��$�œ\������P���PvQ��Wc���@Iv�Ŷ�e\�5v	���FS
�W����G��I)�ǳSN��`��=>��ф3��c�\����lJS��i�T��B��Ff~�� ;���df�����Rn��#���ř99���
�X7Fn��"'"Ӿ��x��C^���/���+�NL���f���>�US<�!z_�D�:�� �[bLB��'����6X�	k�k�����P?��,ԫ��hK�ҡR���{Ӭ썿�<ւ���L���bb��F Z�a���L��S�[?`������,Z2u�y5p��v���q_j_��A�H��&�� k���k��q�L�W��B��$�ьTn��2W�M*�>	�04����!�;T�D�����|�Xs����O�����\� �ۺ���H@��q�?уy��^��">�_��G�<�oBH��y��&j�bK�.8F���,Or2��������.3��3.��ة����#ɞ����}
��I�]�۶����x.�4 m�e�wI�fn�³n�.���\��y�c�5�qj�`��z?�� [��W�����ida��Ͱ�����H����c�ݫ��T:_ŧ������9�?)4�1R�-?ț��J�$C�����n�$���1��I�L�k�*�5��*�k��Ӄpzς�9�ҿS��i����A���:0C8��TB��0�>O�6�75�-�S	�Um�Ņ�+�%�v���z��W�R�u% �L�������T]UC�A�' �Ȁ@�N�_2
�Ze{̿hp�"��2|��z�n@��G����o{y�� G�5ZP� ��i��F
��!�F��Z?i�p~P��jS�8=�s�v�[�>�7@��5x�oM��P� ba���t�&�je�8�Q����`����Q�@P��Z�W���/=� !Q�6�M�.�z[;�l��CA����pO�1��C��;�EF5@�Rx!=/>�@�"'ƕ��z�y�jG�T�a��T�X2Snw���ؐ�yv��O�
uq�_��`�9?�M�`[�yQ�?��1)K(#��'��j�n& ���<�����C���"��hM�l��Δ@���Ծt����`�"2��#M+���	=u��*&���G����DS��	�>֜�����6ڮ�=[�1�j�C^�2�Nڜ^�f��E��j�c>Hp�U������0�'ܐb/�i��rF���~'���_�� یC�2�A��W������КԼ���(W�������HK�`��ĥ��*L��"�4
g�)�;O8��Z���,Q`�뢛+�x��%b5;_�^wz/������� �X+m�)�a�啦~�U����U�V�*���kb��O��o8��B�)�i��5�D�\�ط��-����`.#ϭ��6�Ç�]8�#�ݒ�n�6�`D����^Y�6��Y4�᳔��u�m���Y�[���f&��tIY��!.3��0��(O��%9LP���;����*8ު%,+W*gX�Q:4�&.�Y�n��d�	��6o�pk1�^�~�~`�L��ر��iu�/�̰���A�4H��{�pt������#4��F>�	�"0*����W�?�2���Kw�|U+���
�n�v2Jsq��3�>"�_�� ��1��G*iQ8`�~IEϢ�=d���n���A�B�A^F��#���6k���%Q�����R=񲖕�p���O�]�]�-�e��X�
�qV���}2�[��~�� /C�+Rk ���<:W��q���G͋����J���̈vx"]���|j�Iȥ�ؤ2Y5�'�4������yF�?�}yR&}�p����q�w�ԩ@&��TGˇO���k��uư4�=�v�dNo$i�;��Q:jS�ڃ���zͻ��)k(91Ǎz2�]U��$���_��}з�"0��	dӳ@.�����cn�d[��̝854B>ɋ='m�9`���9� 9Y�,C(.�ɮ�G ��I�n5m���o<+��E��a���n�2Y$����.�N�;��Q��{�j;%_�߭G���W�L��0�[\b�L��� ���+>���zT�De�F�v�Z�,\�ƛ�^�06K�=d�
�4���ȟ��h���7[b�\j1��_��Ĳ���.����ۼs�1��]�p�B�lծ�!	�i|�c4,m��/���eT.-��2�#�%�d��,~?��d�5!�����u>}q�-ә���SҲ�K�ע��U��3��������}�|'WB����B�%�F=��g��_��lm]��ee�/�G̔"�����X�~����z|���������|��0���&��=�&�҆d���?ÑM��\���v
<�4��R(�.N~C���\L1-�j>�
ھV_�)�|���~�$3L"�jdℹ��:�hs�
}���%bÎƺ��]W�@����		RŴn޿3�شxV����|1_�����u�3	�D���>8��B���LC���>�>nu��t:ԉ�:4@8�ٟ�i�����-�'��/wT����6
	��dx���*�Bhprw�
�d9�Г"��l3J�Ej�M��KtS&�K~MJ3�����b�#�j��Ml"��?��y������:)Ɵ����c����j����/u#t�k�N.XU7834�<T~�p��l_�e��I�c
�GD&i��������3l�GQ@-$6bխ'"�=對��~��B�Ԡx���>���҆�/���ܩ�-�H�>Ґ�I�o����e9�"k�|%5�P~��&gP��q�ۜ~���'z�)�KP���B����v{y�%��j�[Bb�5V&���o�baItI^�@fD�@\k��9���Ԅ�����*:�F}(�gm�ʶ��X�����g��&d$z��?� {�a32��)Ȣ�����UU�>��Rt��o#�Vu[^�pQH�� L��N�?�����a���Mp|�m�q2k�*�b��&+��Q=�źi,�@v���ݦT���Mq��}��3>��(F��o����C��O,�ԅr;3ΠI?{f�dŜs��+�a�g�*5C��9��wY�,�ӾKV��7���{���a�b��_^I��$�IB޲��FD��*�3�^?�	���Y�>bG|$A�ണY�7cm����nK1c�Aը*9=��j�1����iv(H����N�'��oK�&�j뼨D�� �.:��z����G��a$<{���g�HFN��Xm�N�D	�w�i�,�d��{z��(8/z[1��㌷E	�h6硕!p��J���b^
]�ϑ-`����C���-� ��Q�>��$��8k��D�g�����tG�E�]�^0�tQ�?x����D��I�<t��u4U���0}��P����� ÐV��Y�d�����;<X/Sk���۱��@���]��> ���]���(Qq�C�/�Yd��u���(|	��΀`Τ9�����xZܳ��2^���I���*�f���P�%�Şh�Wd_A��AF ��#��j�];�)(�L����4&^��B=���8u�ctQ�^Xų>fµ�rE&}�?_Z3�@N�jvࡔP����¢���^���L�ň<��{��k��$��&��:�<6E�	Z�~w~J���dkX���0�Ξ\�Z����?�:�3�n}��9��r���$���T�}�|̺��+h��r�\�����<j�V7;���/�����+h���ؠ��ϓ������͏
����Ԁ��'m�q_�Bc��8�v2��a�t�m��(/��6'�X���f��{��s��<v>��Z�h���2+뛏�Ϫ��PV��w�K>�'*(��jm�:��BMg������Ht���L��h�m�DO�-�e�k�.�לx�D�*�� �'nL��>.����7-��q�k"�E�e�q�� �����������x�k̞Vmc✵�9��_dqRU�ë��rP��~�BW�&��-����m�I��p.��rjazF�a+iC�E}l��2�^�� �i9�l�@�kH��hRP�gC�����xڦ�l���l3�/���͋�B"t=�"�����i�-��Dh�|�(��i����X�^�1�'y��ou?���9�eh�<��?��}eʨR��h��m&�]�."�":��<����]��?�s�^�g�}�J��!�nd�Ԫ��5���<K���Ki;�H�<���5Z���{������΅eQ��K5�d�����>B��WN*��:>�q|i"��ۜ�=����;wq��/#�kNl�r�l��FYH� q3
Ҷ�Ǎt&�%g�םƟy��+N����qO�ﯖ2rd?���+b=�$4����\h:%%�	�:w���S����Y9#]�[��I��SL~ŋB,�X��-�1����~���z�b���O]z�0N������k�7�-�A�u���-�,\� ;�sl<�R���ե��ዲ?�t`��Cl��V~��|, �l��Ǡ�p�?}uR�b���'�I}�)��"W��`���!��Nʃ� �t�za�V�ɿ];��n퀧VN3I|l)��@\��yN��y�}j;V�-�*�'�q�Hw�%BKQq�����?�1pW��0C�ۣ�,��=�����J�����*�m�s���u8"0�����f���!ҁKq�I��*�&Y0=iU�j8=��_�5��A�oFx/�QG�E�V��N>:�:�K���})Uf8�*���v5U8�[o�c��t�d�n�tBj�잖�D��o6�f+�ՒL����(QyC��1KF�@]���Iu_YK��i'�E
���;U�pŉ�_�_T�2'�P?��A����)��^~T�8�sW��LH����[��}w��:���a{�·i��N�/���)cM��NjbF��(�p��X��4#��� 	~,�A�^�\%�׋�ԏ��I�O�������!t�ǽL�8���'�t�#�
��]�� �5�ʆo#}P�ݫ��e�A�R�aK�"�����@�\4��.ٚw�m�N����w���F5R�OO�L�L=UTl��[`h]@�nZ �~�r�u��t
B��S� ��
3K�긣4��2s��g^f@>��x���eBlq§B�#�0ϽcϜ����3&'g��R�9���݌�~�, �t�AbV��$�kq;��sV�%�10�������n�00�XƮb7)8G�t��j��xX�.�F�o��zVJ��*��+J�8��3���˓	dgVWn{��a8|Kb#�p/�3%Ck"2]��K����v�ItE��柮Q*����Y!z^�	�V;uxʛ.�9&��ɵ;'��^�D`(����\�֍�������j*�&��~��'�E���x�uȄ��hw8���%k[�`O�uj�<p' ���{ǽŕ$��9/t��pJ*�,��-����ͮZ���k�ͿǒՕt:O�ȖS�X���>2�4j��p#�yi< �$�e��곜^�G*�N�-p�egqS�\"cӔ��٥��0�L��+H���K&������L_����r
v�jgs��:g�`	uB^�@�=|II%mol�`�y?���o��hxv��k���@v��ӌC=}���ͅ�$&��b�y��)���<��X`���J0�M�L�	N-�ͅڼ��ΒH�kE�Dm������~Ѹ�fn��nj$�Q>9��1�]�$�r�S��,"��V��Z����c����tl-�`���7�Ł�
k�1�u
�� ��;~�Y&��qٍ+N)S���!*!�ݛɻ�8��a}�||�0K;��a�U�c1�\32����7���v��)�V�5,�h��j��iD;����Nn�L˟���;Xq�2��K�EBr���4V�E����<�i~"M����v(5���
o�`m�`~�o��Bdgj	�f(%�����E��$b��ja���@Ϯ��?�6m�s&�6&���:?~�+x&�1XR�>�&[LT�*����Ո�W����:�~0��n����֢����aBd����?c.�*2H?�ҍ�gp���x�@ۊ�P3��\��zC-��6��#q3�Yѽ-���� #��T1�0�@[�so�G���|w�vWϢZ<�8E�\�V'4�di7ӊ�P�v��x`����Q�ݤ��DA��Y1�z��V��t��
�Y����*d���h��%%�B���|�Y
`r��ښ=�+��	S���Vg��lq���w!J��̜w�Y�>(�U����c`��C��Qz�*����sP��7�U�Od�y.���H^�9��,͎���/頣	�}�;� >�c���|�W�Ep�_Ϯ\�Q���%� +��)$�Q ���A}��-M�V��u\;����Ȟ��^�-=8�}i:D�CC���/,���f�>����@ZV�.�*5����g{�%�޺�XY��9��97���Oz.�~>��x�D\���^� ��>��5D�*sD9��$>�a���82�t#��=����Xvu��W�o���
��4E���=P=w�����ڡ����ζ�����V�o�տH.��>�y��Sċ�=�^e<\�9^�@���T�T�~��g?�������8@3o��u#<�*��sz�(fhe3<�	x��@��F��M���P��, �ۤ�9�.������׋��H�؝ɑݻ|´�b����9�-��G��l��XԤ�Gs���i�l���|�o��4�<����t�����h��(C��l. a<st���b_�ܿ�o������?"F��zpq'��GE��US�Ɔ�,8��P���!������#q��Ij���{1<���N�D�E�)��������*�4�7�"]��|���7w�F�J%�l�w�%E�R{V�o���q��9.Q��q�sW9=;��A`���8��/I�*cGJ�H�TȤ_䩣�d�hO�1���Rtw�X<��QI�k� SȌ[y8����h 8�={d����i�> ?�/�%-�Z�>� t��{W~��̱���wi�V���,m�9���9��b�>P�4���?]�m�WX��:�O��c��6O�9^��,R�����笂$��6Q1��hf�iDH��{��ǡ#�K)܂=!�`iL%si�1�(���p���+"��.fkc3h�#<�mi���u�o��{M�k�Ik*o����$����gf ځ��*�Y֫sL	�9��+�B�`��7~��[Em����ZK��S�2�f@�!�1=��_��O�;ȅAΚׅt#�L��:C��I\!J�a�.J�ǹ~���|���t2����F���Ĺ<�ÑQ���T�wy�{��tf���pz���b���a�~p��!C%L�k9
�b�d�Y�VR�#&nδ@��^�A#;pc|��N��ּ���d�J�*�4�^&#������@t��t�f{F�2�G��CV���#���Z���nPZ���D�r�eP�z����Qs�'3�����v 	�e�-�^��,߀��>*��_	y%dq ��y���6A�uJ-
�
ͥͣ=9��#�KG�D}v%F�K�,G ���)=�]�#Qz��0p#�n��ɂ��U��@~J	���C#).$����Vv�Cσ�x�I��)ˢ�(�?@�`j״ZW�A�8�B���a׸�)��%��j���lAP<Z��C�K���
PW�ߎx�p')������_�!Є�,�������{z~�*��"'i>4���G���S��KנD�1�/p�^u�߼M��X�-%�V=�5h���3g&Y�r�?�X�΍��# ��ߟLc�ℰ`���A/6�d�ׯj���η�"����a�7��@S���1dH�5�k|w���4��.oi�`��^6g����DrP��,��m��P���.�Zk�� ��Sx�8U}&�7���2(���I�V�s�d���F�R���q�$X�����\�r>��#�R�{�a�5��٠�h$c�W�ӧ��j\{��hS�Ij��N�}����8���b<G�UV�����"U�s_�%R���A�z<H%�(U�S�
Zs[J���(��N�����,���`{�?�|��5��5h�QM�h�0��j6e�hR{�t��s�C�'�ڞ,{��(�C`;�ʤO�;�n۱��B+����8K����X��˧z�c��/DI�js�"�Z�e�?�~s��e�)c��FE]k�)a��C)o�,�	����R���w�b�v(�,|iϓg�/�� ���9"e��͏��UU���A7��ø���B��)c�KMG,����
6��¢��	��q�*�����3��e��+3�����t��A!>�+<1���m_�HN*���H��AB��Fr�����D�����5ۍw�ʚN�C@һ�m#��L�J\���Zߡ�YZ/�Zun�s�gk��i����/	 �8/��8g%�{g�#bJ"�k�`����;��q0����Ǹ��$���<�-�:���Wz��w�����\�s�!��)�%}�)�-�2g/����>U3�аJ�Z+'�%N�^������!��i��j��I«-�k`(�L^'��#X}�Ƿ�/I�I>Y��w\w"]3̴$_��~�t+E�]<���XcW)cO�G$��f�g̔g:�hC	����V�x�ԫ��!W����F'�N�D�L�D<�2*ADN6��Aa SYԥ����(&�	r8���ѵ����|��k�ݢ�-AQ��Hq���ڹ��)@}��)&�x��q%��7 �
� w���V�-���`N^�-�!-��X��!�%y!h���Ў	�ʏE;hiyB��Eܬo`�R�|�D��)Mrj����o�X���?� �$ ���c�H�%u3AN�9���٫X�ȼ��v�����ը�8L��7��X<Aؓ�J��sa�A�~߻�xՋ\���t�1��߾��4h��Җ��3A!��Y�=�?���"�S�/ZPS�������ˮ�2��O��ܘ/����<#���`����e�烉���n�L���tƷ�E�������Y��e,�8��ގ�.��#ZKY$��'F����P�[]K�iy�F �i�
�GY�1�Σ� Le4X�xE��Eu�o��!��]1��	VFtٻQ�+Ux�7���o���VUJv*�r<��0��)��49iF��i�p�G���c�d�wT����r�����A�h�s�n�7�x&�xrl�թ����a��^�޻��J�3E�{2o��P{���^���{w����)oK2ț޴�nF)dV)�G���Em�3��Uۭ�y@"応\��b�M'��3��$��u���]k@��3��ؚ�sJ��8]���E�HcM@����l��}{nB9�oY��y�6��@PO�,pzR0��:�L����oD�&��j��P�F��ӣ�8���W�4��d��7��D��fv��Ճ�ݎS'�]�w^.��|��>�|z}�7����g��Q�J$�f��UL��`D�.}#���X����[C`h���!I�Z�����㿨j��W�t���p�.�|��ūAz`rs٠�Ƀ�����*R@_�g�.1x�6�y#�o����,�>��Ѕ#ʉK�F© eZ�lG�8A���I� �ɜEE��V�4��zK��q���_�x�i:� �JhAp��ҭd�R:i�i�z��q�׾*����K2��Ԣ `Y�ܑr��Q��I��3�Ȝ�	VrSx��*���4+*v���u���E4�B*b�fTm��Ka�sI�͟21�{)׀���Ǆ�E��?3���}(O�K��XD�1���<�����p>���-�7�W�X̓B�:��c�|����~k~`sކ�g���},VX��љ�yqڅd�R����T0�.�{2�&� �OXֽa+���ߩ"��Q�T��C�4���,b;ZltmF@���InH9���sfmY�~��inuә���S>�q�AD���taw��I6��4��`�Kj]&0���D�y
36�� ���Fl�5����L]:dwQ��i�LP/��t��Nx0��%8�̱���6�k�E\B�G�����vN�W^r���0�v2�5D����Z|�=��N  >�K�s/��-#]Y"�FV�O~Y!���D�/^�4�q�G�]\b˄�x)#l�07�����º�oŅ�L�����3�^m+qu7�υ���q4��&��غ��/�K/Ⱦ(9Z���j^�Q5L�QE��?I	$��-`wҙ1�q�v�F��R)���wCB:>����?����Z�Rd$��_)	$	Ȁ]�1|�9�
4m3�-���\BCKs�\+��1�,��L�ZI�7�=�m����w��MC�0H�7��8r+��n& (1/dM�'H�5]�g�_��7��)cv�k�.�Լ2�b��a�3�;�������E��9���uθ��t�-��D[����Z���WǼ�Y��Z�Di7m5�������Yp�$�a`�=&'l#pX�=d����`7���
)Ƅ�?p#�oU)� �*���[�����)X��z�$蕒�Ȅ���n�k2�(�+�v�u�e(�El��Z��θa����^R��,1��@s�~(�ю���F�R�{��+�PPo�|�E�� f--�Q��Xw\��,���AE��7��ת���MW����3.,<���
s���8�U��E�DmfԋKQ��m5\���|
o8���W;�o-֍9�ɜ�F�F2X��(:~�N�7��lV����t7��5c�E��CӀ�,;��}7�Ĳ�߷kXٸz���:���`JJ=%���7��b��������f+A_ٝ���E�Y8�Ycz���9�*��L�U�������rA���d���GY�* vg��V"w��"���u�r��,"3���9�,�5:eY��|��!���k>��\_۽�hV�ι�x/�!��rP����Z�j�\��l�0�rT���;%I���ḳj�Zo�,K�³F� �4~E�&H�*[<-�Z�ž,���ô,���ú�;v��0�v���f�P��;XY�eo�S������s��BO���t�����.)?�B�O���S;D��ķ��f�Ü]È�����T���<�3�8��ٲ�c=j���! l�(E�R���Ĕ�#L�	a�o��8G
>SH�^��0��9�:�@�:%��y�8��ja���9�� ��:|�����M+�oJʢX�09����X�&��W�ؕ׸��}��3�8DNYB<�mل'n»>􂫔b-��݆�I��٨���OU�{���$y��y;r0���K��[_1ʰk��	��%0;����K�S���(�~�~��</?c�s#��S�_v8��Z)�)ڕ��YS��/u�g�f�1�PIOH�2ۻ��J��V�-���p
���.�CXG`�]Z��
%�F�	L~��x`wXp�2K��d�V���g��K�H�	��1��&O���>&��#���l��m�� ��f$p�]��ؖ���*�8��1�F����{[���D�hr��>�Q�2�k� >	)�Y�a�#ev[�H�9�c������c9!q���xiq[�CT ���k��4�X��Q�J_b�W��r��륈v�w@D@�n���&�N��v �'kʱ8k�UC�*@�p�w���p��y/��� �bu3])v�A�fiH�m�dO�|�ЫN�"y*���z�����XX���Y�� F��+u/P�Ԥ�&A;��D�[}�lN�ʣ&�r�D��N�J��o\��VM�la$3S�GS�:i�^8ɓ��Z4�p�> Gp~�8�Y۽{K��o�:�=q�_T��PaV�#�zD��R����:��#�P��`͏���Y{Ӷ�x�����K~Հ �c*��V��^O��_��7�5�������!���.��B߰$=$=`Z���ڀg$)���*��¬c����Z�Id��f�\��rM�?�
��� N�}o���t��b� s����i�����	���wsō.�M.,v9�k1HO����\`|X���&���q	�w]�Pb�I��;��ۄ@�0�6�������Hg�(����0�_>��f��ۇ��ʂl��
mo����{KF^��v�.F��wޜ�x��)~}�bj������`����*�ޞ
o0|i�֥���6<�S�K߾���r���%z�q7R^ZW{�E�D�Q!f�s�S
L<N9�NA�M���:x�^������&��o[�S�c�S`��}L�P;|mY�H:%���e�D��'�"� �IN>�cl�`��J+�FNp7�-5;�/��
������d@z9�-��߆h��:�1�3�:����Ֆ�5w��h�z^� �_a�'K�SS>#T�D�� ��n.����G�)�q�Q��b'Z�Ȁ��ђ��R߄����>Jң�9����I�s1����h�%�[�W��KQA�1�W���􌚅҉^!�'6o>���M/���ց����'^�l`T�m�A��WN��p���М�k�JJX���	���c�埵э����A�ר���f���]@�=~��X�e��B�2���v�}�8�V��j8bZ+v��S9d>�S.��2���W��Eی��0���s��=P.t���Cf9ѭ&*�4� ��/��jxB��I�u��Y�e�b	L�>��;�������8��p���S���0`��k��G�Q5Z���؆|}֋�d��8��Ͻ�vP)W�pc"�Bpp��>]I!���m��s�q¨�VH��;�MǴPi0nQ6uh��6�t��:[�����ԋ`J�(�s���H�%�z���w��ZEG��F%r!7������e�\�zge��
*�=$��*��	cH�mf*I@5a��&V��k���DrO��B����r�蟾P�v�V-s��r�фU�~�+��)a�%Lu~��x݌��@ $��jw�N����(Ms�B��=Vp�����u���A�Q� ߁4�y<x��Q �ފ ��$��c#��HBR˦���y�rf�,�D��b~��^^�ƦDy����#aG��ucw�F��1�E��>c��lm�����=t���}R�3upd�Wy�<A8���z�J>M��q�Z	�G>����=ye25���75:T4[�uR�D�^�}1�R[����gne�����W��|#��L~�Ezk;���Vw��*۳$i��6&�M{���Ol��1�*��}?4nD4��d5ߌ?�C��9�]f���B�%�V��&��1�b9J�p!~����>;c�E['i�߰*0I�	9��a«��ia�䗙���v,�̧G��s�;��X��Ĳ(���Zc|�bd>����\W��H�\����*�ΈW��Qh�A��,@A#��L�A�b�r���zZ	�B/h����nc�,���kֶ%��WI?#E0"A��z���ޑ�<?}�Mt��I��qա+�xZG�GU^}�qd��i���6�?���v�5\cia]m�o��79h>k��cZ5�V�tDJ!���!s�XJ
wdb#�Tg�{~���[J��X�у�M,���!o��:�:-I�c�@(Ƞ�[�	�o	c��41���3��dО�f�jL�p�L0�mݱ�a<��O���uz�����E#2����k�M+�Y��L���C:�D�O�4�V �&��g�r��Ӛ�5¼X�ȶ��gbu��t<�Ɍ�~e�愑������;�֋UzAX����wMÖ��e&����˥�o���K�H�BzĤ���_枉�?�[��E��s���^l{t�Ɯ�v�'#5��X�Bx4Y�)�]̈́�x�$l��dI+sp��$��K�de�x�>
���m6�>7�Ԗ�^��B)�?ٍk����o�����]��k^��R��y��|2���\�$YP�n��J�?�K�MM����u{fc#[��j�ҿ�v:|�:ȡ綃��?��'FQf��w�Eo���&R��U��8o{��I�`|�*�N�Psl�WZ��8�A�$��:wȈ��aV��@�t��C=�-u���7Z+�V��eK��+��b��/�&A��־�r���>q:�^�W�M{�<�{���8b�%< �ݒ<;L�uE��ŬDt��B�|� �H��9� ��.����W�߂�� �t9� iLW[��*���-a�X =��L`
\y��7 �*�-V���Rz�Έ���� �����3��A�K���"1(Ȏ�s�����wngF�(z��MQo�¼�������
��I�Q�U/>�3�M�p�0�+�c�E�G��dT:3O+Uْ���f�(I*�1�jM8��c�>o3thXA�b��Ѥ�";�/��C�cm�����^����Gn�����,A��[��2��Q9���Q�q ��Y�)=r�e[�ZKf_y�T�i@-rT��j���Se�cZ0Qx?�R��%��Hܽ42���ӣX�����9ǯ�1�������;�ܯ��0|��dJ�`_1��ʱC,�+�6\��WxEsl�v<x������������>x2K�fGF��ǳ���F�
�j�D��.#���f=d�_T��6��6����<D/QyG&����tf�q������y��j$�P�b�*��>/�`! ��UT�8yL�B
��=����_Hд�{��
�d��j`@�}�9M^I6�s͝�$��Iѳ���!TD����Hx�˷\-:��7,#3ب��i�{��]n:	����٪퍌�R�p	�qI)�eO����H6�������'KA:�:��f��
��jHB�ZUg��
&	v��q�gl��?%Q���$m֙ ,��_;_x�B��1��MT��Yvs�aO�ȪGT.	'Z����f�����F~RB���V��"쥍Z@
�y}m�?ښ���-*�|lu�H�'x:+:�}��_�p�D,aE��&*�[�p�G�"��b�0�Dˣ�A,�J�7�ۼ�Dv�}&��<uB�Mʁ++̈����?��!�@]ybm�d�&�0���})��Þ�aC�����_�B��υi����ytK��U�{E{��|�)vnd�	y`7�����a�38QϊW���NC�l�KpCN��6�HbMI�J�@Z��#>���m�� �I�(%�u��O�j �G���qKE���Y�㵓% vt���|o��I)�� �< �=H��8f��� ?�0��&3	AVޞL��C�"3�u����D��`òQ���ކ_j�������`���8d��1k�4��/$	�ܝt�tdny��}����I��B1���]Q5�qG�_h$qBq�=�����[_�����W���'�Bz�b�16�j�� �B=�*X��!�w�.1ɖ1�"�`�����<i��qZ��`��9��n��k'f����^�;��DRu�Av��,���f�|�ʧ�H�|G�2S�X���Ih�Q���ER�)|�����
{���
�fq'���Hz�!6h~���Ad�8��]�34��|*�����1��1ᙞ����t���n�B��-�a���-����\�X���m���[k�ud\(:�|�0�����}NcO�y� �a<n�ʔ�UL�w[����.���f&�r�.��B���Tn�]�q�,�<�[���p;I�j�	���'�T6�S�z��z���|h?Y�mU\֎N�e��,�6W���RG��vD���_�v��:�i�:6Ԏ��L:v͍�Ӟ������ԥ_ʧK�YV{�;w�g��'�h��
�y�����3�D��i��'Z�A��P1�QK�T�����\ /�e��ZR��i�G���3>ź�����t�2����?C\1�'��d���.��zA}�j@BQ�2.o6��7�H��̗��F�YJU�br�0=���O ��C<f��&o¯<��L	b237�Q���V(m�h�j��o�0�aÆ>�4�O9�/9 +nk�)�L!�m�u�H������q�1I-�7�;��z��:$��PI����~.��9�3��Gpމ]&�Y2�)L���բ�*��~�l�C)�M_I#��/�3u�]�D��k�Q��:9l��_+��<	���o�mn�X=�R�A�iz<�������ɎM�?/F5�t��^g�@�����ݧ�M�_�3x�[B�W'����kT�p,1��;n��x���.��<-r����Z��XO^b�\[z���b|Zf���`��r�����^��2n��.in��*E^-Q�;&P����(Q��ro	��9C�5����2\3� O++#,j2,�c����AZ�t�;H��Y���J2N�3:,
ni��f'2���3:c�LV��v���xIjٜQ���J��`�}�x���ݢ������v<��8c�洎�5I�������n/�NɜQ�8����b��I�&�wj�+�
N������rSmE��Q�φ���6+JU��箔W�F�Ѽ���R��Z�u؅mM�����0�D߃=��m��c%���;�]Y7��q���C:$)�`�m������a8Vˎ��E�^M�yx�$��L��U&��8�;^$?9u)"�+��ǽQ@tR9�������XE���!J;�#PGl{���&,�| 0WJ�� 	���Y<�e� ������D��O��q+4�|���Y�Я[�~u�Z�67�z#��v�`�;2`v7b��r,sgq�����G���F
Ε���̰	�AaQ��捠���Q��.ʜ�[.�jE�(��?�?|{��N�pk+��)���?���L3E-��u��!�zo�����5d�',��Dc�5�6���z �6��e3hs<=�vTd����~3������躕����/e�U����
6��k�x�]�Cbf�1-�Źa4˭��'p=]��j��۶H���/���Iگ�HM����J��b�oD�f0���^���r���*�����*ҷ�������U����MCz�it�����4Y,4�B�62���ۧ�QteC�ږ<]ͦ�0 �00q��l��ۺ'Q�v+���G�X��"
lf�_���S�f6ŗ�?S)�L��K�9��"��c��p+j'�����xI�����j4��{����J�n���*dl�c�$��{��OxIC�&��1�)�C?uI�-@�Z�#����S�ʢ"�ɸ� ���ݺ��7������-���_���C3C��\���m�����'��ٟ��a0�����e�^�t��\q
�������oĪ���W9Y�iQ�Ճ����X���XV�ݣΑ���i`��"$��L�~c����`��>�Z�0�ːl�V�_Me?��?7 F��-��X �(6���0)s>�������o<L�&�c[�_`�%)H�|ߋH�U�pG����)^'��X����^��Cp��h<���/Mu���5��M%8�q�T��=&�Š�]p.�M�r��B �T~�C@��#�Ȉ�V�Ds2&�뼎:��W#��X�g6C69qa��-�	m�P����j�ϧb=}	�����Q9�'�?��,m�©N9ռ��σ
��Ĩ�
�y����cc5��Tdfx(b�?�N�\�9���d���r�EP�D���;��Σ_r���I:���~Y���4�����Md����#���2�J20��z芣�@w3tG=�$��c������V�+��3���X����%}��{Z��)���EO��y�k_�%�\7��0a{dJ�W���F�-��x�T����Ɋc�9�M����ʗ�@��Ҷ�siB��lF���%�,O�o�]�/�l����Fߧ�8нN�*�W��	M�ٓڟq
"�N�_P��h!�ab;sR+�5h�n���H�B��~�L��/�Y��K��6�)�L��d:8�j�c�1�Z�XC`[����mK�n����<Qt�Y����vy��'��BBx��]��enhSSײ��oLg@�S-�K/����`R��b��|P'�H"0�2h�Tu.ԙ|p3�Mj��,M�d�QG63r�9>U�P+>�^�q�!<)�hr�\dU��W��V���V��o	�t�c�b���$����L*�r%�_bh���
XျӚ�ِ�^I�lH�|��A`���8�?|*�W��\E�.%<7�k���n`����*QE�	K�]�]���DSt/�w���É=%��_�=◕뵘����'3Pu<Bl'⪥%ک '�8#ߪd,ǸoF���w��7�K|���1fz��[2&���w�f�HS����OJ��g�w� �ڭ��*L�$��)ר���;xg�����g�c�,���%%̿h"J���T��U)˺E��tl���p7�N�D�ݰi�+t�����Ɲ�\C��;1�6��˯����W��ೊ�����t�Ǟ#��dPb��$���H��_�z���KI VTb=]�n2Y�huo;?�v��W�14;��InA��*>�n�LΗS�HN��̗� &v�>F��`2G�L�/կ�Z-p�_+"a�LN�2Iu�f�����ݿE�q���5��듃o�ĉ=�@�P�\�O�~�0��fR(��t���Ig�a�!ow��Z0j)�0a5C��tp�]^! 7�F����|�dbgJ`"��Vw�����Jf?��X���*�Xf����"�S"���at�C�U�]r���6�R�qj�$�x/^#g�M����jr~�b�s޶[�%D�)8�w �ʀ�V[Km�����dz��]��������В.�T$:ݙ�}�-�'�Qqq߃�}2�B��ʝ�ҁ\�Hjn�q�=IN����J� �g�!����Q�~��q�ϒJ˂��H�Y2�wyv��M"]����Cݓ5�!K��|x��4)ԣ�5�� �v�7v� �����R`o���}���J<����������3��8�B�G�y�߾h���h���{�2O�����YRiD�����))F����u2��f���d=���sv���	�
m�m�z��Wz�F!꧱���q;��0a��m�]IP����r��L��O��S�zwu�.�pb�x���Nh�Hq	�I��xd��ǣX��������?��G�6�h��$���R�LR=�ܪ�ry��&�3 �����3tr�!N�v�xD"ZC���ܐ��[��6i�6;��/���z� ��@Q����,`|�����8q�%'��p xc3UC@�����X�?x��I1W���)�w��m�ص��`����6$#�d�QY��|o��	�'������կ���IZT�m����aV�9,s�m�Xr,�2�6ױ��Ԓ�w9"?Ij��:�(��{
ǫy����61��㕥�>�qvqW��s\Y��������Z5����y\W�Ȏ��V���f��5���O�CK�RE,����p������&��e9v���7��@�t����|b	 A���W�s� 7�uK���+�Ϗ��C���q��L򟎯���>"��7�i���P�=�U@��IʴRƑ�u6�@*Ejg]D1�J5��x�BS�`�W��!E���a�����8l5�Kc��Zu1�:t5�ֱ�~���B���J˰��9A�%a#�$.ݒg�~~�a�W��}��`����Nu�5)�H��gd����&����ɾ��%w)[e$E> C2���˳��;��h��"�"`��Da�0���ߕHT7�*g[M0n.m��` ��a��9N$�U� ��c�>���.a��&��qTp� Q�#)�Ԍ ��3u��#�Y�C�n
(SH!WV���I<�������~seU몬>؄x����!v#�<@X�cqnnՆV����]ݝk�Ax�U���6�Q�$�/��R	_�c�@�Y"�O�p��n�݆��۝*��*9�� T;�}�?mh��O;t�}��t�s�X3�������nqhNH�dK&i�I�����_<�N�����IV%��3K�&��=�CDDΨ�u{5�e�{����:�%lK���3l ��(��i֏�� U]����W��v��]\�������.H�|��G���C�-��g`�%>&���$ ӿ�l}�C�<�ȣ�	i��&U^���Z���^N@|�ٙ����@I���cjJu�
�VL<�qc�f�W�ߨy�VUU�z�}�O�#�^u&pUbһ�j�a�M;{��^��U���эɻm�i��������DP�i�����7<��yJ�^�ԝ��:',�+S��~��.+��S)�)q~'sd�Y�I���}�m����g]�T�XCD����n�1�2�$l�!t�v�%d�imo�=��`����6BN�1!ZV+�l��:��\�"j�3ٺ�T�r���ȥ���At�#�8�ȈA-P�B��D�&����p��L�*���p��B��!�1��ŵ^�\��o����{"4�>yH�ir��KW�&�Y�Ù�������2�*́/�<=�w_�rb�zdao�q�A�ɰ��T$yN���4��t���&����F��y�Q���>n���hfX
pt�-�p�@k0B���Ȧ�[����R�B#���]|Qys�P�����=�urRS{�sv�4�L���t�����rN٫�]��Y�u��3�o�	�7̴���
ws[����. �#��LX3r���<`QGn�@�쏆WR�#�����9��dp��m3υm�� �G|�=��G��� P_p�ȷ����V��Ԫ�>����a#d�y��%�OV��%�|#�"vڭ%��������O]�ђ�c���LZ�� ����� N~S��F���)040��vvt�M�iJ3�$]'���l��p� �gd~�`y��&Xj�Kh�����%_
>��Y�^����^��Y�51�t�O-J?�>�ES�i��ܘ�s9�NE�p��#��[��1�%��μ�B%)����q�h���HN�缛�=W�=���FOz�}����z�CI/�91��+[4�ڂ�>��7�M*������3��!�Z2,���ݮ���wo��T��&�P�����効0)� F��8��&��B!Fѽg
M��)�B����Km<���ͬW�JE�e1��_��f={E�$d>FB�q%�[�:�L�AP
�~��z�u��5U���h��ƚI��z������f�h�}n�tWÅ�!LT`���f,.\m�����p#�'x~���Xc\�F��P��u+�!�Ǘc�9������^Y�ȨB*�z{��[n�����'�y�8����9���h�b�wx{|�������n�&�7��U{|�M���qH�s�ɞGݬU^a��S��r�9�y�G�>�������y9�]�-�S"U>W���,�tW��`aq�R��������]������^})�~ ТC�Mt� ��`�\�X��8��!�`y<�rf>�k0�{<,�{�L��;/����Tۆ�u,�P�e�gC�C%�bi��^��hz�l���h�ۭ��O/��kIbuN�����党�Jf^��7�i�:$�%�]�m�Ѩ����.9�Q�IBf�cda���62b�̚����?�q{[<�x`��ud)!��"<���X/~4\�JJ��f�	���F�O#H�9f�M���{�;�%�quHv�mƁ�,!k�p2S�����a
JP~�f�&,��5=�������A�Iei������_:$ �-p\��L�+
����̰ډ_�e_T���r	k�QA~�|.�M�Sv��5���Z�!.�ބ+���=�� �a9f�E�vqn�%S�*��cQ�rJ=T6�][>���j3�Zۘ#��D��,H3���$k��χL��}+&_��&@�ř��H>y����Ր�@Lh���=��{�_wmS�����i����q��:`�Y�$Kb q��v��z��i�j�� ��
�ly���X�����$n�*o}�\h�S2I"�fB�]l�g��tH��A2�e2EP����i?�3/2s�d6�'��:�1������~7"�1+5�<Ƴ�#�@���E�/�-����9�|���+3(�;Mcy�=3��Tvq�EB�'�6�}!%�")}��q���{ؼ��	 AtQ#��t��8@S���}U�UC�W_��G*1?��V���<��û:V�w��ȌA�����)�f�8U�E`������j$�/�E��	{�k�o�g�?[��ێ��_�L:U�d��Ɵ=�v-�
x�zhA����(%��	� ��Uѥ%2
4Zw]�G���g�Y�[R(�/Pd�"� o� z���C֭�v�"t�>�̨?��Է�\䋮����EĀ-@���|��Y�������������IbTi���>7��e�e�]��LiX+��-���{�1x@3G����Pv&^ڝ��0�s?w	�jx�����ѫj�8�J�[���y~ﳙ�V\t�[_���U@+b��}���1�����?��02ʵ�Ph$^�'�r&�FD���{)`���PD_��e��8.)�����WO�.���"�i8��Ⱞj���,���hx2!>�a;�~�W��[�n$U����g�.8��ـ@IÝ�v7'[����kJ&� �QWU�=�r���e�sp��CO��S&����Ix�Ĳ	��U,e/�`�N��+�O���&�K�{�6��ދ}Q����NDަ����OX�@k6>W���8*�1�(��,��D� ����;D���T)�
V�@�|C=ƀ��n�ֳ�g��IW��2aA	�v���K!|<0��H���;c��W][DDFD�Q�
��ގ���k��t���0��g1kDGe�q)0P�f�I\#_���q��hqʸ'�{\PU[V�ʩ�D�J���z+��[/&�ͭi;��x�d�Iq�&���M�ʇ����Z����Y홦���cǳ���!�}�n2�̐)/<��+��a �?7�R}�=�&V�d�{��hWK��j7dW�,�-�g�;h��.qVd��UZ��G�$Le�QHB$\xħ�+`'�k��?��?R���b�5�T��A<�b��Eh�=�J6?�c���[�G�ףX��X~���GRa���,�����5ai?���/���J�n��"_��<Rj�%����Rճ��bV��鈒��f��פAh��,����	v%3+"��(*"4�}�rN�z���s!�[^��B,��E����Lͤo`ׁj!�_�O�|��ei�Q��	]t�	�Z���f�c��o�j꟦�Qѩ��ŵZf�`T�>�`:"�����M�Yr���wH��eu��n4�|W�\(�j��ќD��Hb���a�l-��B2�.�V�W��ڜ��[�}��rC!#����/�Y�ƽ�ɐ(�:P�#���3�����	���������t���OO�E �9�^�[�tC�%���*��E�<���J[�k��il��v':�i�v-l�j�uQ���s:{�	�g��٪Rm�?�F纉k[j�n�5)N0u�Xr��b�n���섨�M���۴T��?^kB����D�Z��3�8QcMp�x��\3 �9��OO�o�XECז0�s�|0z��=�.H�?fhNW��%�K�\Tn/_���ں���ܗ��j��)7�#���9V�[�r�[]�%�dr6�;�ɝS��قǧqh|���.�A���!��9�T��>9�O#9���C�f�?�uX6J\g%��8`j.��ݐ�w3J�
o\&�F��=:��|��Cq%*�
��C�J���6?2�F3�a���lJ�_�%:M�D����f�
��$=C˱�P��|�fje[�b�%��y� $]��sED@��n�QQ��:��yM0�N�j�
�-�L�G��+��s��n�9�ʤ�����G���� ھ�qs��n�H��VM�wt�@������[P�$��Lپ딞���K,�d�b��v�M%�l�3z7@�.T+�ki�^Nԑ�rFYS��v(�q��!ǉ8�R͝�"���5?�s�r@l��Z>���G�3���^\.���eK��(�3��=���*]���m�#=�9o�/����"�8#5��?.A�80BhLz;<G�&<9#`=�2����^ �x�s����b�:#���?+I�m�@u1��,+m��Nj���ߟ�M�L��K+�Z��-�����ԣ9©�<-9^C�Q�{M7`�p���挽��H����9�f�)�I≭y����nF�n.����Y������%t^2�0�.���T�ݹc�^�?!8�I���{�<�����$
�g���<l��=�4��8J�^M��\|uA��	B�c�(�?��/�D�U�vK��!����g��i�:�9$ L
�ˁ�*b�.��i�o�"Ξp���?��VJ;J�0:��i\�F���.(���uL�N֝�M����m��뿕�8�*j�k�����-b�r8x�]���6��.�I��� �Y(r�L����ETe\mЁ�ު���Ml{6��	\6���x,%�B��qW<w�4ٔ�(�߰>�SIc�P�j�S���2�?��

�a�'�;����e%]�����2�r��?T�M�2/`Y�n��Ԉ���_�Sg7��Έ�g��=��p���i�������f�Ƶ7~=���P齞L�SڮA �jӮW�����]��|^�A�$��L6��	�Q�7&2�j��gE��EE���C��Ͳ&$�D_���q^�1��n�B���p��pT/B��E;s��܌�h?@��:�A:�:@i��	�ӓ���xaD@�K��.�������'Euy����	J��7���#)�,�YTVh�������߷�B����>m��G.	�g�*�rht%H*Q3�g,�2G�As�5�L�_,$`)�_���S���[�Vy���!A�xN��⯙���np� ��>�]�w�)<�֫���rc�u�mY������i�s�ò	R���sm0/�c�@(.V���d��wY��n�|?���8ӀT����%T�$`��쬪�h�!W�a�#T~1S�p�S^!"�GP�?4K�D�A�V$�0���t��i�4�ʤ$�U_O��u%$��?�%���/�����$���)��vI�n�v�b�#���M���o����r_��q��D�;�&�a����XC���l�st�ާ���ڲ�G�8>�s-�����"nxO��Ex 	���e|�w[u��e��3Ӯ?`hd#0~9Ǌ�Թ1ň.Dt����$-��W���;{����JQj(
�Kf]E�T��q|���D��w��� �������,��^{"���ZHdU�l�*�E��~��c! 5�{_>��J�^~�UW\qc��4yD�/EC�M�U�h�(���k�J��w[^�R�Z�T�8���W�J	t~��:���Ybb�
.ؘ�g*s�&����Ke�>�J;�)���l�bgSj�`8��gT��:��T��WL���=��v�� ��*:Y:��`���.o�#��v��,N���~yȻ'�pSH&>�3�Uex] 	'�yP�6Ɛ|���p�H.Fj��M�#�Y!˥(�Q����!+�3Θp�����j�O��ي�z�q�����2�NKV��In`�|*z�^.��6��v\~e�(�|�Op�Q}=�mrG8��@>�8��g�o��T:�GVT.HLK����K���X��(��"#�IصE$���	E�-�
�?�����%�v
ȳ��l}<%�@=:�lx�gl�'g��A�B�rU9�9p��A��>��d6�]����6��Ɉ�,ao*�����<|i��Ժ��}��cɈ6�G1@-�O���H5��,9�Hvd.�M��Pa�j�+�Ƴtc!���� ,��B���]�pi4o��z��5&�1FO4����\��&�<_H�M5M���Q���n Ό��*��k�TD~�����O衢~<lp�����M���y�b�!m�]����� G)~ߎ�t[NT_���z��|.�1�Be>\x��'!�\ǁ�4�@�[����>��� H�8L�=a����e6/��|���{)�q�Ռ�=��ˎ�#
�:���eZ�9�E:�Ո�{���7���Ѯ0�c5)�y��	B5;��%��S|cDvGpc
�8K=Kr��HǕ@�R���6�e��g�.������4F ��z�m�FL��sF����6P���x5�4���<Q����+��ʵ�)r�e�� �FP1 D�k��5_��#��t�xi&�(�5�{X[v�V�i���i{ٞG���k�c�����H���L=�(����[IM4�V�h�9��Io)����:Թ@�z�Z!���_yV#'�4r�@�#Z�� �$&1N�S�)�����w��Ք���e ,��]D���t��4�9���S�[�R���� 9�_|L`�,wr%���gh�V3}�#zz�	ڤ>@�茝�v�t�DPְ:�Ѷ�k<�z�}<j>�ף5z�e�d�:��޽��鄿iKn�8��K�σPN:�0�C�,�4����d��-kv������;��rV�=�P�{ҫ�J'�������qp�#4јH�8Y�\�U��#6U����N�O��`&�u�|��-��3�1)�����X'�:u��Z ,�6p�D��Э����Lp���͜�]@k:���[���m��xg�ב�Oâb'�$�֎����A��NnkY{��1�g�z��Y���Ny�l�Z�5�l���d� �v�ET������t5ԙ�O�����/1���Y���q���i� �P7��������':��}��,��,�2����V�jTŕ2"�[�04����ڱ!T�u�i��n٢��m���	c����B�/���B����e~��F>�W���?]�	�`����!X�b�#�&|��d��]6��9��;d�*u�T�U �����pi1��B�M]��T�*Ti���qLX�M,��p��>���*���_!1Η����L�khj	I�ڵ4X�=$���p��c�;C� �o�8����Y9�	���d(Jr(x!'�\I�}�q�� ��5�����͑ʝ2�0N��N ;78��C�$�ES�L^ �^��|�E<�9jn%����(��ݾ��7e$�û�0b�k_Yƹ:�7ȓ��ӲصC
xig`���5tj 5�{�Gv�X.'���V�t�Z���g�~�P�z�5���i���訯��:�����w��6�i�Zt�3 ��"gf:�pJY*��#~�φT�&Ǉ]u�Ǡ��;���
�w��'������Cӽbƥ� ��r*L�v���ȟP���L`� `X���}ޡ��Y�Gk�3�5
��o��>_a�R�a`������"�}�%�:�	�� Vb���?\V�G�w
a���&�/vJ���5�p���h�H+�B��O�9��=���A�}��L�l	�g�'Å�[Fo<
^���x�H���b'<ߦv��Kob2
��)!�pu�p8;e��?�Dp@��ijRA;�F�Kʩ'�lgڻ!���4�ձ%��B)��e����h�ct�]���Z��ɾ7���<�b/�3Cq��pC�?^=V�7<��#�����h5;�3������.-�G6mL���ֺ�����f�fE�T�¿��L��Ʈ�b��$�<����~�3�ֈ�'݄�֭&�Z��k��`�Լ{�F�@, ���Q�hd�9u��GFv���0eD�>h�L@��zom<c�^�����'���pט��)�am]��P��>�b%]��@AE�ȶ�_���+�z� |烋��:<#��@�w���p��e�}��n޹�%��i�w*1~Rd̝�f	��>���]��� ���Mx��y�`�h��2� �?c�
暤��M�|����۟V���">����	<q�o8N�ZW�8X&����FT7�I 8@��$F�4O�gz��>h`oX�+�b���<H�:5�q��TR}u���y%�:��k��|���{�w^P0�|�@d_PT���/�MDh����5��%qjf�E������."m�.$(�/��a�L��7Fs�3oD�0��=/1�+�2�%$��'������!j&R2n�
�K����\ğyȊ��/Yy����Z��N g�	��J[H�6��ˍ!y�j��#��]*��ٰ�L��.�+����ż��r+L�:���G�{W/�\ q�w� �f���j2L��w=}[�����q@f�h$�L:�C6�����^��$�2ŉ�5U�M��6�X�RM'@���;�����T55#�8���dύ��A���޿.�5�h|�V���^�֑�(.�~��W�+�E}�&5�C�bԭɂKS��<��
�I�B� PK��o�2�%�Z&��>�Sn�=�z�wG���ܱlQʇn�ϕ�>�e�+l�|�Zw|S���N������s���~��5_�U�E���E%���k��]�c�a����d��D���/+=	���خy���vg��l�Z#�ZQ�掫� dÝ/ZD9�b�
����i>���7���
PTʫ�P�G �r{F��IbTu�A[���f�1o>��8���
/�8�-�Ж)��1���
���<<�P�h�u9i�,�r�t�(l0����>sbFdL� �is�Θp�M��s���?�0����Z����]F�J����Ǿ�v��ݎ:���6��6�)2�����J�lc�2�@˨3�6o�M� ���u�9e��)&��>�V�)��%�4t#p�Mo~ s��Ơ߬HE���+�4Xݝ�hɑr���;���Iv+?��T�cq8=�����2��aZ�*�f�
;�!��c����?n�+%�q�=���R-��/Q��l��I��u����?��0�6�NvtXH�4��/�1�;�/�rv�ڇ!���ƁZjS�q�I�@��3��E�%\%s�~靯F}�_x"�v\"}�	��i$�I(z�u���B�.'��.<��i�����p�#�����@P��a-�c"����e`�����_�]c	.aD~&8%�܊���WT�g��U�T�P	
m_.��Z޴m��;��4��[xb:�N3ӆ�
*f���lp�M+��y5YN�A'��o��$ɶ<�#�iVo�HA=0�\ı�x����6�{��'�)���#j;2я�Iliܷy�x<̕��r��י�TϵĔ3OF�Լ� T��&h�%�K�̣�G֐f����oiY`����Jk4�*|�*�Qn��E�1�M��N����_�lxE�/ܡ#l�w獫��q�s;���Y�=�Ĕ��n��lbZ�B'�<���ڲ�.�V��t����62�ɴr=�8��Ô<K�`���/ʽ/��t&U!D�c�[�y�f�����w���K��_�^j�J�$��o��= Y�Y��~�u N[xh���7�5� �Y��[�S�.�\�id�áY\y���H��L�=0�#�v�4��ue��*�6�	�YY�_е��UN#�Q���`{�QS,7�D]�;�nx��1'y��m4��s�5�-3m<vѓ�������!�2	�+f�#�ё\A�)�oy�렣�������
���Z��c��E����+2
���m
z͚sĸa ���Qe��ЖW��h�kJ�cBk�o�4�#�]4�+<:�N���M%R���n�`�_�e��8�^ �D	�BO�;$u+:`mn;ap�/ ���:�K<�/�Tn0C�ѿ��Z�uN~q��/ᳳ{�����Eb3#Fo^���
i<@%G�$���o�Eڦ f@�F ]+6|
�"X���r�b�e�� q��7�2,g9�yzN1T��$%H"��AŦo��&)k���h]����YK��$W���l<1�6�(�L󏹾�zҺj�����#�Cb�!�Қ/|��b�x��H�N�|�2h�K���"�ybr-ws4L*�ʗ����.ݮh>e�
��׽����kB��Ĩ
ho{:bX0k�F�-��{��b�9N�Ener|��^Ԗ�Vx�d���8H�`��B�5'���e�y��
v���w����1aQ�ee`�p��1'���1W<����c�t�k�'f���Qؔn�!|[	��D[5����㨆��k��(�%[��`{����U��X�4�N��	{�N:�/A��W"ᧈɳ;a���9�Z�ƞ�$l�4
v�x�(�Q�K`��j��6||)�C�B1$�Q��;�^�0�W�]u8�� ���i�0Q��u÷�5uV뛶6��O�A�a���M���]n�`�O\ju!�//\s�&ް�b"q�rƒ&���1�]��-���m�LS��m(��
���kYm7�V�Eʺ����Y������%���#6�D*������y�ӉP
�n��j�������p�F�)`x̢�!�'0%?�<$f~ؕ|Fe�ۼo]B�f|�2�$��}ʻ>��TmA5�(��!��EN5fn-u1��>��3��xC�$�Ҝ R$R���t�!؈p��ʅY
[�p�i}F�������(]�W������s���$"������vI�������A���&O�.x8��Í�*�|=T�tf�`���J8�ޖ��y�n�զ �L��1�?4�]�Cn�����K݋�H2���#������d����m�=�h�K5wx�܊���ĸ�O��k������_�^c�� &z�U�o�p~
4��-�U?��Y�> ���9���S��wJ�V�	S�Kk�5{M�1����1EL|KK�;wP*b��YU�׼��J��M/~���/�p��.��y��
/�0�El�%�Q\q���ǚ
��~w;�y����6�g� ���;b�\��{��L�����ۦ��\ܚ��R]���.U|��"�ǿ�k�5�%��X��C�&kq����E�s������E�S��٨��	ۤeR��)T�a ��:X^�1wed9�oD,��wF-����uN����ɏ�Q~�R�u4��V�L|'��bJ#�_r�+&"L�AMc&�%vh1֞3���pJ��i��M��,b�����LH�C	<Nȁ�ߘ}�>Æx���K�6��e͟��B�y�>;�),z}k���LVԽԬ7)��3�ŵB*1;?y�N��a��0������bROʉK�𠭵C����0b��v�sŬX��;�����R�Ȑ먒$�ך�H��#�=��K�"�Q�?C��o��!�̻�J�>�:'��Xqw5)�n�
��6D�D�����́�����].9(��=	2�Y�[�H�n(�:~3KZ"loqMXL�gM�9�}�t��Ph�ٚ���A�7����8�����Pxwq���1�1#1�[��N�����_aˆ�#^$Pu^$k��>�҅�(�tj�0D����/�D!��N�
�Y��w�ÜB��Jֱ���p�b�-�lH��~�EK-��K(�N�Y�,�m�18G�l�q�Z��.c�A��� �z����X��sR��Cvw�|t��S��cP��ES�xZ���v/�9U�v~���Rc�%����H�uf��f�kL_�|+&R�TK�����'bI��kм�h���.l�Cb�Q���7�!H:^���J�iAVX��'��-�-��	zZ��_xc\���13�B�g_�����C𑲊�[) �P	U*8[����fk�h�<�g��R2������@O��a��^�g������
�٬��SCTCmG�E��fT��o���g�2�K� ����u{B�jn�q���!�� ���4�\�aڮ�Ҧ%�)��c����kpZ'\�s�#�=��6�A��/6޾�I�Tshgد��g�EtWh�"��߬�m P9���9?Lq 9��Yxx����G&�����k��Q��`�<�F�����G�H��K�E-��<� �W�~tH?�OŞRd8��x�G��S�æ��˦9�V��qmY9AC�d�T�S�g�"@��{�ϑ�|6�Z���(���nL��al� �F@d�f�xMU(�`%;_�&�+�H�K�B�-1�]l��24u��o�k�\�dN/��h�z(?16qy�J�L>��S[���t"q;�g���oz1��ul1������HZ��{�[M�Y�2�Cք� ��l�@z2Vǣ��^��x�-�9!dO���� ڛ�.dgQG%��i�.���@m��� ��2:��V��Z���Q�?�p�����-��g�����:I���)��,uXr�����ݧ�@T�8h�Ws��)�sJD�n�����6����>���~���c��r~�2�ב�'�����Z�7#���T:�	�9!���� ��F�j�-+�Q���3g���!���oΦ��Eгo\������s����Z�|-���;Ta-7)z� _�f�~V����G�����g�A��{J��?���v1A����P ��ZA�i����M�9n=z��R*3�����~�Wﶙ�o��_�2����k����a��IKju��W�L&kyY�j$7y�^��.������D���%/��ڙ~k q@����±�;-��T���EˋyD��{��䑟b������.��Ę9i?����j�-�i؟B�X��L�l�K��^�r�S=����=smw {����"��9����g�[��
;~�W@1��$�������}N�^g}H�GǘN�n�"�9�j�<(���4���yM@9vbo�2�S��r/L�o`x����.�9�7����5�&┺w��^f6�lH$�J9��6��R�؂�byv:��B��,C�όV؝O�U���>��86ǿ�,��RM�!j2G=��d*��+O({��p�����c����H�=����Z�O�g�����rj���h��jB��������r�:�Q�g�"B���C/G묥��V��vAŬ5�c�I�Q*nߤ�;/�?���	��$e��\�q��.�&n~3�m�(���^]��?}���!��cZ�D��d���5ww���rho9~�i!�V�Q�������� ����W(��'��x�K������+�|x9�3�Rޡoʉ��ࡪ��P����>�ʊk��x�A�ܺ�������DS�~ϥ�����u⤏iО�IZ�6��j�mw�x�`��b�FS�B��\�-K���<�$H'�!w�I���д5�N��U���RFu��24�;g\� ��wNSҞ�����rQ��p�s\�a!	(��R/��($FK�v�h<rC�Ce�#!jj�?W���e�S�G	v��i���Z�hM/���t�}����5�����%�@�b�5C��`�w�U7�޹&�f/��xm�W�Y���a[r7	#@!.�L���o��ψ�W�f��*x����}��UcGc�@eZ-�î\Ry��b_�P�F��W���y��-}	B�m������b�Ӆ�L\�	�C�펔�v7R������@��v�Lᙧ�/��"��18C����Z2���Zߤə�+,yCة�yyC�����;����#����gY�S�AB}J�ykn�Q&Xe��g�H(ࣕ��ղu;���ZGY��*!�<��y�q�a���E�@�{?]���FgZZ�(0�;Nd~��	�h�C�p:_q>�T�^�:�fJ��\	�Q�*{9�J+.�F�f�krK� aW�T�+]ƞ����ݜ�%s��QO�'�6�L�Yl��F:��Te�ɸ@�;�1�G֡��f�����Tk����u��K�R���h�ځ��I��5��쓲s1a%#8�f����w��0%ĘW��#�7:G^bQS��
6z���@bu5Z��>�g}��A�ιD��&B��J���r��~��U8`/R�@X!�A���m��
0���pB~�~�z9G%���i��c!~D"sō�����ܟ��|�t��綘TO�����Zp�[�r��аZO!�P�\��Wɽ1���)�]}���ի���Uu)�Ї��1=�M;��A�sX9����h-7*k�����3:�ߙ) GK�d�![@�.�Q��h3i��[���j���0Yt�28S��Bf�]��;l��q��߈j�7_��A� O9�y�"�bФ�p�J.1�L�,8�%ʤ4�:��y_)E&i�@ͫb���)���Vٛ]4���K��=�xS+�d�m��&���326�'hK�6�?U�����9d�H��}��ʛ5���XI��?�&J�ͧ�7ā1<���6���)���R)�Osy6vU��hD�?�T���^�>���m?OJ�=�nM�ÿ�\Դ9���ٱ�m��`:�`�,���,9#S���>�̡���4�xt裯b�`��Q����>i˘�5p�f��q�~��Qp��ghі�:n+]P�S0�c���}��][\�# v@�Gj�/0h\�Zv]�����?i
_�f��w\���,���̤��ON�+`�jB�����ឱ��#�*9<XsJIg�#������I���&(�$��0�x�����\��7���ʂ�j~����U7�aO��Y�S�DX�3��ꝃ|�U�da ��Ɠ�.V�G�8�eޮ�lL=Q�S.o�4�@��_&2�R�t�խ�� ���f]��t��J�1O������l���+SȎ�e��[f�Ha��Ů��J��TVR�Ӗ���S�>�/�6���/�� 7��AU�9�̳�}r�1w�������*�Нk���Є^y�2&Xi���-׷�E7���x��y�7�͕K�}�5Y0��TbɷUtlm���a�㡞
0C��'�A�ܟ�O�t��+�i�p���?`B�����Ps����x�~$� 3��Z���XO�OG���!�3u7,��7q�Qqx�O� ��Z�=U4��C�7��,�T����CG�Z�q	�W���	�tq�!2M||b!#bTpL���t��.E����Ɵ��m�줣_ ��u�ڱ@�|�V����F>s���ճ8�P�����r����`D$~��^���p*�����GG�mX+�W2��Y�\�Lp�k&��]	0��H�^��W�^t����9d�Ő�w�1�b~N�1kO;�"��N����E}�~�L�������[�d].��fQ0@��e0*,�[�I@�LV��%�QT/���mw�H�ŐY��xFv+X�0C��b3M�:��.ĤY�e,�w-��Q �x�7�%q
�A~��a�[��fZ�t�߰��$�q�5�'�;���?�W�i��j�ćI9_�9}���tÕ62�8��G�L̺����5錭�8�0��?��Te653<4N��Z����*{�>^���^s��'����J�c��'d���C���%E���,V�A~b
k�����ƻ���+�����K=�D�`�u�?qr&���X��Xr��,�rz�0�d4�a���}?V�hZ��.�S�Ϝt����M����pe��ʀ���Ǔ����Y��o��w����}R2�x�W�8b*3�|�i4��٫0T˧���Ɉ����w�Vt��
���BTP�1��m	�)b��w=��{k6��-�]>WA�����N^Ť2��j�	�m�g���)=
,�)���أ.����]5�����͏h|�Ad�T��Զ����Y-1�"O����wn{0
\�[x�d�G�"��Mm���gi�����t vu���hy ���؆�<�Y/ƴ�s�7p�m宂YU�;d�'	[�`��P�zE2O��9��Ac�+�ʈ-c�e��%AlZrOof�r@:W�+�vzV���
7-��}9��Ԗ����s�n��d !mW�p��FxeBf���s��/.�}��ATq�m�g*(���H����O`����g�Vr����w�.U��VՏV�����z�P:�/[y�~*��p����d�g��} �A��E2e�<���&W�����5Wl+�.]>İ�Y���Y��W��gi:���r}3H"�N����o��K`U��Sᵊՠ&Xۃ@O�YGU���Q�@�q�w��|�Y�J���ɺ~*'Tq�2���oo�pE��x��g��z�U���R��� �pg�!n��e�ق���Ԭ���m7���a2V�h�E�.��<�iEp���mpG�@��F2]����8f�|_�c���f��h��p�ςf���W���Rd�%��L�h�����K���اT���.S15��;eSvƽ-o���s��W�~q+�!�~x��ù�Ѯ�P6��.~��!�po���i������d����aP�Ai?e��ԲN`��-�DOr��=�ˬ���1G>~TR@��fK���|�(���.t���;���ĤP�I�J���O�	$VF�w��D��e`�䋤@���oid�p�@9nV*�\oV��xL�ǡ��{X��ES:�}�Pa�˶7y�g����@:�*$���e��%����Y<a*����=�4�m7x����L�d52V}�D�� ��0ƪ���ohw��BjҟT����I?��8��miӉx�!Q�	Nn4��#ްU�c��A[��\>"�o��&$�rޗ��2.\�	j�D�ўA-�c���
5�Sœ�KΞ�V7Xi�
���n�f���=��M�q����8au�/���A{wa1�M䀹S��L6���Kl��r+O`�~��ڰ���������s��&���T�{B��NѡZj�
Py��K�
b@�X*�G�[�L��sViB'�d1|##4I������x�;YD�V��q���oH�{-Hw/ ;
�|�go�"������� ϫ6��,��:�x�Ba�@
�*v����4���aRePW5͒�T�5#C�\u�;1��a�"*L�Y?����4��	�X	n�.HW;F�3�B��QiOCmP�t#X#�~p��|)�J�߬i��=)��x&�O��yr��vT@��QR�)��2�+yk]�ݍ�_t\i���z��_� )]����2|д�Y'����ժ���*E
�^)/�xn���]sw*T�@���\�W�|��_������  �H��]��.t���M��] ��ݏVq�0H~2;hk�''�J׹��P�휓�yc)��T0�+(��(Ӫ��D	zdϬu�!��C�];�>5�Ϯ5M.B�nx����(�[Y��6+�3O�w3��wa��k,؜�c��bub�޺��O�\�Q��E��\�WV�k�Vl͡�� ��O�NF�����E�����~Ǘ����?�R\�dktc������Y�����]a/S�*�^tC]����P����IO�Q��+"��Ɏ��4�;Ds�3�Oߤ�;��k:=6�!V/$b�	&��b��ʊ�Z�����C}������D��-�.�?Kt��t�mM��aKO�� ��j�FPs�eM�y������Xr&�&@��W�\`Ɠ��i
>�Ds4���8���ap� մ�k)WA�<�T���S`;0L���n0l^M�V���#�l��5+�qL������zs;TtG:�`�ŋ�0�p��AoJ�g���&�[���Fo�3��>xJSC�{՛�l�Ьm�n�gưL�,�B�&ͯm���@�t�Lz�HS/���tE���>պ�WJ����e��3�?�[Nׯ��4�	ϐw/ߎrg1;�v�l���B������H��:�Q���1灔o7Z� �|\��2�S��@��V���A�| H��e�dN�� ���Hzx"Y�������������>/��b1{�xG\���f�4�\
�W�Q��t��� h��?�� R����7{�|Oy�^�\����D�N��hZª�su���%&!��	g,���R������_t.'��j�3��梂�Y6%��� t��cN��N��9��AF�@P\-���w~[�w�!���:ڔi�N��Z�)V&���|��➷��h����x��)#�dv�l�ڣ��CE��]C�`���	�rY;��}:�(�����7Λ���L�m 0�ʂ@h�jӱ1�Y��s�]�K1LL��f@�(#_��`q�	
Z����bbVf�i� �%	)ϲ7��ɪ`�,��"�6�;5r�����#���$Eco��N��aB�W�A�hQ`� QN�����@�
����^��.bf櫷��}�P�_/�6�/>�g"P4USX�c�����2H�є;�\��~Y��:�H���&��ZG��$6�K%)'1��4on[s����Q�x�D��b���ɀ���F�6�^ܳ~9۴o���a�3O��mw���2O%H��P��8x�YF����̐2�^���wI��J�5A���',Zn\��yq�#*6�P�1���E)p:'Qr���r$�}6gk��8v�DÿL�9��L���O�*�����~�c?��h�~�,�#y���-^��'��yu��ȭ|7��y>vO��pM�̠�a��[�A��_����$��R~OhfP�@K�z�_�W�ƀVN�$�[w�%I}I ���,����� ��G���h�V���B�Η|�AH����%���c3�M��Du���)f���O���=��g��B�����Ō&��ңk?�L�ˑw�N��5��"��ڏ@�(݉�b`?�������Ijj�S���s��TJ�
�e��o�l\~�=�誘���{��p��8$Cxu��:��OK2>1̣�_1���N��5��F�.�dGaK�m�?u�wPxb��[��$q�������P�!�ϵbkϙ����ٻSH	=�`
��$Ӈ��M^���_'ei�i8?�-��^���	���J�'P�Y��j#MoZ��?��&�}�����l���B��\<i�i�ֵF��#�%�ߙ�¸��~`a���/j�~�ʪ�F5���x��l�W�F�����@%0��^�J��sW¸F���^��^As�(���Q�c`Byu�OKYT�S�~�Y�:f�/,#�?��Y�
s�j�_'.���mf��k3��'�\Z�
,���������;��x,z����ݼd���h��>ENJ��H���f��-��@C���@�,�Ϲ��`�ȴ0,���g��4a�3g��M)�|4}��6�֊�G#h4\��!H��?�t��D$G�nx�D�7��u|����&�KӒD�X�xb�����g�?�t����O�L�e�u�5�hq�/�>�>�Un�����S��n[<^��)0k��<��t�p�	[�R�:]�1x�"�����TK4E��qY�iP0A%"��vu�'�sl���>�[u�QF�y�ce��ŉ�-�:�&҉Nc�6MQ˓F��sn|�u��{�0���-?��v�S��P'dI�v�lj�Ӧ?��Av7�<�ȧ�xT�*��m��Dfx�~���]��gC����i�ë66>Sjb�v���&H�J�!�#^�\ �X��m��s �y/Bp��4�t�c6�m���E��*�W=�em�ꃶ�Y�QN �߲����Tq��Ǜ�i�O�Bg|D=�J���tŭ���9�HM�t�66�8���D���S��`'���M32*{�wcݫ�w�;�;I���6ge��:N2-����?)� `��L(XƸ��{���s�{�QJ�"�lM3���(�jfK)���3|����\�j���z1��Wl�x���3�<RgM���s�(����ZRG�aT��5��kD�8��A�U�3�#�Ie��g�A��W����_瘪���ȱ��J�B�i�w�T7Y g�Σ����/N��t�Ry:�3�*P�v���S�#��c��898B�O7�ӀR��@ʣ�	nE�ML������G%KxZB�����T!�S����`��*��N�t��r�9�o�]j]	�l�D"�n��� ��$]@Nq$����z�t��+�״o=LF����I�L+�^O��O?���+�!A��-��T!Q�,���ڜI�s�i6���7�	�\K�Ws��Ÿ�Z�-`#y1��n�a~1a>+W�oS��R_Ȱ5B�T���%�v_���N�s�=�d�����\r.ɮ��Ǵ����JQ'J������i������OK/�U�<�B-�@�%������!�E�	@�p1O�ʎ�P�6�~�8�`պ�$�7!L��������9�����U���P�
�>����
�Rxp\�oMz�����8�+oe��J��c) �(�e#��L�Wݴ>Bn"4��!Y��:�$Ɓ�K#M�AW(�#���y���%$[^�̝�T����p$��3���Hl�m�"�I��_߱�E��ő��Y8����u=�cV������;��ۈ�ЄٌE����0������w�譟�!���d�A]�7�[ވ·{����qP�����:D�[�+��,�'��J2�c~/������j��S�S�����f���l=� ���ٴ��_�1%rj�ݑ�����.f�#3HI��Gr�'�m��}P"�35��gw)�u(dG�*
���]f<�X��^��>�p�د�Bw6��Q!g;�OI�d2�s�r��.Y9V�U����ge\�ϵ�����g� ���Rx.%[Z��s3��L�O����/�m� ��zD�?Z
ȉ����I�퉏.O�)_���P,�����`U�1a������ct@���sJsQ|�V#Xɾy�W�nC��� (�Q
��gT��--�:'!A})6���l6P���h�z�K�A�;A�U]�H)?��lbV�ۻ�nn���]um�|T���@Ĭf�i�cҾ$���6�N��[�It�b�彙J$H���r��vQ�sȐ�v���7�1�R��$�L�w���j�$Y1{iлz���_?th�'�\��"��m|�DZ����]D4��>Ϡ@}��y}7LX4���֥���&4�~2�������3�6�-7���N6^��Mˁ�7x�26n\�M�j�7h5db@�c�_��w`����I5}T�J�c��~��aP�fT!����K�x4�m%k1T@���/��	�8�]��zc&����˴�U+-j=.j�:��!O�g�
�݊��7������FVo���-�;�a��j[s�]��/��M�l-��M>�`��w�n}*0j��� �����w5��A�L2�>� ���avH�|9��e��_!��B,"Cb!�˘�X��~������P/��`�r��O�6O�`�u���\׀�Rq1	�)�oU��n����:��Y0��:?5��/U�!��eTT��&ꕳE�p�L(F��/��ja.���iz'�"����:�4�\�=[��-���r��L��<3@��R�Y�t���',�d�f��z��AH��79RDh7�l$��Z|N�e)a�8sg��u\l"���B��TY�tZKup!`�V$��&���4����i°>TB=s��r�8���S���/��F�Bf}U=����cy_��2W�O�,F�A�䑶��J+�X�x�`���|>�֪�>�hKU�0��.� XG��M���&ҳ2�yg�����0�QW�{�f�Y;D���V]j�Aq�8��٪y��__!�N�~��� ��UǹqJ�s3FW}�8R!�e)-��^��U�,�j'Kj�������87L��� �ـ,��1�P�)T��� �-�D^Y@mȡ��]���a$��s�2D�������ITgf9|=#��1��&�@����=<`��{������4:�%3���PXbYI��F,�'��Y��B����[��k���pSIo��	+�����ib��@8�o�Z�	�!��_��U�p�L�c�5�'�?z��Y�v=i��+�ݗ��&Κ���8��ԙ�h�V�����~5f1q�|cSp�&Z._X$2���r;��A�3I׿��h;V��௟��&��f���I��	�S���[:��:���^>���j���v�=T��߀����3z��#E�t���G�����}����r� �V�T&n������?~�
.k�L;<��L�?�rU�(�
d���,T��`��a~���a��b��:�XE�&��<\Í���[.[N3aKQ�F�6�YN�mX!�?Bu�xU�����t�wٮ��`�AF�8�|f,�!�s���7�v�7H�'\�G6�α�w%� ���$;����r6.t�Գ�PF�v.T�%a_G<O+�:@�.;�$==��0A;
�ì�KY#m�D�a���1n`u��p����U(b��8�1���f ݉�:��?�FY1QF�6h������-��X�0t���V7Ri�ߩ?��>^6 >D�└~l$5�A�~�D��Њ�u��x`A�C^ǽ�<wu���]wQ�$�쌙�Y]�'�*�֒Sδ�=�x��i�� %zkre�X�4Kg�2��EX@$Άx<�Ը{�N�x0K�Q1�G��<���(o�F}<W���7�J�����°�l!f^���I��N�*�f�%�-�:��-Te����x�bc>Y7�w3G�y�g�x����ݦdAJ�V̱�����Ð��	AD<.vETH���8o�g�7���]��>Df���=L����o�-��� �� ŭ��zwElY���M���-h�$/W�m�*}ud�*yv��[b�����3ȟ+_�09&�� #�Yg�ɀW��>nѮT���eݝ\ng0���ɋ�Y��4%���̎�(U{���,�,�g��ځ�E艰��!x���3�NroZN����,S��ǖ�ԕ�H;"�Qdj�WC�;I�^\��i�O�4]e����P䱴Hf��ڻ���$4�`�Z�� ���U��j\�D:P�"��KJ�0����G���/��e[�m��'�[���@.��{�e�u�x�?�E�Q����h4���/�cb�,�Ѧ�~�˵���gd��FJG�2�=5�ֆ�-�
�;kՀ1΢��==�A'�9�UT���nF�w�ǻ;�eƕb�*�j�&y9s�b�l8\�K�� �
�}�(h,�O��3>-H{�ɹ��x����t"q�Ü[��q-��a�'6�����zX���(�ƗY>O��t7hl P��ڼ)5�M���U�X�1i[O}S����2t�!/I��������M�`�.��o��^3��lR�aG��lL���R�PtoXY�!��ڕwJXe�r{�����8| V+.�>G�BG�4�Q�nV��J��aP��W�H%K�^���ٝ7�{�m�d��o�a��޾��O�R<.,�Lcvͬ�r�t���ږ�'�f��v,�#6s�3�`��	��Z
O�&��qY��	���+��@�>�{��Cj����$K+c�@�	�Z�`!Ţ^���R��N�
��p�&�C�ל��zn��)Z�n31�;O$'G�9�7���aT���U��i5T0�׏æ	�Y鹳[�-����O����m���߸,�m�mb��Zx̅�0 �.��E�5��j�I�}�tL�)qf?#�zF|��>����2�b�m�*�.������� ��:�?��KN�_��~ƣ��я�
W����^T6����iv���u�|բ^8���iQ��9Y���*�vvEܢ�L$�{��+e/j��]t(H9��u:?-�P��?UƜ+�|�Ƀ�C�b�]U\\��&2ҋ�f�H��6��Ճ��4�Q����.��U�)K̂&��Qo��r��磾����`#�r/g�	�0B�i~���\�j�-ө#�ԱF���j�N_���>;���u���7x�����E�鸥k27�DѴa�A=��ֵ�NЋ�q�Q��`a=�J����b�N��}��&����w�W[�"'����	N�V("׉��`;��v��nڡ�*�Њ���ig{�zC���u�Ӫ��L�^k��4C����3�RrA�ע�vv�5������~�GM���%�r*�3��a
\��w���_����_��R$(s��M������d+� 5��"ΰ��>�!����_����naL�H���r�mM$��B0��.�Q�Te��ei�!f�Y.���F�ɑ�v�/2 ��by[��2�k}����AsۏL}�\�:
�H����;�.���3��ުU��Mu��L�/�aO�H�^��S�5����V�{��C��m�m�hȇB���&��q�ʗ��F�f���yZ8�K�y}��SU���߰J�J�U�ϣA�?��L{̶B4�.Q��3n���9K.���j�P�*}\�v��#:ȏ.��&���8�ep��g|� ���m'�����l���n�ۥG/
���%�jO���&����%p�v����i0���Q|�X�4� �`���#h�:ƹ��Ɗ�� W�D���vB o�P�g7ߴ�&ll���$t'�0�wѤq8��4<]-���˧����b��s�5���in.=���0HX1ݛrT��I����şt{�STf⿳�V^�JÂ�J5�X�Ξ}�k��
O+ �[$\�Q̈́�;"cQUk�/E��c�� qz	M�n� �����O"�I���X��'l``QD���x��s�7��6|�X��>�+b3j�Dt�'��iur�(�t���V.���jPpN.e�<	:��9.k_���&b)�,Ý����ޏ�@Nm�R6��i#�O���)�Ѱ��3#���j����N�U)-��J�����h|;K��Dmd�x��N&;k�	X'�������,�6뷙#�� V�P�B�(��DP�Y:���;������F�	୼����N�#`,=�%�p"xy�0_��x�kp|۵�7�_g�JH��]#,-����Û�B�S�-�T��i��pUImr�&.�N��*��8�~��nfO�7��޾-��kɯ�q��_������l�p<z���E�M�,%�_9�t�-��h��i�
��~��[�f���a��[�A��d�@z�+(���[�أ
�����}.:+�4��ǐJ��}���S�`�dgfΜ�Gg�w5�޽�@�{�zF�Ϲe�;�C�@{i�p�π��e�e�,�����>2k��XS�=�8�Ý��q=֜712rӦA�{��\)�@׮kJmx(�B00O�Q��iT��Ď��[���/�r,���/���r�S>�C�g[�M�CC�by_��[��$X�6oO��4��)�[�X�s�;�3�^��s����F$5)+�����JG/���,�#�#-ׁ���+��~�T��b�H�o:}�8�X��CB>桋��O~DZ���E�U��9�Ӂ�^t�oʓ�bHSJ�<�HmL����>��<ӑ :�_�%��w��I`6?��.O�����+˒��uwi��V�c*����q���D��
��D�O�-���J">�Ҽ(�	c�	�2�~��8zM�}��6�h��N��->�#��=YV�[ε���8��]v���O{7<�&r۳���p��G9���nD v�4��m�O��G��@�4ܦ|�DJ�ġ��:"���;g/m��KFM)�d��!NGk�w���Vȓ���`?g�	>��m�=ի}�;0@����*�}�p���9��3U��jI4�mX�#Ī�C�zK�$�)��,?�žT.(�<�"��ζ�){R�mC3:/�����@8d?���vC��6L�Q�jŒ�5�W�A|�����Z:�V�w�QIk���H�=�����5���D�E��KB�l �������J\�z����t+K�8��BD��L� ���j�H�]�zp�u�t���/�*���P�9p�5P)���'�=����I���I}<4<�����]^�J���:�;�.��;Z�N���>wr�ۜ�a`��3���9�'$d�r�#g#
Î�4p��[Լbo�]L��1�!Q[�s0S}������}}O�����nņ���s�6�\<Z*�5�� E���W]#�L*=���]�}$���U@@��"e�gk*�t�-��l�O�a�QXb�~�m�h���|T�(��ۅ�L�E}�,��+�C����臭��
��N����Q�͕[d��`?
����J��e��6�U��w��'����;�Db��3))&�s�j2)tyI}(i�p`&�͔n��^���E���~!�����Y��<-.����2���O���
/���!��GvL�f�(x-B.<�+��k 
1P?����sbą����uE֒{I�`���^������A�[�spJ���^��0��d��J�ii]�,�����j����SҲ7�ڠ�{�9�gB<םb����[<r� `�	�?�F��ѱ�d4���@U�Z��aqܮfd��!k}�)��"2ߖy��j
���̿�5�h �/NR��E�2�{�{P��5����IQ֨�X���8����҅W���d+�BO�QI�]ECV�������،�|{��E2�HaNx�Y�:�'X�h���"�',٨L����`{|���T�k�'�`9E1Img4���C�hF� HX8P�(\��IÑ�f
����O�$��f C����N+w�j�V&z_�>�m	��;bJ�X#�&��('=v������)�/�`}ʹB���6HZ�U��v�� ��_1�k����ƅ`Z�l��%�o�^�K�m;[�WV�u�[��j3�紫
��q�\Ah1��-X���6��H ����x�MFa��MX/�bH�k�F�����x�)fb��t�;�U*��X�f��,jW :�ө(݆@��o�
@>&	�J����,��4��;��OiR���9b5�
����I;�SI��@�Ͽ& p�}���%��W�Z�[U���LY}<E{U���:Rڶ뒒F�#���%���,�]4��E�l���ZƊ��nY��p�����_�V�ٻ���%��v��x޼�"K����]��^��J�#���?P��	�O��~�o5Õ)�7 ��	�wܚs/���?P�g���l�.G�t���q�Q�p[�s^]�����C��#k�W+�3����6!����6EP
��;����QpȖ�F�a�����F�@\�æ�,��'m9�	V9�+�𹋦����?v�v�Ӕ�d[�0��� %�mə=K���M�q,U;(�����猃 ta{�u4KeV1܊_&zC!��V��m(���es�vX�S�Bg�>���.�r]�|���8?��p���'�s��})���!�(���!F���{x�^���{]��p�iT��!�,np�|EY�V�Y�M���6�� @�F�^�7����Y�D���A��l��K�#3y���$�]������ާ��7U�����mp,3O��1�<��ՁO��O`���ܗ�������P�SO�o�N�+fqn�ęQT�s���Wg>#����
>�j�f�/`%�t���>�e����F�(���$r���S��	�׋�k��
d��j��j*��(��x���\Εn�?�O^��̠:G�A�P~woYfЩ�F��Su"���-�Svd��ԍ`�d�eN1E(ȃ�^[�刋Į+1ۊ5s���x�p<�jb��j�x*v�,kٿ��-�#pA����0k����kF~���rj7��!��i�'	6U��-o_������f��	��D�N��vNvx��=g�m��]��bv�����K�8�cŘ��k��+����Im@���ř��q���v��v�O�f�2�܍���ьf�Qz|���)���ڸs��oX�չ���49��8}�e�e��.�.��1�O�'1��`�U}TU1C
b�"�~�h~�to]R�/lַ�%��E��Δ�AG%g�f\�.�L�w��p�D�5��*T+�*�vn�������_��tldnB`������;͍�����LiU�ǜ�h��G��mt^�	T@u�(�i>F�O.��{mrRg��@��1����U6�4D���v�P0ϊY������]�}ZQ������~ek0.Xӟ�yl����W=$�k�{��[)��D�ڧ��MM�m��w�kP'P,@������"�����Q����&�����4���ޔn�	��+���x�ח6��f �(T�f�|M���*��G3�>��8�����G�3�G�C��A��h�ф�SMT��*�����:=��e!�ʩ<k��2nǢ����}b�~�����;������ADCn���"0M�����t�ʩ=���	,�$��3����67<�H[�V+yEAnX'�>��1�D�b^6O���խ��.�s�ɟ�������=}�2��*;(��5���P�+�5�o�� =ʭW��o���$~��2<A_qX>,���F���,%K�FA���PkӉ�����8*@[0�q]��'�d��jՎ�~�����eF�0��Rdq�)��f�@�Qmm�N8^n+E ׊W<�K0��>��'��^:
R���4����ʘNOc����5�<�H��h�F츟CA"T�~�h�h�\��(64Y�F��@c*F�k����� ���'`tS~�c��@���/��!x������Т�W��������}aJn�W8��:�O�R�:P�CaM�5�9!�#��w�61-�"�M�#�>��Wg2;��:t��^�=���0r=��bsb�n��h7|�S��yq�͎&w�`q?��2�#b��!)\�=���� ��@�`���;�:��&���.+����
�iR�ͦN���=�O�i7%u�b�}nwRH��͋�d�f\����?ĥ7������u���&Er�Yʠ�)t쉛���e�
���� &t��N���T����wG� �@�6�3�:hg��Q7\V��Sܼ���N;J�W��G��q�
�Z���)�)���%�zk$�GR�{)��m�1��ﺚ�%ʱf��ǣ(?yg�16�}!ę~W_�,9���
��$����ҜT��vPq�������
6p���l�������AaQ2���{f�RF�!��)v���F�����P��6���E�;u�"c�7D���,}���6��M�S'!�Q����J���"}���}d�w�㪳�ͬ;�R�������3̯�x�`����"����J�n���G#E����D=�	��M�e��rp��Ybo����h�~�̣�5��	n��j���}F<����cH�K�{b�=����$w>��F��<"��>�tB�k��	G�&����!���|%�|W�<Y�Ԗ�Ј� t�rw<�lr�}>��z�R�L�洗�!����J���?~� �鏻.0��=���O�����ߨ^R�O�l��+�ߏ�#aX\57��K�$���(&����@�TJ1K���| 濵N&�\a��d'SH��q�g��b���5��1�H�Ϫ��'B*_6�>�؈T|����-;�� y\��xh�Ʈ���2Y��@�`ϠD���]��D�L\v�iC�'��o�ō�����-n���5����QV�m	�g��{K�{[����U��^���DI��x]r�Lq(<�㾙ņ�&�w9EI-�����7��Y�Ʌ��%<@Z_kSA�N�b�ޑ}ح��K-?'�z���D�[,"@y�u�B�H�zr0T0������˷�,"=�з�ʠ�K����y���|��v�) �����݄z��Z��_pG�n���a�o�M�z�0�V��;���hxt^�{:L��		`�&�X���_*�1ݖ�8��ke��`��?�p�X�����[���@Gϴ��,��MC���链T)u�P�垨� A)Xα�(,5p���
R٥�笳�-z$��k�}K�^�k͇5�B�V��l��a� �˕����˟�ͦ]3W=��d���|NH�N\���F�ԧ'��+5>���Ǫ�G�R�4	"I�D�&;�r>R-r���߫,$�{) �U�ң�/����h�<�9n�]�)eH������|Z���Ll���g=�D�����yFˣ��z�	�~�� `���諭o����)VRYSEP��eݸ�"4\1����`+M~����U G�1�%��R+jo�ab�)V�)ZiG�Jy�1Я��8hm�¢>��{�p�85����A'0H�����8Gnn��>�8��'>j��L"�wl{�Qu;��R�C��e���͡�$������#�Fc���AJ[<�W��M\������T���@���ֵ�Gs�у*$ ��6�N�ؗ�B��1	�'F5߱���8u��YIz���l�dtd�?����>9��mB���f�PO����m��?��y9\s��l�����Ou�a����p�D�rD���E<W>�T�r��f���6���h��M��;�s���6� ~CoO�>}��:r4�`�m��� ��F��V�<g9yd�+�e��XJ�T8�J<DΊ)O�[B�7�K=~�T&�hV'�P�Ov���p��ksh�@�l�mZTxI��״��PPR��<��G�c��G�&�	u��=\R��������(�%bz�υD:�/H��4�� ��0^�=���,�Ǣ��ex�X��+�b�T�{��R˪���p׊�10��98�	7�X�����y��b�����H���i�; ��J�ڎK�9�қ������� �zYW]��$'�^})��{�xJ������E���-!�xRز��ƓL� ��бx���i�N���|��^���;���K�[� O�#Ÿ��A��Wh��,��܍;��1S��TT�42� _n��.\v����Zڛ\[���gb����}Z�M��I���t�Sm9��ec�K�ad�o�&Z,�*�P�W���9�p�F_���W���f���V f�|pL�W=\j�_��`4~�
݄T%�c�4(9��hL��s�[H)�f��#z�.�6�3��(3V�Ww�p����~� WuP�v ѯ�rR� YIFdW��� 1&\O7��`��>~2e9��&ha��Ǆr����=�XSU��oNR�_����}!3�ߦ8���j͋t��&[L����3֕%F�L����&�a3wLFq��E�m�|EQ|Ēm���4�di+�Uun�^	#�[w�"*��f� �(�s��j4�d����[��u���5$�_!���s͕Z+�-ֆ�hd&��ȗk��^�	�`�J�N~ZW|PZ��l��7�l�
!��������_��v�b�Ǻ��w��ɜ�Q͘RRX��w�v��>M�SA�<T��?FW/�
I��͈0��L{��PE�L�bN	�,�`�a�b�Y�i����qV.���V￨�!hMnq�F����n>�;�p��i'�h�w�m���H��
�ďkrΆ�] ��m{�C!P�����v���J��*d	[Н�Q� $�c�}��;_��U�?g��u����ͳ��#�U�bUZ�A���xĎ�'��_l�̺i��sYc#+�����˞&@�Ƽo+ˁ�RQ��[��:`p�˞�΢k��@ȝX_�=���y�R�ˀ�z���deh�_��
[uwb�f%��n̓;��oɎu-TyG��4���)B����[�w��]�	�$��z��g�نBmr �YX� 8�7�7|q	�[W�)F�ǋ�l;lߣ����c9wvGՉ�`>���QG�Pt��q��Kw�Z��^w���yDD�u{8�-���ld��0��ն6�������Y���DZ� wB�9M���cW�k��|%����]�����ȉRX�ʿ>�f�2���;K� /�#��g��$Z
"����8B�k^��d�����\�R��;����i���`����8�pJ���w�=�P�޿��5�%+�Z�X�Ҁ����:�����0ؑ�P��CZ%	Y)�\���(�.Wz�u7��?M�-Lѳ�Y�Qd�qKSLк.KL� ���_�WZ�UrS_�=D7��/{Ś�r�JD�n�5"���X�i���3,��J�nÇ�u�eyR���P���i�W�Ͳ�)�ɼ���=Ir�1�U��{����-���ɁH"�-��s~v���"���c��*�D��V� �mtU�_���!��ul: YJ�x�zH|~����o�2(��cZ1q����9{�I�|�2��B��~S�0Y��Qb�m��X��KC(���hZ��aP���"��j���bhYa�8Ŗ�d���:H�j_����S/�kV�� ���og3`�O��h �MAu��>��E��-8��U��ף���d�G~��Hqy��9��t/���r�Ԯ��3� �@<�6#s��a�Y�tɦ'�5"q��CD�=�&�9'J��x�Łؖ���}泙
-��%�3��zz�]D�_�W2����O-3�H �}.�>�����ҳ���a'���V���;�a�'G�2�iB���#�_9�a�q�S���Ǭ�K��b���K5|S���o%i��k�\eg;"F�ܑ��
���O� ��&F��]���
(�sXXۘ��/ι+���������A	�����E�C����p�����˲�/*�e���"� �tYj���N3��w��^n�V}V��(��T���x�	���b���w��d��8xH�6��Igvz|�L�~�a�:�ĠiJ0ū
i-=���t#�Wre}jW5Y��I��=Þ<�f����Xk�C�\e�S�P���G��~Ba�� �����	L���]�����"�S"�2�,����O��z#�d?t����Yu-�n���Ƕ�l�X�����:<U����Q���� u(��R661��*�@����~k,8��΋:����1hkm�bmg}���A�>m����k3D�o���3��Bl@!��Q� �fe���60f��Y�Ǜ;�3n����t�"�� �{�����ɨ�:h:��C�����RYm��̪!��-�����+�(x[�co��!�^�Ӽ�gv��E]�i5��׸}��w�Q���<�8}/��ok��]#�~e`g����h�p� ����{s��m6f��3P��N �
���P*)����9-�����7��6�9*� �!�/>ۈ����ڝ!L��q3S�@��-��:CY��g��s�O~l?B�n��U;��k�β�&pER�M/>�o���M��rY�L?���b�8��r!$���j�D#כ!��a�9��*��"���yW���T��e����B�ȧԲ 7Ln�M��I`c�y��?�NI��x�-~x0�$��A���?֮�i����.�Ϝu3c���8m{���g����夙0���**��֢�D��9U��~�3"g���O��4�ݣ��O��|#��j,���\_�\�8Lo��1Ȱ�,�Bq�hh�Ī��q;-ЗQ?\���HCti�gl1Od���U��&�QwN��r��1�$�2D�#�3d��<2s���a0�XN9�"�uCG[��w>\}�#�!�(r��4'����*�3�iz"J�]�E���Km,v���s&dqR�ɀ$�|��䀗uۘ�Nb!�DQ��ϕ�+8�m�w���o��,K�l+Q�_�A5,��u�_���T>7�v٘I�J���d�E8f��kNl�p�`8�kb����RId�_E6���*0���3	^����˥�����a+گ
�Vy���y�jN)%�U���^�5�e���4�{�<^���f`�zb�ؽ�dg���i�ON��Y�� ݠ37���+����A�<��ßѯ��p��35�SZH0v�ܠ�o�'���miҺ��3=��J��������7��|I�h ������f���J�ySɍʾ��	p�vfo�8�3��]y��w_���a9!�:v�=k-�v���z��_@���`7U��7Ik#���!&�!ӂZcz���%T.2� o�`�k�����(BK� t����qv�0�1�H,.p��H�DbY�G�t�P��(%��y�dAf�E�2W��uʋ?�Qʽ}=5'��	��� G~���6:m���L�
h��H��r��t_�Ϗ����'�/'�4\��r�1�؅'�&�Ҟ@��,�/*��A8 ў�]�p����� �-Ul|�s��A�˵�ļQ`�����L�j�esD��.�4f��4�uX��yk���@[ݷ)`�������.q_i7)�p� �2r~Ŵ��j|GR��9V���ں��w��e��8�hGB�Hm-������ �)���%AX�wq�,tMG�cc�����֞p[�"���	O��|�Y�$H�5��k�zM�>4�"��☹�tx]x����F��k�p�D���d<�\$^�(��ZۚhR���&H������n?�>>����������X�K�{?�>�]n���a���g�&�_*s�j���*�D�ɢ����р�5�3��.P;!)��Mk]�a�iY��P���iwH��4�T��k��tL�)#r�*�hG�T8�p�>�,�b�X��3��HH]�mZS��wBY�;���hA+L���7��71��à�қ?�Jɳ9��U�5�C�K���ń�@<��2z�\�O�z�����:�c�#|�.uN�J�"T����R�&:�旋�J�A�J��BE=_c�s��B���'�}�	6ܯ��u��P�[�$�1��ݕ[#6�M<�̀a4���z��˅Ϡv��4��[����c�� ��<@8}?�?!Q���-ߩ]�qX�b������d� �
��=���G�Q�T�m�U���g5Dxg^�6�GjKo4�bI�W/���ݧp1���7��=���G^sM���)��2&�.y��y�z"��`P��9̝��jy�=���w�MU��N0������k�����W�r�KfpQ���.�\�Cx8��Q�j�J�3B��1)�#\
�R�U��SY�^l�H��F�n`JeU�*�2�������%V~�՝�r'1�I�fVI��$���[����1������~vur)� ��)��,S�9'�����i훓:B��U��+C$���4��̹߭��d@�g��E�Ojm�b���I�{j	��m�5��$�X��'���ڻ��؂b����u��^����.�����"�O�r��qU-��I�#�����^(�ܡ��OQ�����Nl+b9�i��灄>�[߄��l=# ~�1**��g&���K1��#F:?D,��2��Y7)�'U��5B��v@���<=�X����*'���(�(�����w��#:m���f
s��:E��R��8�K�:���d�����t?�#8z��%Ǝ ��=؞6�͸����r�2��م\;'��|����X+=��0�@�����z��	Z�Hh]s9κ�,�����0V>��A���B>��񲽴�y�'�Ƅ�f�����)���8GM�N=q��6��-s~iϲ�jD�Q��!��/�N8�V��n�v��8�����UP[T1E�L1G��1]k�ѡC�����1�p2��x���Ѱ���g!�I�˟7���,���Xc'�[LCM�.��i,I&����x/
Ж^AĽ�l\
�t��.�!a�s&EROM�A�u�S��S�Ӗ�Q��b�Ĭ��}�9qMR>ݘ�(��x�F�&���1LÕ|g8�ɐA�Tz�c�E��_�	鹽��Fۭt���sE������s0���vm��J�r�O~1�H�n[�����w�4���9�˺��hcIiސ��lz%�����s��U�2���1 ��[�d�/q	J� �����;�b��j�B�H~7�4�P8D~f��,?��䏧���\HS��Ydhf/��>%gb�"��blg7� �'E�jY�mu���jz��%T	U����e�w��1�9�:��`ο;��h�r㪼�`%e��E�B93���8��O�х��6H	��oU
�e=[�0�57�w���	&�Y�o�x?�90b�"�V��!,�V���1x-Ag�xy�vi\E5��d����h�݆W��%�/D�;���>9ᳳ3x�@qX� �e�"CۅD�)��,Mw����C}�ԗ��h	#a��*A6,�N�q*'*T�@笮�ם���ڥ��i�e���b2��ᯢ;`�����2
�����L��k��X�D��l��j�[�H�E�r�H��i�Y�F6RD:3����w�Y����h�(q]op�d�ؕX�=Z_����ߟT�C��bpX�M�r�I%݅���jl��g�8��xa�xUb^��i�{a�^��_����rqdO���iԓ���J���``� \�� ��z��"��1�� ;�n�RݸaIԗ�M>W".uH�z<�
�+R<H�>���[��*��u�*�7�_��2�W���^��j6?�I�����%���9�9�dUBwbw�sϨ�e��gxX�9y� >Q֏AԜ�	㎽�1'�Nʢ����3,��^��} �t��h��_��B��te����¬����0L_����MA{ǖ�8'�D�tC�.�&�e�X�����NKŃ��� N-�j~�����S�<����#�����'��*GF��)�r~|����1��[� }�XZ��)�-@�O^�����!d��W�s5zW�O�R�4~nb��r�c[N,Y(�`v|�X�$^G�l��BA ��n�C����2Gb�;�¨��������R�T�-0 p���y�YIRgy:��� {v�tH͌�v	lw���1/e���{���V��{I4'-�v��q�wt.� y3�\������:g�F�ȧ�ٺ�zd]��p��#C��]$k�n��1��Z��q�k��_�v��pU��e:�&��W�FN�x:VHz+S�V���/w����h:O2�mD�%�8 ��~��M� O��C����E=umi�8A���VBQ�{�7��w��XT��	2��ǁd������HD�r	�����G|��vz����T�@Q5eމ록X�(�L�h[����x��Ù�G0�(�|�K���d�(��ՁS�J���٪��IH����-����V�(c-%~�N�o;z����*��=ٶ�H����
`����]X����FP�3���%��jn@�΂�f�����z�o�i�l���� �ھ�~1�&DR�[�K��:�L��z��9>�<xA3�Z2$c=���HgԊ� ?�[�T�ssY�eE�
^�$�:6�Qaf�/7(�2:���94(�^��c|	����N��ۑ����Y��!�� ��b��)9�Lb���8� P�~
�`��?Q3_uz�b�u�*�,������<�ԲB��NU]�شg1=�Z�mˀ��8y�W�pY�,'�A[�+'�,� m4;ǘ�!H��tp��7Ε�?�%�EW*�B7���d�5��_me��"�g(����a!ʛ�.Lp!]
�Xlͅ5�����J�S���@h�Q�D 	�H'ݟ����~s�[���
Ҹ�Ңh�h��D�E�"B���e{Z��~a�e��<�&عQ�D�5J���u,��y� �<���_��zW�.��4n*���m��F�
,��(���{�l�jM_��ǀɛ�LfA�/���K���]���"Q���{$�����$��R�1��/��L�j)C��~�=�o��dL|��ˠWn[G�8U��ha�����W��dp&��"�Qџ�,����XsبW�};�R,Ii]�,�gۋ �Y�H)�eu�!��������ǌ2�.]#�?�6m5ۛM�a������>Xat)N4.��u$*���Z�`����pb���Ԟ��0�h���a�Z1D�bv��*��*��U[��Y���/�=P�7�w�v��W���T�����Q�=tH)����ܑ,�J)R���N<�O2�ߝ������O9S��
	_�M���q�|P���B�!F�c(��c�/��5����o;FwR,h|�hC���S��ܳ:GRԶ#A��-�]"K(x�>И+o�B��PaPФŽZ� ��Cq�$~�Y����zY*3Sĳk�����e
�D�M^cy�:��P�l���Žy'�#���H�]6��̶Wyc"��d�d�;h#��F���{�~6�rG�@�90��E$yˣ��~�d��Z����, jW�������@�����f�A8 &4�ͫd����tj��6��f��ht#��Ĝ�p)�5QeW�Qcѳl�1c6���Σ�G���+��w�L��'��3���s%j��Ɠ67�k������{Ѫ:G��v��b{����[�n6�W�@K��7�4P�zA\�~9�m�	��!�Q�	F��;�v��䉗}�ؓ�Y�h6'��gf$I6��ߖk4�U��'.- V�O��s�!4��f����/����^�%d�_�r]iH�X�u�`�K�.�m�;����U�k����*Wz}��Ũs�~0u�5HPSm��5ף"���-�æB�R�&�T�v#�HUO$�����SEb��|���?���	*�'U�$�1��ꇱ.	G�c�:R�%��7J @���E�z�ڬ�Nw.>V��V�33�n_W,Ŵy�R��#P���
�~�o���$�j�|\��p�³>P�&�߂��c�2�5���~y��3�x%����Wի ��!��#�k೽�+.��k	�T��y�'���� �a��A��`�ho�r���������穢ݥ��b��3�N��	����\$5g�����!|�c�AX>9#τXzp֊}b���3^�,N�l��>����Ǟ�(5���f;s������A%�E��)|�����]�����%�rDTN���jol��&�Ӂ�۔k�-N�и�w[�Z�,7m���QuK�/B=UAW��)C�Zt6���X���6$�ni�>|i���¢�`�1Ba�N˥�,�"���`�}�KP���\���@��Co�=��5t�},y��[�p�1Oڔ�sM:��a^Z24-�G�\�g�K�(�+�H�C�62�?�$���HWӜ�%Z|�PQB_�����AT[.�"�;3a��q,LB��+��^�����BY ��\��6� Ĥv�i<�y�V�KZI��z�rcO���I�a*�ֵȚR���$�d\72��X��ZLФC�(�R���Du^����9hpHOQ[e��뿞�}Y�D,��L���XK���
�������ԅ'
����4�����å�(���B��F�ẕ_of�Q��/��f_��3�;���e�hӑ - C�|��_9��w琎�,�p�E�H!�̬��Hc��_�ҝ�K�6U���!Ln�obX�	��H��
W�������p�?۬穒����u\xl0���FI��j7��O����U���Pl���E����(�gpP��ң~#�W,R��D~$�<\�ݖ@/T�P�2���.��Sg�ː��o~��؂Y�F�;�[yխd�*����UV���[f��_���G��!������KC+�s,�L>U�|�}@�j�Q��Z��Ɨg��>ത��M���.�F:�:�> �ݻ��E�:�e����5�Y<Y�n�%Y�"V��t/�� ���`�;w��!�z2+spm�CP*S�¹��@T��F� T�J�<O���"�� ��{�N��HPS���� �|�3���icZ�U�[�1�ܣ�>w�P:칊������[��&����ڱ��Ф���I��,\R�/g�1�"�x�;yǪ��[������V���0� �oml�Wqi��Y��2�ni"Ϋt��󬡛s?���X���2Jڦ�ʂ,zw�DڅW���)=N����ŋ��c���{�p��Y�`�'6�5����K�>	*4���P�_��Z�#n��R89&(�\��)p�d]C�\��9����b��=��^�N��=�i��}B��ú���[�Ι$����l�}����'d�R�K�e�}n�
�x*���}z-J�p�f���]��/,9�:+L�*Ff\ǫ�e���D�2�,ּ��2�`&��x*��wL�������n�Ү��Yq
^��|{�Ӊ7���S�I5L����y�Dʐ�3,X^��fIx�oS�B\��t�7zt�V��&�������ow*!�Fh�QI�ʈ�t��@%_�	[�S{&��eI�s�<8F�v^�ܛ�ƀגTW��6-���4Zؒz0�W�%v		��|ہ3yJJ����bmP�55�}�7J�y���ҝ���gG�6A�~�@N�	I��!�`�8vN���g?^��D����!О��g�1��qjUp�5����
�@��p�؄W�Op]ŏ��ُ�X�vK�����a6�r�%{���ě�$��Ls������2�&�����*���W�NY�<��Ȭ��� o�Y�rζl���@���>��(���)�k�~�Ֆ0��t�*�R�%�N��>(��O��n��p���(�d��c��1���^�����$q6W/���Xl�������H+�Uㄔ�~����A��r��]�ayyK�TU���%�g�l���æ�{�C�˩��	`{���P�Sm:��a�t����� ��-xkF�)�8�m9 ��KX��-)�gT�Ve�+nId,Wd�^+�x��8����d����D|I=wP_�_�c�d5^r;Ԗ��w'YA����h�L:��w�sti/�6�DfL�	��a�?�R�'�V��a0��9N��ڽƆ:%ƀ��?�����p��]H���T������ǘ*�DT�j�q$U���� �\:ݕ��5�c�|v0j�>RoeR/C��B���P�`�l`�yʱ���d�!s�zw���Z
<+Dk�%ca0,ޣY]Ҕ��޾�~f�В���<OΘ��-�BR��I�e'��g �h��OEJ�ʾ�!�P�i��F�g,���.ww8��n�����f}HX(�'蜤G7����d<<���>!���.��=�|� �/��K;S�kXœ��>b+�X{�91�ρ!]��������{���\ҐF�L���.Jv%&�;Mq����wY�1)|C>��NGҵ�����7��lc0D(���K̆1�5*�#��%sB�����W����ېwf?��'��d#�<�������8ҧ����JG��)U��E@ad\WB�c&D�m��DX�Uʲ������t��}QG87Q=f�(�=?w���(����1Txb����U����сh�����Ѥ=�-����g�K�0?�z�ㄔUz�:rsғ�	E�M���u7��r_h�	���������,�{�=Sp�2s����jM`Ǯ�3̳�*{���\L�nT��Jl?�or�D�Q�e�Z���������Uu,���*F��oL��ݴ��:d�J�%�{G�G��>�f*�R5���8�ʉˇ_��o�Ⱦ?nL6T� �[ʠ�5��e>�]�"�z����3N���\�Q�sn�/�&�6ǽ�v����ۥ��3Ѝ+T����A�/�Z�~D$]�J���<���!��@j�5�{Q�a9Z�K\�e;�<�Ğ\c���2�,��Z�W|�0Q���������ߏ��,�O���_i���x�)��W��yj�Ӓ�Jlpf����o(�T���oe�X�����T�[J��V�o��.��qK�
�C�z�;g��S����_C���%8or�I���j5������$�`.��ݗ�n�����6�bY�|�J�k��(�Q)��r�?bqiZ�N�s���m;��`�c��E����xH85Lh']�a�Q6_�FS朑I5�������aYV.�����Ck.�w&ec�,�A<Gbxg$�5�_�����lhY��As�DI����t�.	�B��TBļ�#)`
fڈNG?�r2Pw�=+�,�s`�gaqy��!�6n���I���mO�9{z�e�{��'��Z=(,N��o�	�*(�{��k�I�o�\K��/m�w�C02Z�)B�j�+qzCiw��c7����2�f�u��øC�>[ʾ�\%��U�I��Xfw��pJ��b�e������ P>E2�W�P�׺f�g�KZa/V�\/��'a�E�7(�7���/�� B@�+��T����qbmj8 Q����-�Y@sg�T��"��A6��G�'�R.�x/��`Z�"�Ar�$`v�{p�,�����3	��R|_�p�`��dh�B�'� [�Z���y��t����T��t�
���Li��S"h:8�_�J�̄;�Y3J�&+�xBu��rG
5p
z�څ�-}�1.b�-�����hĜ_��07*���vM���RO"�9b>��~�ܳ�1^���a5�}ņ_%�b�t���%E?��Q�:��c=�9� �H v%rZj�Db�����7��ɸ�?v�c;'��Ū�=߉��N��f�M�q3[��O��<�AED�n*�K��F�P�?&��2��g��zV_���48^�I�5�AL9�9Y��"B�qS���,Y�m3L(����)��)�c���W
�l4A��� ��O����:��G?��߫ˋA~�{��X�x�a�䜆��6�~��� �Ք�v������݄<�l&�`������"�3����{�Q$N�b5lC���G<Q�`Yف=�h*?Y���#�O��׀�������~�;�~Gb�N�9^P7LB����t��9s�2Ft�^�{H��<��X�xs/#Z� �[:3�DN.Qp�\�?�]ŗ�_����=�ߔ�#�-J�N�`�#���cQ�f�E��j��]�[m�,0?��H��ƀ/��PVd�r�wn�m��D� w)����
���kRMu�ç6`��핊��W�����9F��������n��h��;TV���Ӝݧ�<��	֦��2/g���o~��؋��K7�8��]��y+$h���<ާD.�-3���UU�Ru�`]�����U�|����~�7|�nt�,���V�����ڷ��PVI{~�b8:�K�����I�rf��xB<��.(��N�^/�\㯲}��B.���o-,�����{j���R6c��P������y�4��z]�����
�oP)�|�c1���L�ֵK�O���",�i-�a�E�P �ȏ�����A��� ������+�W�p���2��d���o�A�f1E@�X[�>�ŅgxC&b���|
�!�?a�H��(�&e��(�
ϗ1�#���)��r��+�2����{�Uf!(2�_��nU�y9��)�%�%$cs�n���[L2�n��=yA�d|)A�!���n|ݗ{ۗ���D�7�zU���b0�?�����J���3�'J��k;�<�$<���w���6����� �hPDeP��Γ��:).��{�O؈[��C�Dm�H.�5}���@�	c'8���>���ĸ��'SO(��$�|��;7�~o��h�$Bd�Ny�3��e)�2�tJ�rcI\Uty�b� =^��.�d��Z�t�
{�A�V�|lv@�n*+���&� ��Փ�vV�����}���7�+�d�����߬ Q=Ct,��Ҿwݮ*O7��'c�>��B"���P̥w:z��d�T>�q�an	h�9�Q8�%��BӨ���侇��?B.�V��O����A���҅��p��_�C��RW#�ϐ�Z��eݸM�����[1c]�ty>�Au�^l����AE��p��[���\��{�:�/oN�Y}��:��甖�?['n��eA1�~��Rԍ���`��p�d�����༩8�@͘���$��ꪝ6��E[�^a�ǕB� !�h�>v����`����NI8�ؿ�4"%%�> ��Ă�a��C�`-��_�J"��k������_�'Z
7�Z~�(�0;�qƞ�<|�yX�~��ԲpOx��s'?���1^3n����`3Uj��Zv��DX��.�'�sQ�Fw��>�=�nl#umc�k3�qT�
�F\�y��Q��۟��s�b[��S!MV,�I�rJ�k�5����>@���!�P��~��+�˜S~�*�:e4��k�u�X��A�PuJ�s{�ۋ}��UA T遡�|p�12�Qnk4���+����N�Dv3��F4XF.���-�]0������@k�:)�D��X���Bl�xл�W��ӿ=��kE�:3�!��+��H��#=�N�x�4#7@d6X�΢�Q4�����?R���^8��pW�F/����IB	b�s�^Y��U���+�ю�m�T�4����D�[��w6�I&UD$��z��<l��U#�:��Kf�cǅz&Ja�V�F��p��z��Y҇��������N䂲�#ݵ�� F{h�hZ���]�=�D�C�_�FZ���Kϛ\�I�#���0s����z�!v�͖�����&(��P;E�I�D����3,8�{�[�f�b����$�t`��]��+ P��ig�cmP��+� ь�$(3�oo^���"1ۦY�#�خ��mF��/n���:y{B�����k�Qƒ9;�� �Cb��y���M�L�W��W}�Y���t8����]�B�J�)R������E��I� ʼ���C�/��YT��09,>�m��Y���w- �4�A{ȡ�����T��Ǟ�V���|į�7�q��[���f�ŷ:�&�U��q|�px<�H�������L�9)��6�1P�d���̪�wk��T`v��DwQ0�_�������0/w�|�/���_��k�v���n���N����*�1A�o��$}̞��S>B����7!��|._Y�'��N>�ES���	9�p	�%v�렅����!�L{�i�zB�<�)��W-id����.^�z�.�E�R!�K�e
�u�)��p�c���fC��aѭ�.{�>��S#ת��C��$��Es�*�l��S�<�|�[�c2i������.>�-j��^t�Pj��O��>�W�x=}hr�W����@V���ic�[(�kfS�Sʈ��~ٶ�l_�A�,���i$U�֯X��mFE�߄6xL���V�Aɖm�}� �����	�境��)
�@eɃ�IkN[g��+M
i/F�ܻ���{ӳ΂�hD��y�GYw1x��J�̂��'���X�Q䢛E�ߞ�M"�7|_]���d���sr뼈�iH�i0�|�E���(\�}�^
�ˠp��z�~�(d�v�ܝ��e�]�a�� ���������iI��U*�ƫ7�#2r0�%�O���:R���m����ns�@^/�~gӽ'��ck{�X��)���ż�=�tx��Vj�V�>�G�im0Dj�: �P,Y�+�[KU��,�p�����<(;����L�Ŕ�������2�����P�p�	L��~�J�M&������C�h���"�"�}����}4��Bfqpէϭ  ӃS�?꬗��J�يj���~��z.K۔t&:*�b]|�M&�t��R�I�k�QQ&�xWXeZ�{$�ZZ#DY�dS��7�G����9�
6H��!&t�g�EPK'[vt�n~�`8gr�@Z�L(��&���CFb����&���◛�#`��+��I�F����� ��� .lI�(a�izZ	g�����d:t�޻7>�'��v|SETm:����#���U�1��Jp5��y�����JT�S0T ��[ڲXlD�������&�lz��]�w��eo�<��J�y�c��@n ��2����J|N(a@*[��x@��Έ�2�5m��h0*,~Ӳ��[�gI�K�Dr���v~?z���So {�E�'�D���d�W�\Z�����*!�Z���������Է(��o.�{)nʂ* 1RG���4�գ�f��_�1(�G#ʰ�#��"3.��1���2�����������6)�����.@ ��,O��y���f{��_�ff�:k�h��hI(����Te- ]nr�������T�N��>��K)����Ot(�L��������>����]�ٓ�+�m�����mq�����6C��ڒw�@�A�uS<�kz�>��I����)H�?=�&Ȩ*IVN���V҈�9�e�ͅDғ+Z���^jk����L�	,�a ���~V�`W5/��	Sh��z�.�5ݯ����X)�vShuq���pUb���l��~���!��M�X�>(�$x�1�t�xƻׄ���S:��׫�}��zlgd�1�!��H{��^�����
���:��>���yXz[�>��7�&��>{�+�����X�NW�E�Y��GQ�s���{��u	�c���Ֆ�Vg�W"�K����W8��r~�D���M:hHxz�4�r ��v��no�qj�=�w�����?�ŲIy��M`{�/t�����'i���*[��
�z�-��B���~Ї�Z����)	}T[<! ���=V������O��MP��{��/�)��Q�';�����D�E9��IW�oy�h5���΄0�˘$��>�<[1��Q�s�㈸��V��z�!�C�����u���6	� om�r���j�u�IE;R8GQ
�.ǩ=~m���h�4D~P����]c5׏P���R�:�яi���z�I���J �Y0��j�U5�ŏ�5��RU�T��3ԣH4Xp�:޺^D���y�,��:RL�Ŏ�r�\0/�����
{���/J�T6�<!�œ�z�g)�D!z� L#���3׭�ʇX�Eȁٽ�����z�inE�H��o��z�u %�ũ��u���]6�8���0# :�K�B��&7�O�ᝐ�z��.�Of=��wh��	FF�	NU}��1�xj
�y#4t�Oz�vp��� TS><���l8x1x=�\�����E��~hK���r?���pd�:��B��D��?�6��]��ʴ@�U�z��uڦ�U� ���Dus+´�l��+Q�b}w��c��TΘ�5I
�FY�t7��F���@�@El�g�G�h@��BK����a�`am��t�/Ӧ��\q$�`���a��dE�Ӆ܈��T��ˇS��k-|G@ �?����'.�R�n�QwƢ�(���@O櫯�ͬ������ I�p�m�(��.%)2M���u�ZU%@��}ժ��S������|��<����Y
ϣ�|2σNm�m6��z`WL���?2�����iM���V�IS�igą������F���7O��\A�����@> ��Z=�Հ=��;/�lr���9h��܃2��'e�����ylK(ް�k�U� ������jG������s`=cؙ�t:>PR�$Ħ�Ǩ�����Լ	K�u����a����L����mK��L����:�n�j{6�&�{��7�#���Hb�<{2��L+z:�5���rMسx�g�]ڻq���X��lk	���O��"�N�P�ŉk�դ�M ,�A�q���[�JQC��@��@���Ȧ�ί5$s�k��t�i<u쵭NF�+(F�|#׍���j!�ha�#�3�~����(�xL2ti��L��m�I>[lXKΓ�,s��T��"�u�񐘢�n�JQPzր�b�R|	/�)���N�^��I"��;<}T�5\�$xF�}�"������ji��C�N]\�^����k_�zdR�ZW�����/��X��Le�����B\�l�79b��@j���
onlAk�0e\E�M!���51�wz@X���z��=��M�!�5�r�{��l�n�N!�!B��-NQ�XH�?a�:�}F����8W]��h��2���#�
w���z�JEt�~=lˮ�m!e��ܑ��ɣU5�ن�E+�9��q��hC��fËHFW��BUE�"��iA�P��.w� @2���� Y�tP�*s׃��F}{ �G�,���^m�J'u�J�|����u�F�H�]�B�';����7� ��ǭ�5c�r�����S��C� ��������5���<�;Ve��G7��)8)������
3��B��4���+6��;7����nw�⭞st�9<���X�N�}��S���-x	�z���j�N{���`3�Z_u�����S����|���hl H���i^��m*ψ��g}�驞cM3Qv�w0E@�TY1��P�O��M\�W�	�'A�"F��׈̡D���,�n�B��� :#�
�s}� ��'�	��Y��J�9�-밥ĥ0�5>� �w���[��X	a��t�wmT��d$w\�[A������I�%Q�9�ί�d�4��;.��)������4��/��[T��Pd^~MyO�\��|�WN�!D����+�߃���M*���A �Әn�!n�����Ӡ2�"Lm~_�r'��*��Pm�M� �G �|M���٥2R�S`%%e����萊�+�P��,��Nín�><��|��͚Ī �q[]��Aoб�xx>Hg1�tȗP�p7<������u�u�Slr�#?���L���$؝Db�����G�D�Ƥ���6ưO��Oi�5h�7��"����(�i	b:��(W�J��s5R�֗B/�?��@Y���,�cG�l�b����N�pt�K�M���L�XFX&��9����h
a��/�ܩ����$*�S�$@�D������h�����!%l��I�/F#�dS�fyY�/�E�J�t� ��rè�b6���F� ��.=��	�h�.I�M�`R�L�:s���V�.�cc��ARѦZ����&��S��F^�Y3D?iO�~�;��F�M�i��?���d!UU�!�}�a�y�<�c|�>$"��40fS�g�����HRС�m�!�	���n�%��Ǔ�^�!���`U����6�x��J�"&�:��¼@!����U�U�m�����1��0������-�KU��aT���:��u�U���|4�x#�/���(7R����j&����w�R���l��l#��J9���� kC���o��0�c,p~�w!���l/m󝗄6�6]��DR��Aǩ���N*_���Q��`����n�t�_��0R�`.�W��Ѣ�-���#��w䆭M�>���*zx��o��m\�S��E(%���2���,�Ջ>㺢.J�~�7IT��ACIVP�e�7_F�aY��>�T>�v�7�#�5%~tN�ݹLm�|�T�mk4:��/o�'��i�C�JNh)D���J���<'��f�!#��/����W� �B��m�qlv@��O%��	����Ty@���ۢ� W�{�Q�#��"�׌`�$-��
V��#�8��u�Fm�
�7C�_�縅�tS�2�*Ĺ��&�,���m�{��ߑ��ѓ{�\�<��f�=0hT�n�S.gE1p���	o�-�R�r�3>C�{O�K��`Vg+=@��0��`s=�iO5H2��) mf�t�$.2^�@�q��m�e%!�]�Ã��Y���m��X�N�x$��>�yy�(���<�>��Ƕg��ڼ��r�$�D��Q�׎�q�8na�oy��!�W�M����N?*��n��[_k�h���8z��|&��^f]���|"A�t���a�q���}���2�="1��BBx׶4�F��{��Pz����"�H�|���A��������/��K�4)�����Q�Y�}�����#�n~�ڋ�rr� b�]C��({���!�ĭ��-���� E0�K��2y�d�g-0�_�AW�p�"�,��.��w.u���vH�Z��߾��t%qk �С�N7l6Z{&Se����bTX#��Rt�72I
S"f[V�x^g���6�c���6��\�L���l>�\V�TwOY�\<�X���Y�����l�F�۔�o��M"���٠vHY䖊sJ�{�u�N���8 BJ,���D#�>����.\*�f%�1�#�����%V��j�Ͽu��J���P`)"��'T{S�`��`
��_ Z�+���Á�ծh9b��|��6/b��OG���{���#�ɔ
qZ�*�O遰����4��Q���@�Q@rb���S���1�D��3!�5�p�.�g�`�٣���]B����'*�	>�N9���ߦ����l���6�U>F���[BJ±b�h�~J4��}�Ta��O�[A�V�/�ɒz�)��v��Z.��I�Ψ[���s��|�iD��M:�+������H�����Ƀ;	>��&�Nls�z�h��
�B��s޳l$�%�9��K�mSvޭ,�K�e,\Л+h���w+2h�透?L�OӶS�7�:�c���������Ԗج��ڔ e!�3i�r)�A�߹5 �Ϯ��Ï��3=�؀�H!�=�
dLf�H�qő�2��ORb�K�	a�N:�l�w Cݔ��B��À�R��$�R���e,gJ�y�MA�44\F%������-1�K�x��Ed�*xHx�j}&��o����M�&�z�_Er�ɼ  qK��$(9�1k���s1�.�(k���TL�e��}C��P�C��M@7�@|,jQ�E���y�D�3��H�Lc@���n<�D_��)�dd͟W��R�Ŧ�F�HQB��(��|��<\��:�`�ᡨ��YH�h��E�yG��	�O%�I?k�BǺW��|RԆ�&trt}��������+������w�v��S�Q��Q���Y�(����XOE����y�\]gf!���\���8l��,�^�*��.QL�G�S���������}���u;)P�콝+3@@߮	�����I36�s7�/U�<�>�P�wP�l��a(r'i��in�h���ί�ra�>��ܔ�o��~�chxpn-�E�쫶��*� �F)�%�GhiXQ�A��{-�7�,����Ƙ5��r���������ז�K�Ŏ|j��7=��dmw]���9,&���DuB�!�> #�z�ԋ8�U���/��o~�,������(\�ۗ�hԨ��A�L�/^��p��U$?6f�T�S��d#���<3�oz��I��<��
ַ�e.��G�"b���g�_�/��T�ţ�8D}�!���?C��P�|C%�z��K�A��#�� \S�\�a�������v�輫ZC��y�'k�D�;��	x���PF&vXX��a�x��L��k��QKA�@���� ������7_���8�����.9c��������y�3���M2�J�&�h���ir��x�+G�t89�gE��`P�t',���C(��U!��aAT�>�vI�)���T��nN<��s~�-�j6Z];�D�'C���.���K��1w�Z�&R�1Gkm�R�A�&Sؿ�����;ɾk{��ѵ 3~�����);A�nWQ���OL�|4�1\����k�~�T��j�����O� �Wu$[KJ�?���o�������k  �u�1��L�c�&�';��ߑ������.5�h���:Q�s�%-��?��;]o����lIhNs����}P�
�b�U_��,�NfR��H�����'40Hh����}�D`�2}�V`���\����w����r/O��i�(��TV�ߖC�� �z�S;`�_��,� �8O��Cf�!�U'�=����P�{/g��	�C�	�`�j|J�N$���qnCv�/Y������
���"帀�y'�U����%�a��IR]c��w���F���ZJo�/�[����@���:�3���kL'���O�YJ���2In��cd,�o�ln�ڛr3�-��lNeX`/��j}�`�FZ�=�}�1�דNp��p)M�A)�ܩ_�x"zf߹��SCe�cnO�M�TV�wƔ���B]�4z�Am����]ulFf�;\�)26���X�ov�^o�(@��G���P�!��ns@�쩃=/FI/��Њ�op��>Z�Xz�ԓ? |��f�y��cxn0 |��H�܎��h�����'��׌�P|�E�������mu��|MQ���M���B;�I�U��c�& ]��Ԍ�fs@c�o��_:����Gx=Ad���*��mOj���[S�!��.@y1b��lʼ�v���㣷h6(z�+e%#�'���F�{�ev6�D�C;��5�K��yB]lW�����oղ?��7�p���{l�K��h��(��HUmF�
����40J��7@!�B��H����
]�f�#�G����o�|���{?ʎ鉨Ԡ[�-����
t}�%�y+ݣ�`�4H�VƝ�7lPhc��ʧ������䳯�Kڏ8���a�7���*ݠ�f���Ѝ4m��K�V��{~�v�
b�]��ħ���&𾏈�`x��Ax��&܌_ ���3���k9�^�y�՛o��~����H\���� ��"�(:}��tݶdJ���J���T�8ǹ<��s��Z�k"��M���aApךN.W�f�I4�"�g%�O2ܨ]^;�A��x@�4,UKc��x��ܪ8C��+�.�M2��!�H�&o�zq
�]4!V�����w�Wޤ���ݣ(U�a�.��V;C���4��$���ã��Gy>&� �W�cƼE�*M�k����Q�^\�y^*���uKF-����O��I��2�Y*s�}�l�l#A m_����d�n�j)Q��:�h��p�/8g'.Tz������'�X�F��nu� L�ܺ��V�c��ݢ�*L'���mE�BcJ�w��>&۽���)�ߜ4�RMfC'��y�ۥ�څ)iK�S%���/ƺO��G�*��uML]��|����4i�x���O2�R2�L*�)�"�X�}��HIa(ؒ�	1l��y(9��d%:�V��Nh��dp	���s`�
�F6��1��l�PpT�?P�cX>7b���gw��:�Ga���F�_��]������9�Mib{�1�/������V���_o=��F���7�0�R�?���h��84cHP<��7z�!�Ŵ\5CeQA�P��n�����\EnQl��?����ӣ�����D��|�4g�<S>�Q��2��	P褰z;]��^pb��vV�y�����M�:Ȼ�ՐQ���L� ��Ƭ�`��4,��E뽫C^n�6"�
���a<L
��2�YT:�]_(�R�	���Cs�7p[��rt��L:�Lxk��^��7���J�c�[J�e����S���߶��0~C���i~��y��a �#ZPE�Նk㕺0�G�?9��5xbb1�# ��⪖�W&����2b��1�F�c������� �Yv�d�D�=�J�S[����G����<M�#D�f�jd��j�A6�p���1Ɵ%��;�o�类������>:LH߱�?�DR����
����V!q������U��s�;���`�n�_d�l?m8hMF7c�c�ٺ�%5F��fd~��#mޏ]r,<ñ�:�y���i#r���|�D���*��ҧ�'�tu<���{���׀`��Jr6<G���j�!A��~��ȩv���
�_�hn"�&��Oչc��7�T,'G]��-������O�'�\�r��8�� y0�X��g��!�R�,���%R'a �'ԣ5G$�$z��`�7�~�v�х��F�hP����#���^h�ȑ���&��>�%Y�Ei�I��R��#5���	Ԫ�k*�[��V��[�qZ�&?��<J�Z.���W��V���7㉘�K����Ž��uj����㳬����n��R���}LfNE���� O}����q{G��� =��q���໺�ͩ���sݪ
K�-(��P�-d�1ܤ3����{��_b��c�~n]�֣�{Ӡ{�
�pѽ�x6�bп�r�����N������b��;K�jA�$��P���QC� �T�S�3g�Ş�}��H8Z���c&���z3�,����{�B�E�)Ҫ�g�d���#����hv�8�����E޼������V���)�"yg���V��<�Rz)�R��cF!�;ޫ��M^�2�8Y��x��PO����вw�}�ؒ�وnRl	��_��ֳ�����s�u�����б��U�¥�YBKR�hh���ɩ �s�T���AԅD�t8��^C)\�_h*;�aPH��Ⴚ����Ih�ң�iUknSh޷��U<��k��I��ЃYS�����`"�����P�������X"��ic4'����6�S����[���*�h:�>$���ֿ���T���I��1J[fJR��kP2-1��؜6�;'�sA*C>˺�:�(���-��p3~&�e.��,�~�K(�/�	��2���G��U�?|����"�F5���=�:0~|��m�N����.n��]�,��s6�ks�n���m�o���Ϊ1�> �	Q�[�@��f�lt�<$���%�l�q-������\��MCj �]�n@R<�>�8%�����f̷X�^�TLJ�xNF�ň�k�t���]q( ��g�B�EҌ�א�b�jJ8ֆ���
����7��n�S��m�	�ZV�E��n'�>�SKCE��Vk�] o`�Pd}��F�"�o��h�`��<t[m���Q�[(���||�,���;���÷�����h���2�OO�J@@�^��,	�,.,�����	�)�W�U#�u��׮��{!��M�ΰ���D�A P���F����d>h�_/��`�6R�e
���dH�v�@�_��ѭv!ZwF�a��U�>��;*��M�3Y(j���޻_�7=�S}��&�s�([Y�,Mz��;7��D4�O�������X���d�a;� �8�~�[�F��bH`G�vI���m�~'�uS��nQ���/܉��G��5�bB���e�f���V��|�L�N�zL"�RT�3{���_����H�&���@I����7��^���F�5[�&�{�m릧��~Ј�$�����;S�����ˀrl�f)�a9%K�z���\�����N�/��D0�qi�3�5���EI"�$i�y��i��^��c��՚������������-!�C����XIЦni��(�p9��X�k|�>��fo�O��z����,�Q��I��Ge�@�u+߆� ��0�B����J)ɘHx]%�J��')���9ڜ`���"���8�ݏ��c�v�š|�%�Tg�0��U��T��(z�m�0��Xt�'O~b5���
|h�Q�7݅{A�����Y�����ҫ���Kk�2���'��ɔk s~a�@D�8�s:~��.^���[%>[F���UV�@U�Ov햳�%/�� �OeygG���oVϏ��z=�A.�����u}�h����g�U�T7˔�I�F��i�h���Wyzt!��FG&����o�5���նn�w�4țg�K� @����"�s���/�!�z� �k�6�+
�XX�^��Y~/~�y3�AD,�+O�k���ɨ����bZ8�T��'.�������*��e�?yJKzex�%��5&:f9e�x��vy7R�"8.��M+P2�2b&��e���r|��h}?Z����/���T��d���A�1��q�L̸��-��c�߄jv��-����[t�c�� �����5z��G� �srA$���p��HK�z�n��u�g�����c{yY��NfB��#)}��i؄��8(�P]��t�W��[$��n�����kPnk�O�U�a�=������0��_��ld[�(Zdpb&Ԅ�N��T:����R��>V,BA�~*�O. "�F�}=������c ��b�m���k���4���7�R���JJ>����P����QJ�RcΙ��آPA|���d}����ʧ��N<����F�1����Zm�۬u���@9��9���F��h�O舔���w�J��`�e�.��|������#M�n`����6O�/�l��#����>{�/D��vP6���c�>r�wv ��	\�Ma������'Ul��'�M�&�!k�}�9�1\�p���w��,6���u@{a����=8ytJ\F�?�>D����5K#��L�Q�cg^(xX�~��5:�BA�����=2[���>�]ٌ8�ΟK�o�s�)r��Ƞ�Ԁ�3XZ��%N�RN��K�#��"!1�~Hx*�3~
��N�)��#�k���սȶ���,^��F���&��W��z���b݌k��?-
>��hh��}Gd�d�z<�4V�WL�x%�*ly��[��\Nƌ�v���=��f�lp%8rB�#�[2�=�r�5DB p������T� �.qc	#3�WF���d���=)��*�[��S�����́�H7��'�b�4k#�N0<Pe��VYu�ۄ��/!�?a�t��2�4�{�=8�����ƽ�v?��u��MB�f���ڑ7��9��\�"�w)�̀�����K,�+,�p�]*IEǇ���Y��p��Ql�3#@��5�*�K|��,�)J֨K\H��J]��O�����|m�>��"��Cu�<������!�V'��6n�n⢺�ʇ�ݠE.p��Ǟ����v�]���lw��J�w�ߗ�%�I�2�����j����fsV!&��YHJ�u<3���h,�NG-qh��|�y�	�w�}����<ET�|����,�'y%�7�A��~Z~���ꨨ��é!n&�X��\S/�I	��ڻK&�F�,&�"h:��hH��CL�ݪI��V��uk@���_&G���Wk�$ݠ����͢(7�;�H�e8 �k��\�h���o��F����i���h�	����1�%=O�̗�n+
`��7��aAm$sr�R�l���;zf�t��B5W3?x7c�[_��!�K�Еb%qFO��3�7 ��ﴵүK`�n;�_���O��r�j#6�x����:�*�=�l/o�q�m���-r�����nhbK�3Ф����-꾝0�HQ"�Z�q=#��9�E앫��']��� ^ڏ3*	-���JS��j'*k�99��dK�~�u"ɭ��D_(��%�LmW�'�&Wѹ'{1�>�J��'�%�z�#U:�Y�:���������c�S�H��Pq�B�����O(v��d�9�7�G*ar*:~@K8PH��M8�!Ɇ�_��c@��m7aL7"�2��A},C���5�D�4௞�a�T����5�(�}�ʵG2AI��Nu��X�i)���g?�\��a�Q�]�n2�9��I�+u:;�ǬB{i�H��9B�B��r��-t�t�)P�f���ib��c�cao��<��?���s�S�����@���Q� ����	KJ�F��$ۭ+� ��֗d�d�
ڇI�'ңohMg��b���3 9TE�-��Ō��o6��fP�R�oÚ8�Hm@�劳�&��6C �p�T�e������#��ڽ���x
��^�2S�f�>������_�چ��%��������>�~<H��ǹ����|uJl��}O�X�6�� ��î��]Pq��7�r�m�2g�U?����Col�h^���WES��������MU��
>gO_R�����S���h���g4���\�0w�7�Ʀj�W��K�M.r�e�j�L�"T�o�����X2+�wR���@����r�_�&q-�]�>n������+�h��X���~ Gc��{�;׊L��A�h�|4���#�t�7$���b�ѭ��g�~
~i������P���<�3��4^���ϨQs5��!��k�|��9���D8����1]*���(@��j0��PO�F����}�v%�r�z��� R�"��@hz �?|���M�!��3P�M~�Ƃ��/5�m���OmZiP��Ql�6�b�a��q�����[|�iv�։1���,�2�|o/�ᇑt�L�,��d�(ʜ֡�]�b��}�!P6�B��1e������˦�� la~j ��AtB��0ݡ��z��͆a7��`^-�T�k�{�>�-׸A��MJ�mN��sUx�Q#2�܍��J	�ޒ���=P緑U���/�%E 8��U�]$Ϻ�> ����:�i�Wt��d��*5��<��3g�Ê�p��<������Ix���im��5G	SE\���B x�!������5ͬ	�"�������'e*�1+l��}���6rҧ�g��V�^��_;�o^s��[�r�n�=��Z[��u<���ݵ��׋Kf��C��C7=صML�W(b�'!���_oDCd��{��[p�V��,	s[�ke�ն�k�{]ei���-�s)m�0mh:Q�`�0r����>�{��bƥL;ư4�q���i�O�r;k͜����s�̚�ň�`y�Z����\!�q.�j����aT�1(��K�q����[��c3��pu*�?ɒ�)�ŀ���'�?b����&/Mn #��g�ʑ�ꯋ�^5�8����t���~ �?|xzҽp�h����B��҄*��v��hv�D�B��nOV����8=(��2�O�9�����S��D�d�d�Y&ǃV�D�+|𒧔�3���1���RwUe�"�s1��`���V�M!�w@��N+��'�S(m��fU�\���<����-�E�_�K�LI|�-��ܱS�﯅@q���;�@��n�1�
.�jM�pDL6��8�"��|Z���	���{��?�?� ����e"T��<�P�h�-[�ͺ���G�읟!������%����ٶdx�T�Q2jc���n�!շ�b6WbDh�2�Re�=׊/�q��|.����� T(�cQbg:��~���N٭��e[o�͘��m�U����u!5�haUs���?�<^7�3hYg>|̷��) �DV��\��#g4܂�cRzyf�yH�?"�w�w���,���\do~�ߑ������c�ٲ��)�Ϡ�6�Z8�����P�Q��Wx�_*?BC��IT�KƷ!�n�@��'hk{��3b�Ԡ�L��q<y�J�3B3C����g{N�G����j1��i�&٥���''�TvOI;��ȿ��`̴���r����*34rw���P�7�!�8���*��F���7s���Q'ö�Hj��q�����H�2��t�^�e~I`�O�� �`�IIa>t>�Q�]Q�3c=��k�qA�"�Ű�f)��/�M=��d�*D�ѭ7��B�o��K
��/�,��CF0/�$&)o�� ]�9k]\���$X��sIy�p��(��5�]M��]_ɬL-�egӞ�P������#{��@v��J#Tϓg���݆�� �t�h���u��R��V�Ψ�[4�J�»d���d�9�7�L3��`Tx��^��]eW�Ƚ���*��=��֟��KsS�u�^$9u	��&��Ų=݀�^��ɬg�
dU�m�o��r[@���&-�x'n�/S����pŦ�>l�Ҩ;ٕo���.X������D0����@v��?�ۈs=Bt�c�v�2C�)v��`���X��&f�q�����(�� �jc��;��w��tR8�#�F<���MEǬ�}yb"~���޿zL]�z�*�v�nWeu�ށ&K'�,���般�@����fLx�٘��$,��:7(e#mks;Yy@���j�Y�m��)� ȇt�A�il\ƲÞ�G�<-�<
Q�N����Tvڸq� ^���x�ݓΦx�Dv1��E�qwFԍ�:���ҽ1�b-Ըbg���+��K�������h�"�p�z§hR��G�,��r��!�!�}P ���/��aY�����p0��'J��J�W�=��۶8�?�κ�GWl�o�b���Ј��.�֡���	~�%�u}�-4�\�2�U)ي�.�Sю*�F���sN�wd�7t �`��w�Z��[�E��=Zh�YUx���ἅ,�R�3�J +����a~h���L�W�8"����9iŜ�6�)����[��ofk�2L�??�U筷G�����F�ǧ��� %f�*��wT�E9>�j�mZ�Ø�5�w���O�e��M���%�� ળK �
n)�U�z�jg����x�CR6���2�Q�����ڰ�MI@jGť�����{h'琽�},�6a/�\���
r-{ENi�B���k�4�@�M��za�ہW�@����@U�b3!��chFl�io@������8g�K�_7��U+��=?�� b���e�q	�O(���/��sy48G{��Y�6�	����I@��}� �����P��p�$�D�Ł���x:���=����w^��.S���A����l$UBU:/��Ã��d�˰l" p}08� ([JC��'�c� �ğ�\��%�<<ԇ`u<�!��9ff�Mgzl�Z@p�S���aS���)a�><7?B#Y42uJ���Hc[3�1���v���F�����@7 E�]�Gg���f�$��p���v�f���~7���مġ���+���m��<L1�P"C���=�o70ڃ�5B�0�V�<�`j�������&1~��e���YI��v��n�]�:tO������.e��m�|�0	z�`~�"��3���*e��J�;�7�G�B�W�y�	��*؎^��z�+Z��N���uϋ1.-����d��X���~����2J��7T��<�Ll��J�?�A���$"U$`��������*q��fd����V��PO4%B}�2���������k��v��D?����i�ЙGі�alB�	'�R1��'-�[ �U�\����'�j�s����Ne�����V���n�p��	�B�td�LC����0�h�>F�`��6>�;�6/��j�zUzw�e0�2���Pb�l~La��5�Ү�B,/5GrN�pUr��@��Ω��T����Wj��]E(��s�ʦ��ܳѯ�A�)x�/�]�gl{��Y�ͱ�����Kq�xG,!��*�mm��'�����t(e��2	B�i��W��5k�=h.��VL(�\�6���p͚�F��s�N����Qc�@��Cy����ՀW$JYg�1o7�IM���4��yY�oƄ���8�u����8W�PG���U�~3tUOm�Q��揪ğ;��n�k'��P�y�(��D����9A��h�o�Q���������'��#u�l���؜n�7CQr-��b�-��I��;u$/���L���`�Y*���&����Xа��|�;��1���ɶc�blr��-������h��ݰ&*72��{������T�睙������Y���4X�U��lQ���1=F�d��k�,����D��m1X���h�|s�eVFt"�A��5S�y����ۉ�������M�R�_*��k/8M���)LF{�1)2�]������bx�uz`�Ccl7�.�5�P�-"�"�����B���&h�K��o����ݪljoS��.��5g�K�K�3$˓�G�
t��{@� e{�!���P��|lX@�z+]�3�9j��M�M�����z�?@f@7����O�@�.�/��*t�z|z@� e����bÿ��'a_ ��9�m�\��hO��zNZ��#���閎CyIn�8�����R�@Vx,��^����q	�y/��a�Wn��Ҟ�.<�8�ݎ��F=�S|�Z�Nu�Դ'�:�ˮdR��wSC��ğ)�F����F[��,JA	C�y灻�+��n��m����E�g�B�������K^9jvμu�GtA���I�'�HZpN�KŎ��������"������e� n~�I��Z1�}=�2��w���aǠ��B�qO2��m���OC����ų�զ�#l��
THf��]"B֝�А�h
��&��c����	k����6�`�H��;�*R	���L�����j�E�j9�[*�k���s������$�	����㓯����5��?3Rf�HhJ�̗#\��!%�k�'�9���_^�-�n���Z���0E-�Yo� 楧���E�`c�\\j�-���a�c�Nd����0�uNt���~I��ط��Y�^����ozP$v0c�;��Z:d�N´�a�i�b�Ƙ�9m�'�I����4%_��s9͵�an&���4_ }�����Êk�|�k(��܌�O��u�o�n=�������3tG^�n��G.�(�c�^�y���5�e/gx˂D0�֢eY�7uj�6ު�Q/�5Q��Ң�s�o?n�.��r�L�)��8��ĝ\|��^��Ā�:�0���߮R�t����}�k���]�Q�n\�1žb����D�V�	�n/���W��N�Dy�y�^���t�}��E���}�p Wj�.D��b���#�w��J���jQ�v_�-6����(��	�I��m��<D��bΈY�A�ʽ�]JB ��>Z2
�J>�s�젒U��s�����?�c��
�ILC��o�y7��n.�C��,����x�w��T��%4�B���_�s�t֗SC�5d!�0�\�*�P��C;Ž��5gC���L
Uh�1d1q$��	Xz��[�m ����uٯ���p�P8t6�wq���o��F�����*Y:�)��)����:6۶Ȧq�����S0c�.�eU��{�P��HW ]D	��m�"��e��HJ\�{�X��!9�0�}������K����gB���7�s�o�
#�Q�pg��2�ރ��Z�]�V�a@��r���vG�]I��`��Kи5wZ+���S�=�<����|vh���07�MBZ.Ѯ#&��ͅ�k�+'�T���p���p<�`"�h�[��.cБ�����a$Cq�F�C�@Ǚ�si_�k�T�D\]'U=<d.�#��&��_��V�v��J�@�k���	�7;�jyM?�>��̔٘3pH;#���%�(��c��X�vn�������B!�?&����q�te�s+W�a$��#\�Ć���T���?���HGw2e�ݪG	�Ȟ�
_�������=p5��`�����Z��̸�xZ3ً��w���Q*oV���s'�>��d��P�A��z��M]�g��YfqP�=�p�-CaS�d��\��8q���L��2Ǫ�"(�҉߿wdAk���R�ױ.+��ʡ��~�B��f�a����)�Ү�\�v:�C`3R���1L�R9N�'���E0\��j��6�W�F�W��立�D�e����ȯ�T����*=�b@
4hz�����]:�����1�Aw�&�o�Q(t��_����-y\z&������O!:I��@�����J��T~��Ec�uП�X�t:��2(�A��-R�-�����-*�u��~�B$&h)����G���5�C��\�R������DF�UW��\K��^�b�9����"� ��	�D6Vz���L2t��3�|��zM�|Z�?�������r�#Ħ�T�m�6��e%4%C�P��p���hl�/�Z���e�t�����z�� F�˕��)k��Û�^�o�O�'��Իw�}���ޤ��hY'
V��6��-j_VGh^\ Tf�t��y�����3#)S�0�㉚4����7p�qeԹ�h.�d�s���'F7������(Phd��Z;��)��8�7�O��ͪ#&R�z#[��wBb9a��R55��R�Jgy�ae4�iA�v�"3Zh�y��1���UzP34ܶ��).�6zŇ�&[9�0mE��C_�C�S�^��	a���ȏ�k�%�6�F>Ww�7m��%�[>��s���,�_��o>�f) ��*ʉ�jN�-
h����SH��勍�bT�������3&��ڐk����6{�-�IYnyk�\	rx����#Y�Xq�S��K<�T�֯�?�TD��{Q�KO|o&�p��Hk�r.�N�X�X��|w*,kkAq�肁�}�@<Z�g�;�M�'�in��6���)(,�3�Dٚ���o7�dʲ�1����>L>-��ʥ�x�	���W�Ih�E���+"&WYm<�Z>�TK5�����T���k��<׾t-4�����?J t��J�ZC�����L"M~N�e��9�u1�*��i������4� ���G�=�~������)���7�p!�������LF�[ C��Ï�����_jc�O�g>ei�	NRPq���������v�'h�-�x��)Q�K&(�
�~�7��y��ѵ�c��M<�Ȣ���V���׏DS� SH�����R���.f�H܆��s�Q*'�W���b�ؽ�i���r%U��ߗ��4렿|׀V�i���ߚ��*Y��0[~3������vӺ�,��^�2�N�C����=Ff9!�R��-��a��O�ſxk��>��'4���c���4�Fъ����jc�}&:�0wd��w�������t*%2����zZ�I|��?�j?�w>�)��ש3\�S��M���;��
��#ԋ[�T�ݡ� ,������L.M:)�'țp��V8��#Ej���A���19�4x�bѢ?Da4Kc��b�xE/@C�0�=u��N@�$�Xi +���kA�;a%�q��O43���h�բ�J��K&YsM��0���׮3|?���E���:�ϸ��w��ǢM4��Tٙ�W�=�!o����� ���=�I��J�Y�-�f䉣s)cɩX�t�_ώi��e���%\�K�z��'���L2�ћ�q�в���7��W���'Iّ|7��������)9�8��������ò��6��r�:́��%��BO�4N*��������p�|r2Bf���)ƽ����л�I��/as]YZ�z;ߚZ��M(|J�z���÷l	F��C��#w�9�>6�E�A��[ ������s˶�L-�7\�����J�=��荄�_MȽ�՘�����˝BC�*��Z��ٙkb.��l��-�>l�jOYڢ���f�A�al9��'
8z`�Bp,��tY��n�b��?Z�+ܩk/e��Ι G�UE�o�Y�ӛ� �2<���Vd��5Dz��]?p�� D�����\HeT����
x�����Y�4���!���-��r�6t�J]f8i��D�"���튦aaՠ�9�=?�e��L�UoH�G�pu ��Xhz�e���O_���<���Y�~RH��2�	����O9ZRQ?+�P;� NG����D��7u�hK�1��{`ô�ni��T�������%+��i#�c�N�e����j���fN����X����W�q�+;M�-rL�7 2�Atj��"1*Wy�/�P�Hn�����v���T����F�p.��s�	n��lnG���ǟ���t�ń/�c���l�8�~�mݜ��x��g<�5����k��7�j�F$s%�^}�4���>��xɫ
串#qƯp�F3�������YN�]�����Ƈ�I���1N�2~��2�@ ��>��cR�69��MK�e�⿦$cS�){	5Y��
�9�Hf�VԆe�y�x���ѦlI׾
TS��T�F����r,f?BO*��U�[�q-?�0�!����߾0~y����/�����l����"����*�;>O߳�uo��n�'@��_�g���� �"���r�k8���Z3�20�?���Km��5b�C�ih�	�����	b� � ��+<my���U���(����܎�
���Mey�P]
0z7��kb���p��(l�:�yh	�X�� ���0J�������k�7̧�P�����m{�|������u��{=��S����J#9�"?#y�õ��a qSR��g��Z w�2W)k�:�!=9��=�"�
�!�/uGc�j������'��"Ͷ}�F������oj���q ����I�꒽�|��W�p��)����H��E�Tb2/	�y�ɯ���/$��wC�Uᓱ̜\�(�~��I�e<�Y��#7���y�����<qY��L�Iu�M{��QS^����devbv���b�z3��X��-�r��w���~-��Sɨ���Jng�2��̢�jt��v7��t'Z`YO*�A���r �������>���w�=�G�M�V@hvf�!�� �L�A���v�A�5����*D)��s\|�Z�_5�ĢT@��w�l,>�F~|�|����<l�P2�4���7<^�<�&A���a�P�F?��*��lm�&�o�*yG�%����������Iun����T�%{�o2��˃�ex��^ D��uV;�j�b����&��/�{�<:-!R�H1Z�B �3#ӌ;nH�\��U|.v�zP5�	;<߁�1O��er�o��h5�F4��DF�b�C3�5��o]�#{Y0���ݏ�^E��}~ћ��$��:^N�$o�$�_6��͕�Z����ڔ6Y�)�'�����v �'����Y;R�\`��`�1�'h��2��y����,�m�ߝX���/�5=��΅xƍ���|ި.0+� nxla��Y��{/=��0�	�}(�A���Tv@��X��[��|��8�;�H��ajO�G�
t"|S���'ٺ�iu�k|8E�E�d��lGdQB�� �h�_?�-뉼�� �x�?n����8�_����W�BD !cZ#-~�xF���z��1oEWf�]/X����#:�Y�bb�2��q�!��Ɉ����{�}�hc~=�:��9�s\G���+�_;���$f�r؉>��8M�F�J���P�6FV6c�B�R7M�]?f{\���4�?g�߼N�W��߶���dAC��[��L���o9uy�4�0�bP�������_/��D
1�R�D�H���Lk����L���h�{`���\`Sl5���d��t��֏JR�:WP.R�EOb*���c�����k���%��-�6	�|k`u�6��
����J�[dq���K;P>^��W��^<3Nv�.a��y�=o'F��6��Q���[)L�,2�u:�4I2߱~K���UC��@��x~뺾O8k�2$�k�~<X��8�
�}�[�.�����%�n��Θ�P���n�y���v�v��|K�C���:H�t��+��t��w> ��*oC�"yy��Q�X�S��<'m����V#9������q=G�Y���������o��� k*��ȥ�J�� =e���73ܾ͐AY8<_Z�:Q[
@>�}U���~�Q���S����`�lNGq��קƟ(k�����?�Mg�wn�2Uʵ1vP�񀟉%N�|b����ObE퉜��	c��ə����3���H׾ҁG��$�A��Z{��)��B$�`�G��4+1�#��qŗ<Z��}�����5�k����A�L�)��f����
�% k�Ɲ��%o*8Ѭ��[�Rmt埫"TT��[��E�k�إ���duW]M2���(_X�A�͏�;�=��Hi~�H����n��+�9���}���W�����t5�}�٦})�dwA�JA�w� 5n���)ԍ��S��{/��{�����0�3ַ`-���\�����!��|U�h)�K0��@�ǀS!LR�B���ӝPo��fR���h ��ɘ}&�f��cΜw��Z�sqf��KԢ��N�̶�5��\�9ؤ8�9{}ڡ����C�cÔ,�	?s�����a@�i�=��ݰ���{�OLǙa���7���#Gbm0
ևM/~^�h�\�7\s��=�4��|gh�e�� ��b��'E}�;�"���2���`KR��;Cx�V&����-%B�wU��+�8f�G��|. LY�[��Ӫx��9��m��u�ib���W�K�r\�x�@�=�de��kQ�p�9!
�f��n��")3c�ͼ�;sru/,(��/
��ɠ�FS�	���8f�"�Y���y8#��wr�))�X��`S֮�ȹ�//o�7Y�o���Q�3��(�s4?%+���+����u���S��XY+��(���93�������HBgP:�l٘�,��Z�״��/0�2��*Aȕ3����)�5���a���z���hd�=�yv���8�P����On���{_�����pv9n(,��(����	5�ن8ϝ�M������5��y���.�H+�e�M3��ܵ��r�����x<�MbX~�:�=߹�+�I�_2�>Mȱɬc�65:5���!��1�*Jo�VC��
.�VPp���MK>�&DRf�>�)��R���-b���b�Pi��Њ�w����BO�e�����)�٫lˊ'
��.��~��3F��{j�m��%9�'�oK���y�oK9�`G��1���4\���=\�$��=)X٬!ב���b�u˛S,�"�����鱭��J�O�&�Q�r}���Yl+oJ(�]WC��H_d^���՟I$[�̊�[�yz` x-�e�	���I�����wE�z�2�N`�-l���|�iT��A~"ȫ�Zwn����j �1��X�C���'4RkxJ��Y�bgu"�t8��z�;�Qgp{�w�_v�z9����n<o�j�iG6�?h�xl�D��p2Y�\��M��|sj�y��j��W�W���(c�+�]?ܜo��X5� u�|��[Q}x�K�v���L{ð�;�O��yw�����%���~G~|�Qb�+vE)Xrv�I����nO���Cj�nyO���'�9-����e�
:��b��:°�� l=��-�L,�]�NV)>U2>��P��0��4`\R���WA�>���-ᷳE�-[�,���:��s� �����M�wO��O�M���9��#:љ�#oh[��ԥԺ�<�Rs� �򳓅���\��dbE�*� W{TG2~<�����.x�v���HP�����gr���Q�ِ����hI�u$(�� I�M��J�C�-���={F�O{��@�`Pp
� *����������6�Vh��ѯ8�?$��5�F�'�:6]�F;�f���`b�ļ�(�_YfQ�w�;}��el5@� �S�����h{xwyg��D'8�]�6��!�<��j5�~3��J�b�f>����6�����Sߛ�MX"6UÃ��v"�C��_e)a�Y%�p`_(d��A��u&1�c�n�4�U�H�Cɟ����6R����dV^C`��E���'�����Y)lF�lJ䀋��y�;d��n��9MJEX��B���q�uz��<4X����.�
g�gf����������`�C�*�,w`C6U
0����t�I�D�ڬ�|�t��܃�]}r�kã;�9������ҝf��PKh�R��K@�o�������_4L3fJ�x��1vs�����2��e���)�׻L�e����O4(0��;=�Y*-`���V龦:*���1/�%ԁ���
���m#�^�9�ZE���?�(
�IN�(}[����cZ����JNd#�l!K��]�W�"j4t?5oR�&�����2~��F����X�%�0�J�C���t���u�I��~WBQZ+��U���6_��S"����ឦ�����h�{bbb��v��_ ������o/�@��W�� �e�T�(�l���G.B�b��� �K��`0�̚]���Sj�0s�J��*���;v>���i�eW�&�|Ta [r[섢����y"���!X�|񜴛.~���4�,OX��ø�_v/Ȯ{׋f��{}��Z:��aY���o^����~��C�(2�Z��Y���?/M�2R-�͒c �w~9��8�Q��
���89��Kڶ������$6�##�GB�Yډ���}z@9�{ؾ̱)��[�~	
��d�# Y�\TeĹ�(?w��5ޑ�8#��z���P��d����x�{S<b`5Z�H%��T_��2v�@���8a�<6��PG��;�upÚS���K��]o�dwd��Q���0>�4w!l<�} {��� G�.g�M9���s�3��y�RPU}��F���! Ѓ8�/]�����\�ɸp�B��V�eXRF����1%X)�Mԙ�7�Q�Y���b".˘�?#Jދ��Q�r�s�c��s�p�����N���w�k������+Sh���@?���gʜ�����|zq��7޲P�#
�	w��F�y��`w��{����4���F:L��^�����mr��s�>�+~�<��2����r�n���7����+)��?��V�(�c\ϼ��]C ��]�!��p�Afȩ�,��~-e�V���l3V�HQ�~m�3����@����Ϥ���=�p�}s���#T��a�	��*����Af��������ti��;�y�����w7<��-	�Zѐdp��7����)y�X� �Ю�mƥe��rD5n;޻n&T�T��C�p�Y���(��5�*��:b?�Z���uX(A�ސ@ڤ���4Ț�����ZnE�����̳�U4��1V�HG���R��3�{7q,�Dæ���z�yhl�R��Ӓ�e:�}�L�+�S$��O�|OC���/ld��0�}��8�ʴu�42O�<6�s�aFՂMX�ų���W�٨�|�R��u/=M\?��hʻ=��U|�H�&��8���2�c:�L���[����.)����߹ߑ\|�N�yk���r�~W���}����*;7LE���L�"���d����b�B�SQeUZ�4�<�[&���F���AXP4/����~�p�K	����G��(G��
n�O�m!C����Uv<}X�у��W���1G�"�2�s"~5�.w��b@�r�jL�ձ�̰"ӏn%�t%�0{�ٖ3�H�=5�j�M�;�	�$��>�&v�;Yr@��4��F�=��q���KId�p'ٵ��Ov*f�����'wŐ��g�ԬK�ؚ_:w�V�������t�k��V�P]�~� Se�m�W�~'�B�ix���Q2u=�o��oS�NXi���p��D)3PB}NI~�\p5�2�W3x�P��u�-A��_\��??�2�38�y.�k*�>���?4�3CsoHWV�h�Į��$AZ�t2������iG�����]�\^2>rd�����~`hE����	���Tr�G��>h������U�"��ّU��^��u딄��ɓNa�z(��l���}���b,E�hV23D�k�������}&9���S�+�-9]�Z:!���1�u�q�	�G4�B�qZ;`��m��ܑu:�U�����&l},��6҉�����L�	�l��+�����i�5�!*�O�"��XT����
^Ia%�d�>]P[����ԍrH�+_�fj���.��Rrw�w�2�~_Y}(]Z�{���*��W�Ƙ��sz9�Gx������jV�h{I��zd�wT)���u��32��*J���k���;�)��pGߨW�XK`��d{��:=�@=��b��B�8�.�X4�n�I��u'�=�\I!$=�EwJ-v�wU@�@��ɳdN���Y�RtY��%O
���C0��.��l�^���.\�~����{y��,���B[a�5=rB��1���p���:j��s�3S]!'����X���3ւ��v.�FFl�=t^s��
����q��1�\����ߕ9�Ω�Nkr�^�&\��d�6ѯ���NT�垨������t�Кy�Ei�푠���� �}$bl"?h�ٚ�+d{����w�Σ�:s1���x�ڐ?�X��X;�8��փ%K�du�m�U��2��嗛}�l��1>�L������C���0gP�YHh�O0a5�f��7����Ӊ�R6�{�{�����~�˥��+p�ZR�_������k[�w`�tAo?�H�� ]��Y�M~c�t�4�Ϡ��-_������x��̪}Ur�i����!,Q�#�~)���fO�k��`N|��86J��;ۺ:-�%q����
��i^�!O�ؔ�iLiC2��"�6.�eٷ�v!^b�9�%��)O��ђ������4�f�f���ʡA7���Վ�0012��x3&w����2�a�V"����z��(Sh��C�]T�@n��?@�v#v�����>;�w�{|c��qqq�:�����wz&i����y�S�e�;h�V�t֒J�k��e��Qb뼓 "�2W/O���G UNw�캛}��![��2[�����g����)�L7�h�#9�����S�^���V��S�_F�'��wkˍ�ܚ�5�Ҿ���'PK������\5�l�"<6��B�Fq��1}l���ݻ��3d?>�͕�ֆ=���J�x$6	��lA8�>R���`f;�l-ϳ�� e��{K�Q��\G��u(��/��>Α�x�I���?*ib 7ci�Fc!	����\�g
�H�YT$�ǵ���ۘ
Kv���yej�P��=��&�Hp3�*�q4$	�8=y�&�}e(6
x�lw�~���+(3��j��_13A��>|��9��P������~[�b�9'�۩,E귊�{O ��Wɟ½s�K�o0(5D��Lƻ�ָO�k�,X��s���GV]�	~��Mq��v�n�#���/�Hx6[-��<;ߴ��垟��B�G����&���3�A�%(g.*���j�l�iP�'������f��K�fo��9Q�3vުLY���8�ݧ��c�+!q'�.)o���5�]Dܑ��7OOAsOhb-'��q�/o�-����\p�+t���˃;ȷ�&���{���*°)h�Jc���M;~^@�?��l��L���I���Uj�աP��
L�x�H�	,��2�1�e�U����4��QIC^H%����LW�TOZ����y7�NI�OA�_^��0n\Y�>GnW.0��v��E}6�L!�Q>���A��̒Q�z�����Fe]��uۋu��K!�h��%�ղ;�G��F�l�1.�k�=��0�{Kw$�X�>A�M�Gi�W��sgݨ%�c�q��[/�(C+ [���K��h4#��S���x�1�0O%��'I��gV�W}�������T�3`P���[j� ΀{Y2�XDOV��xt�y���z� �%r�)k�w��v��<L�p�a4}�
��u��=M/n�nC�\�Vؠ�i7Hg�93����Ѝe�	r*�$�������iK����z;C9��$�� 0d�a������Ce԰)Q�/�Ї��o��.Q��q����]i��z>��V5�y�y�4gB�J)�	�|]��,�x#Ug<��W��.�����^�E4�8�O�D��ն)�ߪ��ĥ��xo:Lϛ_d��;�,C�M��CONNB���C��+��Y���^�X@�#ɼK��J�����>V�������¸lr�������t)Fu�hlm����#�����E֢�7��<U�yZ'
.��Ğ����75���9�.0� �l�,����zXu�i�<�6�y%�����}�}o��34��ĭ%��<���ы5����;�+l"�6$%#K��p�#,䬬�$$�q���#����^�h�C��k�OҀE�'��I�����ٌޖB���ŗ,��FęP�D{W���O���PVj3j�G6حy\�����O�h#B$ï*w
KEdG�"˶F˓�f�5Z�����6'Ɂ���'o�����d��D��9� <S͟�����`�p�h�l�t;"�����57玽�,Ǒn�DK���o����J ݹ/��<�1C�5̷��LZ��6�H1���������`2tr��s��Z�}G*2���,b��<���:p���9m:���g��)*1�ր��H�����F��]�h��E�|��"|f�a�=��k���Y��#20Ա�#�Ve[8�et�w��B�\Z��p�����N���
���f��0q	��O�g �Mw�sC\%���86a�u��f�1��t�ɻ�lw���<%�dR>��a΀iׇ�Y�X;���I����ޒu��[��H}�Z)=���M�Q��N*��59~.X��ס�c�T����
���T�'b.br���J0J"´�a���C�e�l���<>��DV
#e ���,��hO��ä�M��S�čx���}�O�}���ð~�8"�| ]U
�|D;n��(��E;�e��
���
ܸ�O�:�J%�$̹��e(@Ykэ�n�a�̅�C��ə�^g\���R����bp��)��=�G�
^h���g���8Z���r�!
"0r7�
�]�4��m9h��&��\<���^:ʔ���V��'6q���޸B��:�{%��@7}b���� �meh�_q��I��B/��#F����@�IKdy�=���ג�<�{��E�Д�[=�b�F��5���<�}{"�]��ā�y=�`H��+�K����
��b�� ��e8)�;
�9/��#�? ��*ӯc�}�#)(�*߬��C'��,Ӈ,{[��1l�E��ޣ	�L�ߒXL_�e8�>�5�C������L�Q�(�C�C���P��G��;��h�O9�Jl_r����Ƅ��I�Z��v�ʨRr�W�ꗬ�W��;�[�z9�xbf[�Q�T=�~�d�5/@Z����%!�ok�GtE��H�ز�0�#�L��)�1�g�*.�n���k�������s<80x?b~ی��䴾,>��Z������>�i���=y���GL��E
�g�fl[�u���f/E�f����"�qo�kgQ�ıv�N�����<�MK`{������@JkO�V�+GG��2A���sɳţ�U��q,37���g������}�Xjx����`���B�L<3]�r*�!�T}u2'##�vH/oD��R]"^)���3j�&r�)n����G��2C����\�u'b�'[}!\j���&�B���_5T��G���������_#Zd�=6_��� �ک��>���5�q�r��d�b�S"ڐ���1��λըp%��V��u��r'M�s%G������ۗ�m�:���%���M�GinT����9�xg�	��u����o�%-o�1xG�f�A��@�f~�vosl'ͨ�\�RU��	�n�h����<��ږ`�v�q�F���`�tmV�@f<�����ـ�`Иt	=�K��{F@\Q�$xZ]�@�Pt�9,'$л�@�W'g8���j�E5�嬢Ɉܧ؂A���N���1iv7(H{׼�V!w�Ѩ�.7Х���'4ǿ��M��
zW����-i��2�'7��(`��Y���Cݼ7���;y'�r�-XQ����;��8�DP1��c��U�O�����K]Q�@�%����C{MM|�+�̝M���.D�+}���:�gPg�f��#h���`e�kM�*B�O}�q��X~�����D�D�1�T�J=����i�Gq�����*1�����B��/��%��Y�����;�
>�����̠�Ml�T�x���������jv�]�hl�^�(���Yj�x�
�?��:��Zw��a=FA��6�2@���	x��|�E��J��a�n���!�5�钓�2��B�NH�G�L���h�]�QG$���ž�irY��%8�+���� ���\p$���(�ѳ3��?���X~\%T�U@��=� yMc�N�N3�G-�Dp]�
�S��UZ��z��[�K�qd(�� h2j�|���s�Ñm���'�@J�>�F���*mZe*z�LP���z�����[�֟Sl��\sF�H}N�?u��N��-�M~��Oզ�^���I��@��EL�59!g.3��b����*R������aQB��5?�I��ɺ�@B��ͦ�
]��1Z;Q�[��Hم�Y����)���*�z���|S���)+�:�G����#[\@Yy�T����)��%&��J����K�����a�R�!;��Dʣ��a����^y4��=����i��F�v����{f�ƌ ��h�*X}%�]s�_�0|6Ǎ]_����}���Ƌ=�VҔ���C���\c��Ɏ�ZE��_y��8vY.w���/��E�H��H""���cHӃ���y���+Gu7K�8ӥcjy��b\o�M�]�ޑ�z���4���LW�B�<��xuT�:�&�r�``=c� Ns���P1[��7j�_U��=[<���Y\~�폫�ϡ�M'tY1A�u�P��X,�I-�C��> # �Gz!���-����UjRML�O<��q$����Ћ|c�b�{��HC���'M���ߪ��흺9b�p(Q?���-�� �Wn īf�����q��%32����\�L�7qiɳ�.�;�@֗�n%K:���w%._�+�
���۲;��h��\����Q:���A����cw/xLLޭ�o\��Ã6A_�Z�M���]�ǦF��'��FY%��N ̸��ۭ�@U<	�|�j����t��HWl���tg�<#��0N�x-~8)R4������ϡ��%�+� �3����l�%���u�(�"H1��@�#`�b�{�fa��N7�7H��������$�?�g�	�9���� ��$��Y�[��b���@B�6��)"���gS�!\�
/�~�35B�]�7�u#���AWd1[���ī��*W�@�n��9�BuI����?�;���b�Ŵ[���**�<�e�3�
 ۇ��7.<���y�D�\�n���@=݃������"V`�z��;�"��2;Q�eo�H��}У���;�7�^ZЦ�$�	)�������<�[��Z�u����ݖ{��/�})�Z���J.W��#	�|5�;�I�*�X�)Qd�s\E#�P�2��mW]��ɳ�1�X$y�іs�eʁ~)�c�h��r������q�o�-v" Cႉ��@��D$�V��~�6~i��C���ٙ¹��1�"�f1Հ�w:\�+��wyU5{rod�Zԡ��R۬���/, Zv ����o�_��%,�`XVSy�=���Ip��Z(�v2�V��6*�i�9T>s�Z~���ǉ�yH��a�e�
 ?�n�d�nu��a�qq�jDDֆ�Ձn��^1 ����Qm�׳���19R�D���m��q���*��e�v�d5�&D��=�{�E�n�R�E5�F�/���ر�-`L��|��[��r1��2y	/��WAf{f0�(y
�UK��8y�ѵ��ی�N�����>*BiBQ�_�?a&��x�e�˜�n�32���Z���� ���3�͒'®��/��,��PL����fB��#�d)OAQar����\RVl9=���:�'ˇh��c�l�\UC�gm0���@�=0$$����_gbG}$TcM��4�Q��K2���zu�@T1�l�7��,:R�u��q�w�k�^l��Bs"[��q�iP�B�~?��g叮�G(���^e؃��/p�4�J0�t�%=%v�"Y�h:acc�WMm���>�7�C�i��"��[ְ�t��f����`�.�+Bcމ#���?�Dlv�������K!��,JW�2!P����Տ�]��X��a�� 5?l8E�H�ٞqu�7��4@�^2�Ty�S-����( /ԓ}R�0�V�CPS�Қ}��jZ�0d��ߤ0�j8��Y?���E}.��w�$6�Vw��	\D(�.z39i�R���� �s���9�ل۱��j���T���P�	�T�`
����y�Z#�>�+g�vj�2�|��3�s �Y���6�s���$����̇Q�>��A
�V���R"n��Ǭj��h{��y�Ag�f�s2m�w���Ol��1v�%2�����~VA"��X"������R��Fd��Ƕ�1��j{ �������Up�[��=����j�)JH�^rn�Z�_�'P��Z=��ae��
�9ΈA�Q�7$��A�	�7�&��k㗩l�Mm�~���
��H��zT[u<����ǣ�����nS��_�Z���NO�s�,p޻!��i�v�!_,RPJi�2<�=�3��wMp��	�c��$/6F�P�3�k�ո*k߲�co�YK��qU5_�������˸�0���@P70e���d��)e�7����?P͑��@(�h�����:��{p�M����pH8�1�i8������y�������P�3����` �Q)��d�&�����1���nv������y�H�<��\I������ɓy�� ��#��N�z�
��b��������n�,���W�W�]iGL�3��6e�j�cڧ�:�$��T�Ee?�G�u�<�c/$r���٩+R�Q�e�f\EZJ��ߊX�ot����P���D`���SZ�⻍X�D4Z����w��E�P�����^MD#m�/�%��C& $^�F,�`�!g�is�*w�����䋞�Z��ψ�9͌Q�z+�$�X~~=g�ŋZ4ѯ%~/7H4��8���֨�>�Xe�� T�&�s�k9�˳!7��~��|+/�~(��C=k/k,=Ek'+j��F穐�9�����c0�K�5�jq֢�U����t�ί�f��պҙ�_nt��Q�G�HGk���'!���wŇ������02��>"7cg�-[�S+�{V�"���'���z��z�ʋ+�"F�R��p��l�@���@���S���$-S�O��"�yX�����ޠ=��H2�V6\M�V��uɬiy��
,Zg�_��h�K�ƭh;G���KjN$ɦv,�o�l���1�zypZL�C�Ƶ��u��٤�kx��N\m���9��^滋�����u��^��p>�����y��-�Ӏo��_�vN��aM[�7���}�<}5�b=P�sd��c��~F���J:Eѩ����m��r"�D#�$ bmt%�Uz�ߡ7p��%GeB���.t=`��g���r�܄��Liͮaa
�uZ^�Da�?��`�0��� %*7����(��L1?N%n,J�]��D�"�4� Z�ρ2g ���%:Қ8�1��f��������nQ��A4��:����˴c�|O�+�gF���넠�N�TL�����J_�F0�N4q?2`�I��])#h:t��i�ڸ؄���#�l�٩ ����z�k���`T�dZ��3���`���O̽��V�@��o��0�2��oX�#��%��P��cH�-5�#�Z�#䲀A �ֲ��[����d��Ɓ�D�"����u�M����E��y�U�Hy��`��߉�4��L�M��~�RZ��m��0���踨��8Ye�����W�v,R���Z�g�Ʃ�uJ��~&z�0˲/�Ǐ��|�^��]���?3�T�7��l���c21(���ĸ���z��HU�쒆I�"��VFu�9�m���I����=�|o{�H*#�lL-���xKf>2���O/ݜ#��T�ԙ��5)�%C ����1�-`�FN=|��u@��p�Fp$������9�%�ˌax^y�r��[��gB+�� �W����h�Sp��XB�puO�����֨`�b�*�����(}=�MwG������[v���FH���6��"oR�Tn����Tn9(���<�!p�eӓ��O�<��(���߻��E�r���`�r����Z!!ɩa����X�<�����Ă��MM s�����"A¹����u�٧\e��xk�A��(CD�$��̶+��̒��Lڃ���ʄ��/Ǚ��8����>��es�e��vc��-Z9ґ�E�??Tv�!�<����L�=`�Mʽ��Iݓ�}+5P!s�E�[���{�Gg�(w�ou�$���C��(��ܲ���^���N�P�+{f�*��p�����-�6���	9->囁���>A�{�oY��+v	��L�/�2ױ��tC��/���06�K'@���AI������OO/qY�<s�8U��Gt+��͇b�D���\�˃������_�5$amX&�R��<Vs����c[Ă���O��Lz�b��/M��3��h���sC�^����(��l"��M���
�z��_[�l�T�:���8�U+����>�H�^r�_���$,����hf��V���O��tY�<�g�/��v�Ё~�J�~9�E&���iʡ�a��p��eӤ��c�AҞQ�a�k���\wA��HY�S���6������p��4c��}e���^V,�Q��m8s��V0���p(���\��] �dL;Y���@Λe�m&K�M�,�RȐ��̽�{�!ܤS�X�N�	
��x� �P�PS�j���w�j��(;�Y:p����l��
V�*!�����񗙪��0E�w�ݱX�$���dJ�;�)��qR�n���T;A~j:W���-��>�� m%,��\ms�DiT
�/�j��f=`��h�#/�W	��A�K7�w�%��������X�1��%���`*/��~f3b阹���W`��`�ۣYd���Nl�������f�/'c����X+��.��6��ZV?(�iP%��D��3��t����+}���RO|D�B��a���V�`�k��E��o:FL�E0�ŵ��:v��v���O��.)?�Ც�����P�P3� �"��r� ��i\t��A�����v=��U���Y���
DW۝\υtYi�K����H +O���sC-)����>�Q��U\�����o�Q'K���!�B���$O�4�1E(@P��/{
�(��c|�,"#;��䎪?��W���BAr�-'�G�|L�p7#��D��j��ʩ
 �T�J���<aſ�r���b�m��F
{��l��s�����t�ao&q��s�q'���ͽl��=������S"b.�ۑG����֚${q��C���l����;-s(a�^�� ����q�Tʾzf�Dpl�,³"|.�5���҉B4��j�� �?3�2ڼ�*\/��Ϻ��OP��EF���ߦ�0��7�Np=>����G�y�r��d����o��[��i$��dG�+_3�����B=��y&>5UВ��#�-����ˍ��΀n�����)&g+���%�D�	<�>`>��$��6\(�W~;"fC,)�W2��TV� ��
4��u5��eMW ��q<�,��EW�+w��| �R�eLU
"�~�r���o�y�\Ҝ��늎m�Wժ�7�vjC5X 8���Z%L#��%X&Hv�A9e&5f�ޯX��i]��L��냟F�%�m�$�k@f	�	�=���q��r�AB$|�r��<x�T��� �z���f���q�wk�f�jw:��ɘ�&�����6�*�?��O�F(��e�*��h̟fϦ��}����KuQ���AQ��8�q�^~c���u� [��W[�k��Y�Q�@�+��4B���!:M�~����f���ad�2�}{��!�+��~]��(���o�^@u����#%#���ɰ��3%�2�����a �6���7X���t�7�$ķ��"�]���T/*�ȁ�.�d�K����_�9�v)���h��	VFl�-��� }ءŉ�PVU��@j��
K@�C���bs"��);u&�)֯����ٷ�,P��]�t��%��V������ud�ː� f���y�g��7LYQ6��um��
�'�4���m�� ,��Pҕqh���a��"��{��K�E�%IRR�"/�@�۾0��:/fʫQ����{%3��d��M��ͪɝ8���c�-�F�ߢN8q[����p�g�@�b��>�|cte~����,�ޚ�:�mF�+���+F
�)Z�i1���" �[ec�'�m��m�ۧ������%ȨW�Qdu�m6x$�{~[�n`f8�um�@]�Єm} ��L��)c�#yѼ\ k���Sh+�}�%���+.g��pZ���+:'�0+}�NѢ�o�t�	RK��{�|��^���o8����H(~E�����G��7�,�#$.nU��m��-yl��H/A�I���Q$���H��"�y$��V����P�pq��rHe/W��F���``vå�f�j=���}-�cP�!@�3��P= ����8<�/+���(��d�P�j>e:�)�A��C�����_��#�B�*&Ѭ_�t-J��ԭ��qc�D/R�G���D���_��Yo�4�O�x��P�O.!aA��މŢ��pn��ا����SK��U�Xݵ�_+�D�A5w�{��R+��lg daŕK�]�bu�w�?j:!�5d�6;L700
\��ԓS�44�H�ɱ���+�{:��O.�f����~�rL��!XzIխX���M'B�&rn��?��8���6g������h�J��!��քm9��(QAO��Y?Э�t�=��ݺ����6���z��
������*HYdA	�C�~v�$�ihq�J߹��^K;?^��[��}59o�%mi=�Vқ�ܨ��0�e=$���u�*����-~���MK3�㞻��5/�9��d��J���_6ع�@>��0�kV��l�a�����w��'��Vd��]��"�4��7 �ƈ��͗;0O�%*�0Ձ�b���+��!�"ݍ+�X�����][ghZ'�
��z��+%7D*�u����aK������b&���H��JZk��V�[����h�47�'=+�r�����0[�/&�?�I�`S]V\����b�ED>���,/|ao:���dqp��T�I۶C7��I�I=��>�Ձ��<@x�fл��vWnK��?�o]H	w��x�w���u����k�����1pc�}�h�]r�t�1-L���NRr�����PE�E;�QGn�(��mA�.��x��He_��e��@wX*��� ��0J)3�"��~�͊l�bj�\��XO|P1��Y���:�F�꺊�#k���Hn�t.����Rb� �k@��<~G�(����R�d��U�@`mJu9��_�\��0�^�f"�����a�FK����6���3���m.���~3�<O������^�jl�!�۱��8����҂u�i6�痐s�ۯ��
�d�
�J�En"S(��e�H�5�qAˇ=6�N�/չ��)������5Ia(n������x���E��A���;�z�U5WB��bgM_'��G���5�3�siL}���S�FX=5N�����V+!�r��ơ}#�W���k8c�7��\Z6m9�殜� R���MT&���/�I��W�%��>kI�1���oo���ϑ���.Nb���Xg!x�շ���c��ҵL ��c�D5�E�ו��/jiWNZ:����`�Eaڦ|a+������ *�%��D��r'���ܼ��"blװ%����-Y��7�>���&[��7_:���y�1�>$h������A�
�m���1W���Q%NJ���)M�Ѫk�s�� ,��`��D��k���9-��7f��RmT�T&b�)6��߮\�\Ȁ$ҠP�Z'
|i���T���K�9�Q�H��bFq���]�K!���j&��b^�傉�~�߾>�׹�e��U!��0��N�C�u�x����{���ԫ1Z�q���t�{2B1=� Ƀ�bv*�O�M��+��bξ"���H��B(�:�=UWI�I�+��{�8n^z�1G_�F{z��mYG�
�q0_�M��	���"8���3�E�6w�tw��V��\������(gd=ߌ�	��c�@���P>{�l��^cb��j`X����1X2[�H��2Pv� O��AL��<�U��r�o�^,*z�YDx
1��.K�%PK0�*�N��5fԦ���7�$X��L�-V��q���K�r����ȵ]ͭ3�֘�h5�.%��?�4ô7j���}6f
 � �̿8�XO�$�f��I�;�&�B����W�����,�O銻��Y.�K��prvmdc�-���(	��;�R5^覔*o��O|�TY�������t)crÂ��8��y-����m{�cɥv�]7���W�{��n�g��N:
���9DBr]{�<k�~��J�9��6�'R�J<���Q��K%�q ��၅:6?�ي��}H�f�-�Bu4�7����Y��5�����vO�~n|���`@�b̲�Jm�a:ҭ@	�ե�������[�\��V.����Ə=��T�`c������+������d�6�B���1��V�a�lY�7�ɒ}OL!��v�0Jt�NPT�B�'�m�(Sd�k�Xd��e�K����0�ә�a����Oɓ���/��uM�nҗ�5RY��-3$\��]R�N��h��M<�io�{�.����R��Ѣ;7jR�����y�dp���w�'��67�`T�iVTI"�����X;s���`�!o�4�Mû��Q�P��Θ�
2kk	�[���}ȟј�#��v�= ��M�.Ǚ 	�7�|u$(�/���4(, �����C�����w-�<�]�9o�9�t�3����2�1/����{'��7�hQb���e��+��Ӧh�( ��uΐ�/��6��(֤��n����rV�BE�ʽRC�\s��4�q)�E�΢Hz��J׻�ǿ��W�,D�[�������ĵ�+Y8��9��')�����\Fv���rp�n�㈋�!�e�f��0IRy��!�nM�[`�7����$��3�?������+�J0X"a7���h3*��O٬ݞt��L�f�8�>g�������*�-��@� _]8��R��z&�:2��BAsơ`���<��~�v}N*.��5����G�QcUqU����.��'e���.J$�캇ij�-��������N2N��)$��Z�$Xs U�lx���|F20�{������#v��'����_���M����v�ˌmM=:��1��(�L�Q�t�]K�%�,9����x�(��˷�箔�K��=Y+��f0���~O�*��i����x\$�8�=&�o@�p�2&�C�_�)^��-�x�yxˍ�����B;�PTmz�>��:�r�_.�|e�����A��8��{��#*���nT��*�
�[ed�D6�p��`)�~{����w�x�C�찖d���<�u� }k-�u/�]3��%��tK��ڝ:�}d�U0���w�>ԟ��������,8_�3�
�����z���kECSeX�3�x2׉ٻ�a$9p0�'p�y��u��e	h�\$k����]���\������D�Pb÷H]�?`�6��9T�
o6_\���/k!�R�W������6ս�R�J��ݜM���la��ݔ:��A�,���/k�[�IH��)XL��^)�_8�gq�)�J���.݅g'��*?�ӷ�&4=��a�������iG ����H���.���r�zo�Tci�E7BOE�����}��e��ϯ����+�n�d���#k�ѿC�\�\��E�^����SN)�H�\�
��OT=[�B�p��+���a+~��C�NGUk�#
�PF��|�/Ǒ�>H�O����W��lW�cnpwt~�n5��r����m%Np� s���?�#P�%��(ht�D=�����Q�Hja ÓTuo��C�|��@!#� �4�H�G*
ig��+������w׹�ĸ�WE�=�j��|���"
q{�������J��h��/�����+0�`�덯\�xIV��b�2���l�o	�Q����u
?����J-HOk�+t�b�j�ߋ��Y��S�����4�_Ԑ΁w����<M�c���HP����|I\�%��A����(�{�ٝ�{�1W�u�*c����}�x�m��%�_�H�T�+��!��\v��6@�9XOr�	��;#�8Ib!�W�ݖVFH���)#X�kT���Oz�E�6��5�N�R�x�Bc�sj�c����\J�"�1�u����Vr��-毒��,G��7��^�8o٨���/�PR�e�����.!���r;��k]O_>/lb.M� Z�Rɑgn��Me(��V�3�{z��n�UM�@)�7z��}8-������t���
��5t�����$��=����P7l����9���{�pP6p(�����)��׈��c�V���w&���豹ꃥ3�R��OX�Bڟm|�~�����`�(�c�e���;I�mk2�/��Ğ���Jؕ��Lo���5�[B�p6X�!Ėb��T��*�Rlj.�*�TXP	��\/�ԘU
�W�U�����\�mXU�d?FG=S�ta�Bm�À����?>|����IP�}'}�' d ^5N�*��͛é(�<ޯSX�ιh�x�#k�FR�sd�Ь3M����`Oj͑\��u�4����H������������Jn�o
�{� ����I-q*f���n'��w^�*�T�&��n�j�LJ����qrX�z��>��7#p
�i������'l��d��N�p��M�}�V����}%Z�N��x�6��>��w�ڽ��B�{��^7Ɯ�O��b�b6�����w3�w����J�����I��=Ŷr��+MO����c�6X%i
�wAH���L!�3Y�峊��xl��c�}_F�5���5��dwh��QS_�>��w�|1��x�Oc�]�E<{�_�����üO�	�����:�}��hC�c�~�2H�[�$��k�|���5M��"���ͷm�ߩ�9��詶���)i��}�Nl���{�K+�NH��F�Ệ��͒����{I�����i|������Y���a{�~������iH�B�o�d���X?�vm?�@�M!���/^��9��x=��QE����B[�y�Q��hR�_�� �X������ne���9���|�M�N��X�ae))g�wVj�`S-�q��t谛,S�bD̦�*�2ӿUA2��Qpj�ݶ�X��<�5|E�1�:��6Q���8���Z��G4��)ȧ�eN�Kh�/U�Ǆf�Um���7����2� Gd�H*=}�?�{��,�zI�(�!o�t66f�y*���#`�%2��>��Q�a���!�(뻬N�x&�4a󶀜;�e0\��OI�Yp��{�e_���TU̦(݁��P~,MN�H�0�f�#)��xY�E{������v&}g�����8� ��K	�q�]#t:��)�e�x���8m.���u�l�b�m���������cn>x��A	� <Vϲ�uqs��!ϱK7��DH�B����z��.z�������gj����w2���S�%��h@�����^�}�Ĳ��&`hb��	��꽠�@bg QOSW6�8�e�-�4�ɘuLxy�ƓA��o��aJ�b�L	c0ɼ�+?#���ހ 4A�f��w~j�F\/R7E�>���;�W�߮�x�1m����PJCC&����?f�&Ԁr�˔0(�&��s.����~�Y]��|�#N$���+�^#�D��G][��v�!Ez'����,C��%�,�[p�Nob!#���.��������'��2�ڿ��1xo�|�j��Y�ǡzB%ģ�5җ����:m �zZ��LҨ�]�6P<�����C+a=�ãb�p��`'<E����fe�0x�xGE�T�����J�U�?�~�2P|
R��$M�&JTV7k���6�F��tb�A[\ajT�x��V�2��]+��j-#/�5�M{aمRV���	D N/JZG5���hk��Mα �l�~o�C�ay[�,I/c@��Q���.�=�(�5�-�n� ��H�_�u�<�T��������.���&̽;=��f3�y֤��%��TRP�>p�����&a��	� 5�c��b��淥W��{´ǸeA�b_f$ZC!k�����gKN2�2�N{��Z/��gƔ9��@�ȭ&(��iiM')^��sו�=�(���k��H�i2���K~���M������qҡ/��ꠣ�USv2����c�	��2��˖�`,ދ��G��O��m����Xo��g�#���w�XJH�|Ls!�=R|x��}"E�q;����X'SP!��Ͷ��H!H��;�h���1�V�ErY�ԏ��T����"��-;,p3���W����p����<Hp�iHSk��2٠k��TD&-/�
�08EK�F�E��C�����=�l`e����H�cn�M}5���/Щ����T'?�G&YȘ�S.GY9)}����`%�z�z�3^Q�t��r�::+��`sċ�;QC����g1���	i����M�Ow���hS�`ǩ����'�Փ�ȳ��X�1%�5�����u��zg^%>��a"�w�Ii�U��/����SҺ�5����j6��3�)(� 6��Ҡ���E�M��~�Ƈ�(0�2m[z]��}
����c���zҦ`\���>�v;�i��j��z�$�{16�d��.����a�N��j{�"F5n%�}e���k>�v�B��`E�@v �tgvٛ{@�3=�i2/�p;��ܣ-�?��2���i�y��\��G�R)�)#}|G���O��!4�Lɮ�U��"�4���R���;�	Kl+r������������~D��k����ž���Ԧ���߫[���Ѫz� ,S�(�rW��"�d-	�`{ө=�i�#Z��|ɽx�(�R�l��0�-O��!x(�g�͜���e�/���5#�G'�ui���۞d{�gy�5����k$�V��T�z\Ravq!1�����p���|%55��|���m�ز���)*~. �̚�g�O��B�U@;8�IY��$V�/~*��7�s�,�e�� g!_�v|� �iٞ׶x�+}�2�&ɻ�}��=]{��*{ȓ��J���v��]a�-m��V?նP��_��Lw�u�R^����He!o�@���{Eitc7-4�!�'m%Y���]�P�I���χ�Dә:�u�X^~��?�"�Z�̥����`$\�@_��&Fأf�Ѫ/�>���"g�r&�@��Ԟ��Q~�^�$��H9wͮ1Iܑ~Q�p���;$���`ݓm�RAPf���X��\=}�M���z��q�@jS0@8`ˆ����aI��p3W��9�/g�O柺j/�����=Bˍ�Y�#�-���4�Z�'|��.�z8ū#�ĿP;&(�0ƨ��Y��de��� ���ez�=��`����e�HT\;�����ۨ/ժ����">+�wt�[ D}P��^��D#Wd��{��n�.�ft�Z�'��p�C�d��d�+ر1���>'��8���T����fHy~��9�Ë!|�b��d���+���9(�f�|�j�[��E��~6Tm�o�	-|ⷲ�?V��(�5���V�Nu�$��c>_1z�I#'D�M0�>�c��i,D�����ٳ� ��]غZ�����.o��=�iuˡ�%�J6���aʫ���){�n���B-X��z<�-󃗱b��;PJ�F-�L������o���Y���J,,�n<��β Kt=X�S<�>���Ś�fQ�J��3���~���*7��A��V�&$x�:�b��.dLFw񮾋���� ��)���d�8yU����"e����n�.�bxg8���;�����&U�Z�ʿbBp~��1�JV8:��q��7�L��R��z���팈�YJ�m���p,sz��e]4)H<]�ɣ�S��k!��]�|1����}��܈���[�S��@�� 
���4��(��i�돓*}!<�x��Ua�H��쑶cW嬻F��4������0������ݶ��P�!,R�F�-|�( Ġ'%�!��[�X����+���#I	��w���&�k�ӥ�lS,AC�~�N�mNM�ou�P%7�YX�����ph^�p�bu����T�"-�����>��^ݮ�{�8d�����}��8�Qʇ�L��W7'�N����9E�E���g�bdS?lt����T�"*#U�4��J�>�bIhK�AA>��wj�@��m@\I$���O/˖�Xwc�hNt�w�ygR�	��m!B�}�˩�$�.:މ{}�!k���?�ѡ��ʻl�K_`�s���A�Q�1���h���m2U�"US��x��E��o�����5�S�m_1s2Ŷ�  ���˭�m��j��`�����(�ƅ�˦�L%��<��m��Ga�{R��{gΊ
�c'�iW)?�.�AD&���@!š�/^l�z=z��V��wS;�� b΁�y]�����ʕ`K�����톜��7�+&��YV�y+$J��VR�����lBf,�����r����ve�Z�PW'�b���D("��U��t���?�u��o�/[F9�|��
ڸ��zR�l�Q����/(w@���(��|�v��6[[9T�-���������1�t�x���:�-2�EJb�rr�!t�򎋱y^��j��=�vݸ�,����fٶ�����'
,4|���	o^f�P�U˂��F9��)ps��&��lC	VQXWE�&C⏻r��PO~�6��kj�f��6����
�v��MH�	��P��+�JY�1W��ܜ�xA��7�n�k���B�D���$U�5/�]�����U(<>�8�>댵�c$���V� ���EM8�1
�8Jrx[�(��7�����}�f�[�(�ߢϒ������)eK%XdM��4��J��X���=�OAY���F����~d�0!�'/:5�����0�z�tOUc̃G�b�3��\���2s��,6T@���P-,מ��x2��5xc��S�fdb�ʡ�S6��+`���Q�E�{L.��t_/�t�{��I��=�����6�Q�#�w�z��;T��r�����us�ҍ�)&[��xӴv	�>N�+�d��CàJ,�&u;@Ͱag�\mt{�$HWȼ
���EM~�\�9����2>�p���8zt�g�!v���T#d'lLR
��3G`�ʌ���HJ3��Lx�ƌW�T!�S�XɞR�~��b��N����^�hƿ�}�P�����霪j��|�m C&���X089�����JۦiJL��������j:�)	��K>�S9f�HH�<f�z��N����=YQ�G�~W��Zi��E�Z3l�D��X����	���Ϩ-�6�uH�_6��9yc���6��R����c���,��� ���qg<O_�J��? ����	Y۫�R
x\��3��*��;�P�6��Y�HݻX4�U��h��C���)�?� 貶��af���Giw, ea��Th��ݾ'C	����%��2R9��C�nW�h�2y�ǜ]�����c����Y�w�b�T4]�q9X��-���2[���;���g��Z���q�ĆIk�v3P���ܷ�Ɓ�S��;\�ӯX��*3ړt�~�5��'GU�j�"ks�>�ƕ�rz
9Uǉ:b�A�B�U��34�y�<
����bq0�w`�>�����W�9A�����*�c%����A]Ӛ]��9���u�(�ߊ��d��F�ؠ��ڏ2���م��u�D������ٔ���;�3��pm��\=B[�ƀ^�� ޮ'r�W�yuk�˚6q��lfÛD2!E��:����!��V<�V��Sqk.a�\o��# �T�w�Tr�CV�'��r!�/5���\��Ȑ�����,B%z0c�ofޟ�8x���I����5��<ڴ����������ѹlx͋�'�����(݁P��,���p���!a��[��`�1��Ke&��Lv�b��)� ��=�]�e,�{�� �"*))�T�'���|bZ�9��nzl�	ێ%b���Y�6�Y���$P����.nP�@��6�*�2�y�2��b��%�q�1������<(1��|鑾�gۆ+r^ç��3�����I˔����-�&	�bT�feU��2s,��O�,_ �x�X��h]o���&1���;� ����~i֭�m��o
Ι'�Nj���ki!�)Q��u�����Xr�A`��xjp�����&�fud:Ĺ�m����٠�FQ
���8�'��G��g�=��8�@D5]��Yl����0��*	Ws�dY��>���|�9�F��l��aat�d������9�ԚL��n�렏dU]&;!?�8�e=Y�63�vD���B?��ewVP�	�Ҥ����h6H
R��U�h'Lg���͢3,��)�g��{����-������u���.�7��?��x�\5SY��N�M�t��UZ'�Oxy�����r_'5�p���O@���ZJ-t��,;R��4V.|F�U���ѿ]OE"oe�C51����?�Q7����^)$ɬ�5��Bz즸��R#��c��	O��p�4�)�����쑘ٙ�(dWR ��	/����W�����ɩ�ҙ��\E�ڜ�&A>���8�&�]�H�N�;��*���G�jx�:(�-��ն�����+Ͽ�fw�-�`*Z]��$���M�鮊2�N������Uڴ�[����Z�e�]
�,r�/��r\�#��Ϛ�n�`�q�a1�%"�n �x +wӾ��֥�|�;��r��������8/L��c�p���>��F��d��y���)K8Ϳb�+�s$�%|m�<���eǋ;�*Q��m�b�!玦��0#@;�l)2[���춼�n�ɜvTy��:�� �9�cTh�����}�}[���R���]+Ӡg�9�q��>T��e�F�bȟW(ʇ��t<%��c@��A���X`Ŝ��4q����Z�mw��d��U�8���I.P�߽�`�ܴ-�7�S�9�ϱ���P`b8�����F+UA��ҿ��@#\�Ɵ�
����2\�#����C$��N�s��=�����g��f�R�g�_�nP�Ӏ��abZz��3T]N]xe�	�h3v�Ȓ��	����м0Ҹ��Z �,��ׄ��_�0d=j�����,f<n��S�;ĝ�@�o�}����RY��ѳ=�^�s��i_!$@���A'~����/Q��0�V�� ��D�1N�My^��y��[n�T�}�����W_�}}���V�[OHj"TX�g�έ��Z12Q�W�R�D�Q�ߕ<y=������y��������S������g���PBlm��+�g�+h�;���w�y�;E���#��66���<O��I����.0,OC�(�;f�4��E,�Q ��M*�� H���|��8�딦|M
�o?&�%�I�0�@q�n.�����=E8;aa��n���';:�Ҝ/�Ʌ���r��������Kf�QziDFJ�`@(��t������)o���'#����#U?��o��-��w����餝�� �&7�#���Y? �-���,�����K������4>�$^�e�X ^�t�ϟ&�b��Ҝ�'�۠,�;���Ƹ�x�
"�S)F�|��;dB���+�䆢kaI����_.��*��_����da��ɣ�;0�K���W)�l->��tfˠ<�w��x� o�� |P����p%dz-KO��:{[Ye0g/;:֡q��}�������͙��s-}O�o�ԞSn^.�� ���;�{����������/��5]�: ��Ӡ~�^�ߤ�d�V�<_j�O$٦�ZƲj�T�!���sX����&&���e�:�1�fS9��n�M��2��Q�;�����/+��h�]�W�"����G��ʨ9��x�l�k5܍���Q�_*��O�SC/ �Hv�_�?�������T���DHF�面v�$��� 0涥v�2M�s�_��‰�u�H����~P�A��جb��~����*�Vlf����˰���sL��2��{�E��YUW*ˇ�'B<_�=u�����<7���~���
�k�&nNp+���<��J�)�����-=����P�G[2�r��݆Y��QR$��ڪ|>�_ݜv�8g�|g1�8*�wr(�Z�	��)ջ�ל*�������n��d_dK2$X���?����d��!ꦃS�qn�:L>�3�$��6q��Ky-ِkg��
Ʀ��j�_/�K�m�bQ��BR&%σ�j�$3��%-��V��XK�B��J+`K��i�%\'�Κ�����:��c���/��c��氇���߄�rUn�y=K�<g��:�XP[�/�oΎ���F܃�V�'���"��eL�Q��QQ����H�+��o=��')I�ySL�dEEĜ��G�ES$�=RHq��i�p�E>���⫂46_��QT�%�c��j�1�2nf!w�a+��)��.N�G�b�rՏ�|yK+��a��>H��"�n�L	igM�KВ�҅\�譾ju�d��gh˛9)V�u�����H�����a��GM�NA0f�"������2�$�,����]�"sWp�$ϵ�	�E��q�k��F�h��lc���|�-��5��fo�NQ`�Y��`L�n���/�Rs�[�;�R�;�!���sv����H�w��1]c�Zyc��#"���P���jE{j\q�$N������]ջ�̈́�}��IQ;�[�ZA#T���}԰z�js���f����ę�n|�\����}�_ӗL��K�.d-AnG/ǥH�)g7�t�J�d
h��6Q���(`_�+�h-� �׸;�/K�8�r[� �	(e��<��2�׺�4�B_O�V��4����9o�m�+-v>��⸋=�IL����h�t���8���b��N��T�sJ.��P=����ʴ�+��`��h3�Iޞ '�����޾�F�B bnj�W�+�K9��P���ǀJ�R(�W���|��3nrr�*�~�ơ�Q���'I_8;��uqG������/J� �B1�f�S)��ja߰8�Bw�^V�\% �Ċz����EkD<T��X��]S�|ؘ��j`_r��a�$��_�����農eȱ]��+�7�����m���+����e֒<��W�L[������C�X_uS)w���[����n���M�dF�-���	𸬦}U�Y���18� g�D+����-�[X�2E�.�|�0��V�v��mb��C��b^�Λgb�q����/�����E�}m�EqHAd��r�����,�I+{w燳�=�[��b��7�aߟ.q��u����	���u4����]z����j"� ��Vʩ,�I�c�R��ܲ�"���M��+7y�)^�Ԫ���(R`6�wm�i����+vX��? ]�w±��PѢ��U�Ľh�� �I��3X�7��4���Omg7�Bl�)�d����&rվ>�#Ư�A5;����pX�v6ξ� ���oJ|i���!x++��\�q��5�À�s��'�/a�i[`�+���V($�Q��,9Xq?���1܊.�wncl����
�;ar�%�L,u/ ��1`��P�S�W.KV���e>c!9U���t��s��]�WDC��A�H��?v�쏀������ƀ8�.J�i�1<�[\GC���M n��Z���w���O �6}6*����] ϗ�mF��:n�\��/�Ӯ�[5%o�wּ}V�/�Po���@ٌ��8�+@�oM�^/��L����ل$Ə��3V�i>�չ��KT��<��!G��Oh;ژ��-L�OhK��	G���,���J\�	&��g-Y�U�ۆɕ�w�줋o������J�f�ɇb�������,�L������/V��zt�rr����X%�=e�Z��3P0"c����/q���-)�jq�c��S�s6���>?�H2;��_�k]�ҭ|�����_x&�Y42U/����I�{�O~��N�1B�Kk��X�_�,<blV�K|�O�g}?�|��GH�s
���И�'����:�қ8��Ǘ���R0���f�����5` �\N&����l�;{Ϭ��̸�m7��ٜͯ�=��"��C�6;��-���q�A��4�!>CNFoe}����$}�$ړQJ�qSIqۼ��T����<�T���} C.�2�&�ڌ1!Z}=����i9zTZ��E.��i�������&QI�������
�@=���񳦶-�s�A��S%��鏢�/c��Ǟ;����{�5��-6��:��>���Pޜ�Z}Ъز�땯���+�ˮ��s  ���4��F_�8^ٿ�kJ�/0Dr �ܰ��V�Ր���B��z��h�"R�yO�����0xZ�]�:�5�=��Se�Is��-/> �3'�{�N=EU�f��8�JzN��������="�[v�4۔�J�5Ak�
�雛�@�3ǿ�3�2��H��Z5�ɨ�h s��}P���1v�� K@�q!��f���&h�9�?���(�ս"�c! iQvX[���y�`�5�O44Zx1lv<�Oeg�%ӱA�JG�����+���ޔ�6&���1=|������Qwٍ��L��*}���S[U�����n`ܲ�wc��ޗX��l8�}sD�2M[��e����n�]�OmʒvS�?LL�f8���瘛�Lc��n��/Z�'G���*���!�i��/ pD�22q9��������	�7 �9G4����.KS�)�wǰ�����C�����D���жu �J�6�85�q<��8��a���B�������m��Ψѓ�ZT�u�m�9_I�#Xǵq��9�<��g\ 4U��/^��<����b��Y ����l�����7|�̂���Ǝ�4��i�?��x�V�mTA�E�Q�/ٖ9
��t��
��{�p����n�W)�Q�4Ƚi�<�*kf��qR�<����C�΢8�1=0�^�7(���Gʚ���FҘeR��2L�;"�~vӟ��ux!흡�����\�"Na�?��`*t�%z���w��=�5�0��; , �H��m���Y�8��lIb3�����DT���L�!>��Wf��ǘj�V}������w�ke�D���)���������3����NS��O���p�_Ƅ�O%z	��O�������C�2�U�,&�ā Թ�bce&e�r̀��<Q�YD��Jf���Ƕ�9��&M
"�)��B��I4�l������ţ�4Lfe�ם�]un���;"2�;�*�e��}b7=���o�Xv}��ㄴ/�t|ש�(��i���S;�����@�$)ڊ��+d[����m]�uf�k*$�_�RG%��k�u������SS%N��
Y�g����F ���6���?�:���m��Sr+�m��q�%ěm܁��D�ܸ��r�nc�w��c��o�_�,�6�Ƶ�$ s��}��y��\l)��~3{���|��.r=�8��g�����,O�''��ce���.RhK&�[��7��)7�re��v����uzR�wK9�܏��h5E�Ľ�E���n��"��7��_�LD�#1�vq?~2�h7��}���h��"��?��yFveCڎ�ྡZh���rx�J��^��_k�g]'�i�	��G�}���Pv%-�MS �	��M>[S����ݒk�%k���J�V��������Zy%��fs�����h��i� �9{ �O�!:ebX{�~���ī�w�#��JC�>QjT�s3�D�B��x"ٷɿ�Q9vJC�va�G9�N!��)�Zk?�^�d����f5�`�6�cή�~��p��jzYa�8K$i�=R;�$L��)i�f�L�:�,�� a�Z.H������W�7�n6�ʈg��+w��2��ڲ�%�w��%ER�~aԬ��M�.@�)�����!��d78�~Q��y|��E��yC�9�nkw�y8	��z�csdgq��3���-,��g0��ZtA^��������e�9�	�h��#D�%:Z�p��}�2x1�M��+�I�c��b2����n?�m ������oW�+���j>�
2����W�A�G��ש�/�N�������wS?�"�c�V~_)d��-,��h�@[�t�7B7�V����_����qwGr��c-���E�L��I�Oz�=���w�_�d���y�jBc��S�&Om��:7�S����K�	���!A�:��gg�
r�[���B�wX,�ިL2Ґ��*�e���SCpCM�Rt�,5'V�����v�Y�.$x� }i��c*�'��H���݆���V��LvR?po�vjڦ1����?۠�9|J�bE:�4:u��ߺ��@���B�$d�q�U�qg�?�\��g1g���Q2ѐZP f�Ͳ_��,�p��
�U�M�[���ĩw��ޮ�M�m����Q���V���S�Q�k��Iׅ3����2<#yr��ԓ��ɞ���~�-�;I a֦���G_���Of�W/<��i[��"f�_;�m���(�N����m�+%>�͞횁.���$�^h��'��e�A�D"�_��.fY�}9�1��zSi�b�n�>d���Ԙ���S����aN5�؝*̦��v ���i��t�@C(f�����k5�|d��v}a,"�S����+�	���7ۆ������'���X B�Hj�"�R�<
���b����;7B�~�~�ɞ� .#i(h��}*���rw"�p̜����,�W״XC3�	d�l��Es\�4<]��	b�N��-�t'	�E�K,EF<F�Q�2��Ƞ���f��HI��UF��iͻ7���V���'�	�+#Z�7س��ZG��j`��e���ѠxT�+c[�9�1�UH�gѮ�̎��S�I�O�#�@[���|Z1E퉧���T�Ćv�R�~-L�p4�"�.6�}��VC#�/��{kTw�;����,[
,۽��&�L�o���:�*���B_=z��q�*h����]�_\ ����9���2>��u���0��ű|�S+HԷM89=���U�!��&�L)\�j	�F��!WK'\Ja���p����UCI?J�x������ 9����I��ZD���k���E�����'ܸ'��A�E\6/��d���8_�c��~�yf�� ������48GO��Kk��UWy�]j��|��0|n�4�y�sF#�W�M� �Щ��	��4
91�T Psn���GZ�!G�TrR�X�9�� ��R�v���3����v6�r�,��sg+�LC���82�bc��LR�X'+�i���(���A��]r/�7���Z�`{"u\�������s撦�Ԕޓ��� ��#.��zl_�B�r~}�U:a? �z�_�?���+���7��zf���ӕ�hӋ<p鹋��:�i9���jՑ�o�}R<�,P��),'FG� 2�ϱ
ie�)ƹҝú٥|��l,�\�!�#�n�9 ����3ڄ��ms�R�	F�!�	���=Z�6��@o�^GD��<w��IN����wso�!�;����T�_^���y�x����x�t6����T�
_%r�A��Qp����]�;ڇe����eg+.mުw�z��v�V �	mu��� c��e���v�Vh>[�����.M����Ĺ�&a���s��)G6-[PdiV�6b�j����l����Q � ���@���>������5h���eu/N4��&^Q�&�����ds,?�5dGU�戂�S���.�H�HA�t?d7(��J6��S���C��(��T�7���$�z�� ��/��y�N�?���������<���r�GO	��i�[f6�FtP�\�17��,<Ϸ�� A0;Ԡes3��ڦ��O�[?1
g�3���kO7XT4ޗ7�#��:S���i�tPs�	��}.t^�|WG%�I��u�[4%B�P ���/Q���Dy���~+���9'��\s׀�P�,�-�5�J��!���%��_���٥Y~5,���+0?��~�$���
�$�I�����ҲD!}�����ّ�r�Y��(uy���CʝSW���`�u�)��v�:k?VV4К��/��b�oT��`5��BV�&`��Y�ܶz�v�l���0���n��<��ir�K�d�g�bR��V��.��IO���\Z(/�J���Q�oD�����.��[�{���g�kr�'d#0[�;[sF�����!���%n cY<y�V�����߽%a^�	d�� 7q�냖'O�z��4��ެ��{ف���c��
�r�����F�n#���7�y�]��]���;v�.���v��/�$�+�J��$�����};?�"Lm�0�i4����6yr���'�+�BZ/ӳb޿$����(??������83֮I��2�(�[�.ִP��'1�7��O�96\�rI��ڝ�Ҽl0�w�4.$g�cRT��X�ۼ�E;8���X3���<���쀤:8�h����0�P��b�{�y˼�Q<��u�?C�J�
	�7`#��<���׹.�Sl� 2ߛ�Tr1�A5�}�9=GR���z�O\_[fTS-q\�z�7η	����:��I�z��<���M�Z��=X���dQ�����������W' �Ux|Ӑ�kϝ��T�mAT��$d�}ڏ+'Ӓ=��!�v�蔴^+��kĲ|*�q��~�X|�]$Ϟe�:s Ai�j0��jQ����?3#�YǙ!X�Z���w<�咴��5�'p�j����m�p�2m�
�+Iu@<]D�B>�@����5m�/� s���q��j����҇�3E���ٯ��FD�g��.B�� �1�G-LL�Ο:OlK����#lG�
j���ow�D��r��_���௚�)'Hȩ)�Е?e?L��7��~p�*@_��P�D���6,��Gؿ=l��[��S�|��w���9Ov��Ʉ_�g?�w�4�+�q����8:����eZ�Yd�]#ˣz腸�I,g���_�]L:�� �K_�{�ӷ���Ǩ�|�f�w��8��N	�ؼ�g�zC��	Z(.OJ�j���V��}�%uI?Z���;=l�	IM�\�Dh�]�'�r}��lpF�ɧ:��X��BmH�6�鄳�XT�m,��@��۾��R�B'�6�Ѥ��>m�X���2���#���ߞ�����-�c��굫��"z��;�Dd�3�킻lO�`Ɉ4;��(�qް� 'J+�QLP (����M�zb�t������q
'W#��-K�)=m	���Y\���4�7��zG�����>�t�8�<zb��7�i���kb��t�
NZg,2���f��[g#���-w5���6�'�wwܤ�gH��\�����"�VQ�H{�ޓm	KB/���,����H�˴��y�aL���6f����.�e����]y�ҼG\��#
�����g@�P�8����c��U�H���ʥd�G�q�1��2�V���b�1�bҦ�CS�9�Ҕ��85|.�ř�Sˇڗ����v�-����.����<ޣ��z�N�F�+-S�iT5�K�h�&�w�P����<o唡�;�.'�����Z�m�d�ƵTQJ��Ck�k?��p�W�L_��nE4���Y��a�������@;"�f|�=���YS,�a��_,���lH�\��o�v�6�X��)����2�
�5Q}��P�U�!�)���O�3SZ�t�����w�i1�j�j�9��["$�~X��	+o���u:�)#���u��j_�\��!v�������Q�q� �9`�`H6���h�eg�+��C�6p�3�3{�G���@��:����<�4�]7r#���UFCl�v��D� ;;�=Μb�b��/����*��C�e]-�ZE{b�J�AF��y(�w|~p)	ɇ��L��P��	���;�G{�>�@�l�j�A4�T2R>�M;�/�!�`n�G�1��3�r��h�S#��"��r'���0�������VG�-Y;��r������kM#fq���녖+�GE-�*�KKv����j�ʬ���0�Pwk�vT��Uv>a/��׶jA��jU�[A�6���)7����pֺ�c�"
�Hi��6����i4�<�^rV53�UbѺ��ʹ;��0�Jkh%1�hD�nFn;�{�B�?��,|O=4��L�b���|W�e?���C!��Q�zc1ך�?�T$$���P"e4C����+�XA�V��:Gg�~	��M��g!��D]=T�ֶ���?�CP���D���2{�Q�3������ܹ�f��������9� �C���l�֩�T�����	�
�0j#��.F9�7B�i�A�yo�Rg�#�r�o�.b
H��3��&�ͣ���Hi�7��ױM���p��RB0��{�q�8Ԣ+�dte�	��'M�c7'���C��.���d=���E�Li�Le���	�(�Je@���=�o(}��D[�`/c�dtt�<�ևK㵇����@=��mϗ6Ao*�E�"� ��4�Ѫ�����[Z%��E�:)x)'#����9V_j��M���Č�V��X��	xX�ǦL�a/r;2@�t�bH�q����x��`�!+S�Tʖ�n7hz8��$����$��c��%D�c?촳�5�eg�"g��2�*!��U r`���]󲆫�4<���.��^M��~�}�Yd�a��%8�:��N�(u����D�W|o�9�'Ҿk���ɦs�iC����?fG��?�.�^?����#o!�	o�RG���/��t!9��-�A��O����x�%�t��P@���˹�c���5�38���)	��
^%�M:�Mz���&a����P>���d�m��6�!�~��@���Ͻ�q�Z�[{�,A��$21�m��g�$��u�C ���Hi�wy���?�j�9��:�Ũ'p(�׋�<�N���Ω:+�J�a��й����!�<]~���ا]�����̃R{&-
�K����tRO.T�\�!9ݍ(P����xI���v̈�2w)�IY��ȕ,M7m��ɚ��R��R�x��1�6T)-�TJp�$���HNrI���v�Ч:+���Rf�\�_����8[�(��m��$-���2��έf�U ������1r����4��g����>�,���oa��R���8c)Q%uP���L��ei���ƆkaR���W�ʱ��ˈs��+\�I!͢�{9ZZ4�_'<���S�+��Q�okp]�Pe���:�{i�A��8���e�1����y���Ö�ds�k8��P���=͢���IRe�s4��;����k֦��{c����w��L�9�}�a��q�x�t�I���N���X^`�0��K��GF�W@���ގ@Wt^���v5��3�F%(ɠf�Z�ҁ���/1f��)����:L:`l0g��:#�+nNWSA'�� 3�Q�M����p���7p��ր��(�h?��Z��vY)���0p���O+����.���g\A�̺�%.�ב��.�c�p�Z`���#�<�
�`���P���S�_8i��i��U��5�	8�A,)?�;u���z��sT��ʧ�O&�<�ID�A7�� ��я)�T��e������*�˵�sy���JU�3�$��z���ٌ�$1s�/sk�<�������:��XLF�S�d,���$�9"�����C]m֫��LVa�C����)�t��%e��BE�&�c@*%8J�����˪��8 '�'�E�Xk��U�q��̐-�ΊEvIfFRO���1��X���p����RV,8���|�i�@�����Al|;��H�s�����~�\Jl.�\��a�k7�3Pp���Mh��5";��n��"�E�:0�*Z`�� 7�P�؟�ʁ��j�`��A��U5nA;�	���h{W��ˠ�v�jbJ�E�^�H�`����8�� >��j�8�u��`+��ν�u^�F��$�X1Lyغ��j97��4}>�H����R���8����~�j׾������8Ԫ*��ñ�c��m��n`7�.��+�{gī�P�A9տ�y|�sSW$Z��EB{�DR�� �����4.~s��-ߊ�G�.�sX��dP	��uo���O��C��lņ(��J�o�pA#�Ȳ7��Wi�m'�d�CO�Q���k��-}��4�#wfŉ}�Lfΰ�CZY*��u_Д�$>j9�oX�-�~�H��������n��=nfH��<�(�1w,��P{�,Ph
:m�D���]�
��P�"�I� A�y�����(�dS�t��%��;"��uL]B�|c���M��r�C�jϴ�\ �������?Q� �j���⌓���){}7��b��� Q����DJ��;0��;����*R
��e���!������f]^�!�;V+/%+Qp�C��o�6Zod?vQv`�/Qá����z�(�D9��omsP�z�0�DE����ز�+5��+�O�uA��W�Ύj��(E��M��ҳ��;-�7n��W_���	eWQ!��Vd�{?}{��E^�K#���XJ�c�ƓR��#N��f龥[�=f��2�J����?|'�C��Ve���mk�(��s�ފ������� {�ul �i�  ��h��/i4�LO����;�B�� oI#-
�u�||���1gHQ���U&�D���K�	�j��CPJ��('
K��b}�	�r�'�����J7�K/5P@��л(ѡ3QItƄV>w��D��:X�ᕥȿ_nތ��{��Y�̄��Yd��ŇK���?ܪ�*X&	�+��� ���P��|2!M0z���Xd>�E�p�""F�R
+m�N*��q���ּ��#��pqԠ�L��>�G��L�j:��1߃�	�xN^B��H��<�i ��84 pRt!��u�R� 1�Kv�C0�v��xCg�tق����!«�<1E����
�ߓ�L.�V�?�����H�2�������������g�G�u�A�Z�ҝV��<�8<��qx�w�6�CYm�a���H�dy��}bt����K�9y�����>���į�#P���܌o�o��a�]��іz��Z�1�,�Z�����H��]��މ���4�#V}A�����}Y���ӿ� �w�X�Ey-t�7<��ZtM��us6������.5�S������>q���E��%�����ۦ'���Y�q1dz�?�`�M�נM� ���nº��߄�I>�[I����}�J����	��S�SiيK,��%��R�<�OVp�X"���}���hHfya�����9t�u�5H�� ���5�1q��!���!���p�H�c!P,��w��e�ݷ��Y�\�p%)Q�/�T��yt4�7VW���2�lG&�2����4'��<��p�� �m;]ߜ܌��h\W���p�V-��������盐>����i�O�ط��A�m�$�uF�ض{��ɱk�t�E�ۋ�A��!�����7�?V�9�c61�~��gL��<GeK��t�b��!j�����8h^VbYCJ��K�`� ����7�.��-Ґu��C:�7�������3�=I�'D����mE���!����wf:�h!\djf�͕�z�`�e��q]o]	Tm��rC�@P;���bc뚦:�o�B��?�WJ,�r�I}Up'�8/ ��$���� ]gX[�����	0ʋL�S�����$'|Z���+�����wY8���	�Ɍ������?��^���$�8��+�0�=߯������i��cn�8/Gx�8�;�z��%o��Շ�����Y�s��,�]�`�Q軤���0u��Ib@USzd���ە%�C� c #���(�]�,���إYE@�����~��[(�r`�-�zj�!����A̜���7%(�ǀ�,�[�YҦ�Õ�(�M�>MO-����Dbf�z�� �i�H	�O'Œq���U��s�{�,�Q_�;Z8r�ܱ�,B	['����A�2'��#t�֥P���a[���� �)ӁV�D\�:���h�ǋH�C��$6kV^4AdE5xw��IjS���L��:��陦�G�ks�;��<!���*%:�=��/����!���K��X�X�`�L���s�G�����&�m)3��w(�O��q��Nx��$(��=��|�+
B|A0��#��G�D�QI	@;�7���]:AG��y4�$�C�`�-��מ�8�^�1�@v�3�2I�F���%����Q���S�L�M�F�v�i	|�dS"��������K ޟsF����g���7JW�|h}6�Y,�x���&�謠b�����C��->WU��J���;�R�]������'q�[��g�=����$�^V�C�^�;Dh��A+^ �jpD���b���X�;��8�UD�o�±ڎ�����ޞ���˃��v!$������Ⴭ��|�?��{o�d��+mi�]�ȩ}�ʦ�޼3�����4�M1�ɉHS��3S1}�W{���wTQl���>��!֒;�q�Ӿma��&	��>�W��?^tP�P�I�n8��G{��l��;n�@Jؐ����	*����%�S/M�:�zģ/�?H^���k�}����� ��3G"�+�S�\?���;�i�1Cg5�MΌD��3�%�w ށ�`$���IH����o]��*x	qOQ�w\|u�F�쾃�Pmµ-��'X�j,}&�G@/��]��ݥCzF%��K%��$���Á�I1L�S}��e�>B���S�C����������x"��[��}�b������<�m3������8�Q��R���.�9M�a-|1��9)�B>�@[�	��p
s��)��������
ub��\[�����ҍy��=��BU�+�{���<Ĉ� a�W���P[k��c�6s"^~���� Z8��iQ��Q��G�� ��G�`�ϛ����-��J`^��b��<Vx8
QW�b$~}�� t�B����"̒�h{?ʑUU$3��:�d돘����O���Y�c�Z�/�DE������9���׶ml�f>��
"��Fh!-W#Au���K��p=������7�Nꨲ�h"U��ٞ��Ub'eϷ��~��\�ң�@��X��@q�X�W��� �5gк)<P�k�يGk��qw���=rD�|Y���d���9�!y����\&�l��0зK�H���ت�q�����j��<\.�1k�cq�EWp0'B�����&�-��|Q,n��z�M
�r��D����[�s ��<}�����2��{�OcP]���8�A�YO�������&z�������h�5*�m��ɩj�Ed��x�m��Ȉ�o���GQPZVү�����Gn�VwQ)0�_~�VM;L��4hl���^���i�9��&��D��JWm���d��j5����L�2���<��7{^;ֶ�߲��8��!������8k���f�Q=fN�Z�%��>L�M�eu�`��AA����`��A7�t`�-"ބl��O*�&`7Ń��b��J5�˗r�pJnI�Ȉo���gj$�'�d��T������DN*�cP>����r(��]ŕ�y�(&qPB{�ni&6`[	@"};¢o���Ss!�$lc�0K�` ��B�Β:�λ��kw���M��v�s�C
�DD9�M}ELv����n�6NMs���4��� ����i�f�~�T��l6���0�蕅-��`��i C|� ��m�_&��傁��AZqg���y���1I�朷��G�=��p�w%�iH.g�{C��UX:�7As��Y=^n���ñ�ٍ���_&2��	�>�?���٨ ���b�_��o��m�"�d�hP��}�kɴ�j�6�'����!C�a���������9Y��̬�Y�r/���ė���\�\�J4���D�b�>R+H�\���I�p�S������h��2QO�j�֦�>�Qb�7=í��Hw�lL�Wl��r�j@����%Z{�1�ؔ�g�7�¤���U��O�%��!V�NN:�Bbr�ȹ['�֯��{4�ټj�A+܃�����$�1�i�9 = y���䊢F�-A�n�/xzPc�^(6�N�@#sC��ݞo��Gv�08�ta3\쫼���˫������ �c��b�������\�`��2�`ץ�]yM�i��(2`OA�7�!�,8^<���B�Ū�rC�G�����K�T���ڈ��c~�@���L<,�ΪEǫ�)vC#T�l�1^���VZ���n-�\����ށ���߁I�ZwZ�����j���p�Б��%	
����@K�.}&�d��(�un��F˼*�{����Y	$u�8u������Bx*�0Z��Z}�����_�?��E�U��Kr��;�i�"�W!dZ�j�'u�"���p@^��_�A��`�����z��ے�~�8� Zb��t��#�3e�;� �qƮɫȅ����BU���=�!����d�Ca��"X��yqՀ��W{��vϟ��$H����E`�t�?W�{'W�q�Ⱦ>��eO%>�]���ֳ[|̂i�`%�̑ԯ���s������0I�٪:-aM��,9�/�h����TI�)Lx��vU&ދ��!3��,���y�b�5A#x���0�	;�S�=��-��(p��[$`�Y�+f��*�*T@~E�M�*9�8n$U��<=�s6x���4�����ʍ�)gYI�{���S��\2a��<XMr
��M��˙��bn�_PF��Q�H�bY��f�"A2 t�h��ɡ�O�;���%?[��O*o^�I��?�o
�=
��s �!���t��ff�ӣиRc�����t��a�.R����-�T$�E�3��_��]�o�%R%˸g;��[��7�s�҂.w�#�	,>	!o���:���[��\�~�ef��z��!%?I�$,%x%E��"��`���1�L��oK�{��@�2��O�U
F�R��,��^a�<�S�Sh\�Y���z�q ��8�/4����:�!������n�����׎>%�b�?��o���#"x;�)�4�o�F5>��T�ʀ_�{��D��Ç��i� ��э�9m�qV�y[���Z��P(�B���u����c�����'O��Zy��Ѧ`��œg84�)��I�� |��n�pm$�۷����L�����\�����>��x�K���>�z��?0m��tM��������J/���F����l#��и���(��4Bͺdk�o�˝�Iʃ�Tt3�B
�C�iM��W�P�L���(���(�ij�P�k.�e.�	�³�v z��"#�x։k��#i�Lǥ��l�E) b����Xk�;�R[Zω�mL��|����Cpf�7��Qڋ����S��zB@!���A1��O�͢GǺ����$-��d���k�.�Ĭ3�i� v��+O�~���v7-������А΂����� efq;\n7=���ѩ�U�X6a����]��yG�ǆ�c�w����a����O5����s�Y�@?��~�q���;�|w�"E?-�7��F����u.	�w��'T�]����<oDSWP�d͹������K��o[U��^r�R����@���&V&^7 ���M�ȢV�?�t g��Բ�D����Y������Ϥ�D�S����_&x3�MЌ�DM���^s�C��x���Pgy��!D�z��&�H�5&(�0ڞ	����Ԇ�� �6�b	���DDdkJ_�(�pHI%S8����S�0DZM/nh�������;��2-sP=��i�m����ٲ0�pCH���Q�og>-.փ[���_���Ɲ�����ԯc䠡�.��rq6���}Y��j}�ׯ�VE�J��=d���#�PtPiU���C��ǈXD��I�M5B��a�F���a�>Z)���i��KV62�<�49�b�\��.�m_˻$�I,�mW�9q^����Z�&e%D���b�
4���t#Ԑq���(p�c��B�D�=�*�N]y�W*�B��/�
���F3s1V'C�آ[��޵ĜZvBkJU��(�xx�;���Z���3�I#���P�� ϰm  ��a'IU-��Բ��HFo�k�I�7�x�^qÆh�O��U�P�Ѣ1��5HJ��/�W&("�X��ȷ��X'a�>YiqSz�+�t�g��߬92��RZ<�U�Wge$�!r9��WX��
������؊����^��OP��z6`��:�~�Gk-#h�^��v7��ɚ2���	q_�Q��a�����Ӏϕ����:}���-ʭ�l�/C��8xb+���VxoOm�>��w�M���P֛�*AV��0� �'�F)^�mAT#��
TM+x�VOC�Z��y[�N������D�����A�Ϟ�a�['9"`ۘ�5~�|+����n:_�z�V���p抖Q�&�4�!0�H�y���� eF6��?� ��S�R����
M�!�T��t6(����s�@���;��b�"�G$e�����E$AP+�.6�#�r���O�8�w򎃲8��>���ZkR��)�+U�=�V�Q�l�m����^�xxjN�(�0'�U՟�\��?<O{O���͇<k5HK�Ej:���G����d���B��N����Ou5O�ʝ/vR�Ƴ���A
:zNG_�m�Ҭ�6��j�\�N�MYJ���-�y-Ұ]��"���+k��H�&B����C�Ua��?�n4Ҝ�g��-�D&&q]���֚���K�x�[��Ô1Eu������V,��[&%h�&N�[���y�U/3*��APћ��@"��:�;Gp�����ވ���/H�)�/.�k4�R��N�G�!�ݠC��>э���&��{�B��z5����}q�|���@)4�T�\9���R9���L +{�ؙ7�֍�V��H6��P�N�`wD�`3)/if�vk�'q���D�"Ґ��YXT�Y&�il� ��2<����+���@)��Gϸ��M�PG�Z�o��qk������X�+�L]��E#&]�����?S6�)��@|uk=��4oږ�UL��U4bF2
-یI$eZy�%&}u�Je[d�"���,�������SOx�
����q�!���g�^�P�i̅�E�9s����	����(]C���RM��|}lܤl+�p�O�UΪܜ�;��M�:�{<j���nյ�T��i	��u>#��y������K�󯿌Ϟ�O3/��9�(6�|�A?B�^H�V֤οm�֝�K׏V��[�}$^��E�P����G ��V����B��-0�)^,t��83U���	v+�l������ws�{�%��E{�a�^��1�&����a��%�_-�-�wB��ATO�<cX7T7���Λ7F8(�ڤ��W+�h=��1���C��D(U���#Gs��H4�,��X��u�OU�W�Q��Qo���7>��($�������٥��~P�M'�m���4J7I�0t����dJ̼� c	ѹ/v��̲9C�S)���s��]qK��q��/Y�ۨ�Z�	�(f����:���G��i���ic/t�ld�W�ͿÎF3�^�q9��7S[�%���z2�M�D˕>��$z ���"���c��J<�����Z��{��y�ȺbS���UI�t�Fe���w?�����vv����3w +@�z�Ô��	�
=TO&j���P�Y9C��@_9c߉����Aɘ���*m�O��uqۢ
��!�Ǿ��Yk�υ"��9%p�hMy�����ꝟ6�ou��I��03��t�p$�q}��||���u[�^����;�'��a8A��m9� {	�E��b!�)�q���RA`�[ra>��\�GXƕ���<'��adn�S��R����a�����Z�`����m�&��0"O����+�U�ԗ�FF*�:�	�z^���t�>g��E�O^���T{�kS�\�Ui"g��CSө�%QJ���Hf�f�,?�+2�J;��P~l:�M``ǯ�h�C�C�u�������}�*�+ ���B:�H���ˈ #����縘������S�p���,}J`���&#��f7<�,�t�74b�� �9/^��fq���(�
<u�>�X��	t+�\h�:j�V�����
��Ckΐ]����!t���A��v��5������6`s�șIa����x�vl�����آ?H��s��d�݀H��o��کE%v��y}�s�PC���$ظqW��M,mXg��uq�RE4�M[�M���]fLw��ŝ10����I	�S��i_bl�
���S-%����Dj��d�H΁��6����y1~*8kUw"%�3W�f1)�}�>�&1�Z�J�21����yV�����[�P%aDE�ˌX<.���nD`�	%|֜����o�8������᷺��Ӄ� �̮���
�w�Pv�G�ѳ�LpUΙfS�&[�R���c.=ך%}1,Կ�j0� ��6��o]=���}j�Ԧ�h],,�?J���8��R�?q/J��zK���W�[�"�0�Mk��	Z�3��1��b�=�R�����c�q���2
vR�-��x�!�*��i1����O�"���qx9��q˳��RТ�|���4w�gK�i��h��e��$pB�!E�ꮹ9��\u
������yZ�Za��ß���dV�=t��)=���.IP�B��g,��sd���5�=�7�� �!��*=�,��L?J��A��]�*��j����:*P���e�!�5y�._`�3nA��d�5�c'�@�����
ڪ���88�쪰D�z�*�����K��dF������	�+"BB#2]<�|�}��u�x��G���W^!�oMB�1GvT��<4�
��	Goi��˸i�g񮵻z�N̚]A�����.��{�,��w;�Mg��4qԵS��m�%Q�?"紀h`��\1+��H�P����Hz#��c��~�6^Zu�G��@���D��@����M쐠�M`��)2i�LAL���h��#+Qݺ����;�	�[�2&	�����&���
�~8�֨^A��~.���ί0����s��.0�!��ˈ�#���K�6n�<�A�#Y��\;�BHy�8Nrs�(E3w=�<�׫���|�+�2=1U�gD��.��Iݭ�Z�;���F���i�{��j�ry���Y;)�ωF��,W\�2������}O8���L|?/ɠ	���	�V�!�ߡҳ��L�[��������O�[p��g�+F�W򇆘�o@zα9_�(G_[�JY�=V?$GfÏ�?*u%�W�JWv�LZ���g� ���.�_ c����D�
�d�S��V�|��26t�6���+y,=�7I?s�'�> ��6u��=�Mpվ��i�Tk���R�{YɴoK)�q�<�J��"�.<>�����[ ��^fL�*����)݃�n�/J��+i�Jڧ��'J�OeN�4����Q�-b:/�N/ �`�ZlǨp��ݠ��+q?�m���π2��s��(��\��躪u+�`�!�Y�?��l��Y������Vd��h8.̐*�u��8�$���^���/Nc#Iٮ�_�TU{dV D��^�(��>��N"�{_��������?���U�7�P\���@@��R�!�������F�;�/e#�=}�.��h��d�xM����pP���Iwn���-7a����Dz�{_-xZ�C�"�p�V�2�(ȿ0�
M 83�m���
	�?���'kqD�@��ē�@�U��!�C&�~3M	�X��ha��Y�-��j���z�&�����&�\-��Ȫ:����Tڦ�ge4�,8~��
F����>ge��;gԄ��7�#��7fv,۔�e��z.��,&�����N�'��Y:a�֬�U�H��7Xm���e���D��r���p⌅D\=�.6"U���[�9z��v	Yy�8���¨��M7�3BQ엲w�A vV���ŉ:D�������{�*�^�XXRZ�	,dWC�.�ВHϲ}��v�#����&嶠����Bq�Z	n7�a�đ ��Z�������=�n �#:�C�0E���N�3��~�@Upd����� �''�Ts����u"߁qF���~ڔ��'*f�e �$�v鏈%��B,�ɻf3�әO�ccs?um���-õڏ�\ˊ���B��pܥFPT �g�,�:�;�E����.�N��M�*���@M`��7p��G��5�����{#Q#M��'$�p�������]��	;!�"��c���}���}�Db!w!�Xg/�
�5�����5s�k���	��O��Chf��\\�!�0köQ\xJ]˥d��u���F�V�gI�(�mq��/(�i����zJ�C�3����xS0���~Z	����nj@�p?������ZǒCn�C	��Q1E�H�'�H��]���f��܀#H��_��x>��0e!+�޳g0����TN3�F�����pK�R���cj��Q�qW�+p���e��0PNb4��泣��&�dD�h?�$���?������f�n�ȂO�B߳�Բ4(~�n���X�a&�?�|&lr�v3���B�B�x�5�MȄ���-�j7�`�
}HwI"����Y4��=�B#�oN(2�9+�`��b�>zk� T���S�v�4.+C8��T��E��cF24/4D<to�� �r/�d��jk�x���ރgy�E�܎�p��>y��n����=*�Q.+�9K��r>��2fپ�~hŘ��kP���ۯ�y�k�Ϩp�����tL`�����VGD�������j�΂�c�j�r[8;��:C�+����	�j>�� v.��f����ZP���iJ>� ��o��_��O�b���E�_9�"����}�k8�\<��E�utw
���3"�0�俶����#���|/�[Y3�"�����%�`��-���)(~� ?��J"�=�ǧ=u�����H�� �>�'�碑=��3T��(��lhe�=����W����)�l�D���vԢ�8����-���)O�s��y���[y��}ǰn�3���j�z%�>�6��y�� ��?���
h�a���Y��,)s;�A���V��BE�$�9�'�H|q�?@��t�Z5�;r&��K	����s��O��<+�������K�S�I�
 T.����_O��g�����L ��)���%����O���[����3%�P�Jt<�@_rvF"`7~��I��7�'Ζ�j	�_�{������&V���"��G˦jM�@�c9I�e���ԙ����h��s?h#\I�;�x~�=��˦�����Om��O���gZ3��4��vV��Uٶ�SE�Ґ׀e}�Y�Qj�fz_QE�c;�O���$�W��!^�����*H՟���v�5F�4*���� ���q9xkm���8d��`���l7�e�矓�2���%M�7/W��s~��&��)�QY,�8���ģ/�мwІ�7����{���A|F{l�K�-���G*��Pp�5�`�6���q�@��G9V�;��������֬�I~�aɌ,�d��Ë4�Rk?�KCT4�0�đ��;c�7,�*?v�p���F�L�~F��O ���Z��u�Y֪�SՄg�a��G�O]�G��S������c�U������2�M���o�bN��1�a�+3���2{(��FٷIRe�UP/D��_����2����޺S��1
|�t
J��y����[�	�'�qd�qk׋����
��4n�N�	
��)��.�%B��;��`4b��05�EB���A')�b��E���Jb���f�`�ܧs�^�}��{��t�[G��O�p���tL����l���Q�U<a����%�Q�����SI��ސ�ĝ��eF��yz�����]6t���H�G�낏���ݒ~��ب�e��PgG&�Կ3��4(ڔ�����:��i���) ��Ԓ!@?���UO�74��8hO*�/��E�j�>а�vMw�R M��خ~�)�{2���@����ft��?}U��O$�78A��3s��������	�I�H8�Eͫq��NW�����k�Ճ>Qz�n�X_fQDϊ��P���WDK�k�8k
�����,/,
n�!����%T�v��ܒ��߭����)T"T'b>���?΂?d���K���S?�.��s��qK�.��f�������I�X���-Ar�
��kg����xp���1��'Sr*�Hoh,�ivZ<��ʎ#���X}eK�[ڏ��[�O�2��~��Z�G�V:/��7
���F���9���Y�ʢ��T��mS�Dzz�̸��ʴ�[��
Q̬�c�����OUIP�T�����=��t�Lkr��sQ��K���Z�[����;�h��]7�Z[�^N���Q�):̏�9N�����8W�-gG��j��Es���9/���f9FT;Q��GH�h���6x�������K�xN���������k 3QL���2i\��+�Lʴ���n�i,nb�����������T�������**|c�N,$�	�UO���׻x���ί�B�4�8���X�ݐ>p�Q��E��fN�Ѹ�]ɀ�j�zd���$�2�����V9�i=}�ò�a�O==7*��A3�~Ѫ<��92_�T���G-c�n�0�"�+�))��D�&	l�}�<��"q�D
�$j�R/?�@�pW��<��/G�9�q�<�!6q+�e���K�|ӶO�k �k�������2����,�v��*�j9���1����
j��楢�r>�@<��#%��8%2��UZҙ��φ�����\�x*)����i`Wq�ё�$i;!�[c\W�v8#I
�Q��
��)�4�Td2�Ϟ���[e_<��QW�6P��&<���3MZ&�P�Ml���M��4l`����-w`5���&���u2$��Τ�@b���@�E^mOi\r���/��MJ\�C(�{cemX�A��R�d  T[��K �xu��Ө���Ta]�'�D��G�VËƖ�"8.����d��l�<s�>�m���x�&u���I�qC��A���U��9����������U��=�F�R�w/U�Īrh����짰��4��_@c�����u��'Y	�D����(I��"ˬ$[ߧ8 Vr\e|��k�������_�g6^,��9H�.���9 �� �1r|%��� L�r3��R�܊,ݷ�˝]�NEk{�s�KX��F�:Q!]\����S���A��_�6��cW�=I.���:�.w�Qxha����vg�m��D1�~J�%�R@C�ᖟ}��W�`�D��R0��ǐ��b��K���j9���9�m%��M��n'P+�?}�2��SO��w�l�+�\bb��/��-���8r�+ u	!ZF��A9�qcZ|��G���T�c�"Y��P5|)���@��O};g>ev5,����H!�4�#��a���=�����bx`W��/9�	|�P�wLo����6R3�d��j�{�M��	z��V�F0C� �h���M&q��8T?U��nʛh��W';���g�jX��+��Ŕ���w���o�Apa�٪ɹ5��:������ ����s"V�XS�����/_}��squV�0�Q��y�KU���:�ǧ��3��:\R#2��EB��;`g�)���G�/v�2Z�u1i�wgϸ���~��O��";m��wf�iV�q�a%=�p�iN����c�]�NP��]����eJE|.r�U*����K���r~~�I~���d����ƨ^��ϒ���`	����O39��Z���G��_=NX�[�� �a�� ��3iL@:�*��I4�d^� ����	�{ż������6`-d��(��Hv��aG���#����y�bL8�>�� ��C��AZ>&Z|�����A�c�p��+�F3��n��U]��9���K�d��pR\5���P{f�N�B�k��qd��Ю�D���=����R1F��E���Q�Zh\��.$fi�`~�:��@��^�*�D>��-�l.L�)�ĉJ:R�y�Z��
,E?�#m��{���M���u|��Z:W}�>8��+4Ig���/���vp��R����t�P#۞#v�e7X�1���I1N�u��\�LF����B�8��
q�fC�
��.e��y�D��bR�K��Se+���ܷrsm��#����#�~��y�/_����K���CI}�lA��Q�����V�.������<�l�r��t�|�/��Z�-GI�XU��@&�?�Z�;=���v�oq�����\��kQ�NJ�����r^�����Ci��c��ǲ�Q kH�n�³c��=M�-���`6F�J����e
i��}����|�^����l�6���Z�����>C@�����R�{]���0c*��d�r�s" Q�ֈ
�(Ѭ�����v��-�)�m�~�b���3.��S���	{C��3C' ���ܼ���3��Ok�tG�/%,.��J��~�(�m�ǡ�E�:���p���kIяf��9����1lr��Հ�gL��r)$5�L�6d��=>�];���\��6�,j�PDߌqV�� ���h��Q؂}�'�wT�j�m�8�]*a+e���?Ÿ�U�(�6M[�~��Ta�*��F�����+L�7ǲ⁲��'Gw�)V�;�|�K�"��C�C��s���X_�i�r�J�Jr��o�#.�bY���tr����|t�qo7�\��fk{峷O����J)�D�Ġ��h�P�ϼ��/#9G��M�	|oY��Ϲk�����A�����(��R�v�_�B"���,�+	&7���j��+�أ�s�0����׻C>�LPWw2��j5Lo]��Τ�A����s��"x��+��8Pb(p����;��Z�;Tk���]�)᲋��s���kc���xsL�N�K��/���'��>����_�R ם3_�~Me�/a�:	��-�0���/�&8ž�m�"h(���&�W�V�#��9dܩ��[7MG�}Cg�ޏR�0Ҫ�ڳ{P�"��� ��m���!M'��(��5��?�Y믶�}	�Ѕ�3_8�+�܈��=y&+�M���C�
���:�e�I#��3$��Þ��'a�p�"��L�΀̕�3�GS�883�<{�D����O�c8��ht\ӂJ�R�%���2E0���[�,�ua�wRYO��*������	d�:9n�4�G�U�,���z*5P��xh}��쇗q(T�%���k{o�����W��_����Ky�,4tӈ�q�sz��ǚH�g��h����^��F��J��:�2������y��̀�dIr�*��TiEj�	����Y ���:���Mœ�~��шMe�U[粧���]���5ݞ*� ���#�ճ�`��dL��r��:=PTF���o�����?�HFÃ��/p�]����)�Z��C��LUß����Z�" ��
�c�rF��X�f�qoTԮl��AH嬣��C�j1S���Q2�����J\��5�kT�����n󭈽=���'|L�Vt��֨%=���B.G�ߴ,��p�Z�w��פȍw�8\��=9}5*�O�%3�ő��6ީh���X����_4k��d�i����o�S\��_�<~)�� X+Fo݁̎��,��T鯞����{!+	I-n�ٮҾ�Eч�ܘY�% :�M���� ��H;+����7��.�yq��i�^�}j����EZc��x�e�cc$��f�ok�f!����;�>'%r��A��Nm�P�!<<`K'ă�\�_V���p��w$	��)���"���R�1��_MƄ��Z���;y�N��y^'>8�
}�ڵ�]�����U��+h@ɏ��%Ïo�7�>9�{/�􎷞.�X�١3��������'<s��k�R������z��Iw�\�kD���t��u�hw�+�����ȯ}���}T�Es�3�D*�}9ғ�����%�[�����5d/�r�B�ąe�����F��vƚ����{��A�^��zV���Xb�Q���W����ݍr��b�	����D�^M������>�5��@�#�/BE���0�+[�,d�t�*�j��+UWq0lg%���Рm����v$��fᠻ��P���%�*t:�v1��MЅ�!(7Uz���,�T!�"Т��М�*!��c��<�sC%iF0x�R��(�ޱ�=���s��������)�����$�-S�@5����8�ef���סt���9�����m�Mz��� ��2ݤ����~�d5����MǛD[P�pp�F+�}.�E�Ƈ�|(v�fÍI5[V'	Me���z6�>L8Z�;6�M�ɉ�S��S`���aA(V� �Y���8���2��I�]ʮ��#�q�g�����-T��F�s���z�&N����{������@5��f�\y�RU��[�_�����Nbdj�z�����T�{ ��5�v�s�4%f����?��V<�u��́�:� +��k�����r�c�f����S�� �PuH������~��|R:��?f�#��>c��4���^��_�@���o>Y��_������R!ĺ�(`�T%�t�#{��_ѱC�̣Xn3_ t'��6!�x<�n��W9Y2>��u΂#!�)x	v"�H�-�yꁨ���굴B�;�Ì�!�j	�"��Qa �zM�b�Bmn�Ĩ6|a��A�u9z��M�`jA��I�g�}�X�X�ց�hj��y�I�Φa�;� �o/�^��p��[�M��˽��mڋ~�]t�H?T�����nK�c�ˠt��2�Bf�.(�:2�	t������S���GrO>k�e9��%�Ǻ",�����U���$�?��`{YӸ>�@�WY��v�sO6���O��G�8�O��J�����C:���D��_@�P�l)W�yjUm05�$[���K�� B�N:ѓ�����y�B.� D��p&��Qm�M[���o���l�So�iO)�1I�~����O^�s=2���س솖�.��f����=�mcy���|!�,�>�p��D���:6^��������ܢ����M�A*���9��Hz��\�r�s�Q_��ԱA�7�53w|g\Mq�a��.'�1���0�L��%�-�=�8x��j>hok�Uv[5ZW�B*�X��g2���(L�*�<!GiA���78=ܧ�
}���U�#q˞�|���,��@B�Hi�1\�44�4^d���璙�i���L�|`o���(�����6�3z�S���̊N���Oy��.�S�#�y�{(b�q�f��08���PT4�3������5گ�j�xC�F�Yo�&��4�b�-
ƾ%>å3L[�fǔ�X�t������G��y^8N��3�) *k����e5��'Үv�%vu�C+T7��,4�{�}�����u��w��@���hYrf0�fY[|>x�1��Hj?��5�+���ֆS��1�Ww�x���{D�!n��|�CI`l�v�v$��㡥� ��H�}61M]bο���I�&ί��Q�PJ�����6؊0D���F��������q����I���)�p��/����u��'�����RK�;��8P��kTI0���+
���ޝM7�6��%�P�vE�|�se0,���P'���*���NS�z�3��Ƙ�%��#7��&���Cb�Q^�%����UN�mx<��^g�:$���/�}��J�I�4������V�q��M7�¶�v��j�y2�T�ť��E�̒ڍ}��q��,N�����!�i���0�g+y~�~8n�=���&�ó�\�C���?:q����=L	Qݾ�(��P����zܯ೟oh�lNI�����rˌ
f��߳�D��Q-T�ټT}�9n����MzS�]�3cF[����_2�Q��*z��m���#�%���y�����L�uc'�{�⠙�)2�����`'�Bb�fm��i�dh�0
H�ϭZ�ƽT���W���ep"�K���
�3`�%��S�}F�e/t��~D�Y�M5��^F���&!��7z6�9#B�Ha׍*�ѯ�ĥ�M�Z�Xe�x(���p�Kҗ�: יl�_��ى��d����m�>	��v�\��k�D��`�,�}z@	�OS�fN�~ 5�Ô�p�v��[6��co;-d���n���>,s�Niݲ߽���ާ�����4"�Ø��J�zV?��!Ԇ����sޜw�v�p�],^ʋ��Kj��,[�Z�G�h�*�d��Γ���_o�&���������w��>Dw8|�`���!��v�^?��Vc�s�s�����8�9�Lpf��ź�@ã{����l��M���m��υ������ev���~u;P@£^S(Qq's&`������4���#�F��]�����p��C7�"]�$��ϻ��3ز�lh[��ӌL�\���Z%~B���[���d0�(͛>0���'R��b�CbYx�;2I�$U��`g�6nO^�x�-%� ��R�r8C� aLŪ鰽H㉬�y� \>�/���e-w3�v*7e]����iEV�Ǐ��;����2��{o��Z7r�O/���'���E���H+!D�qqQ���9�=z�lW�Z�.]�y@]Qe��,e�S0Eܥ94h���������b{��Xp`�^�Z{����D��N��z<Ib��[��brҋ�:nT�F�{z��^Nyu��WX����IJx�X�/�V�M��ʁ	��χ(֋x�'o�3�C+�"8�.���c�bF6f|�f�؜N_:�9��=��w��t_�:��=� �Wn$=C!��<��Vc��pk�<em0�����S�A`a��V-�)�7T�w<.���\1S��,p��w�֤�R�ඡR�Hn��N|�H���Հ+4C} q���șᘻiR�L�G�%���Vu���xѻ��XRBV嘇�
�e���#h5�8��+e��et%ʝrZ	�H7� :1�B�^�p��X3lӽ�q��~��Sғ��,�u�p��k_٬�+�X������S�|=���q����i��,��y�s$���8��D�Wۮaw��� }>~E(6C�|�5����>�ue#�`���%��bs��鎺2` "�!ڄ�ya��0~t�K�;��\@u����?f���\`�i���A�t��vj~?��w��U�m3=���MUX(!,i?�;�Ґ���B=��ă���ƿ�lE������9�������ڞF�r8���T�~xm#]9���xƄN�:��|�Lx�Y�A��		���[�
�=K�"�kR����k|[z1.�8��I�qAI>�^��N>QG�����~��<�`®J�1`j&�X0zۨ�#)�I����F�8=8�Ҋ�����)g�W@�����Y��t^�[>DЈ�d�u��%i:Q���vzI�ߤe��Bٲk�\�XW�s�^� 9!J�k���\
M&�oY2�66b���IWpr�	h�,������ l���w�
Y���(KF>
��[��&�愋m�Y? ����u~�������O|��W��$����������]�{��<z��۞�6���J�&G�[/��5�����(�F��P��b�哼w4����w�t���'��p�ψ�N$��3=��F_fA	w��U�"4�5�˾�4����kng~�J	,aM�ʚd��X�耇�0yD�&�)GXUh�i��5�_�e���$:^���dۨ[�j��i�%���ӟ�QCQ��vw�$�hܨ� 8L�|2�����}�� Q���9���A�ϯj��zF�΋�w�crW�L��GA�i�Up-]�X�Cm������Ï��Et7W��	���4�.�/-���4b/m�B`x��`�OHEQ.��g�6�r�yD�|bJ3����Emv���:�H ;ʼR2n�j7W!Ng^�j�:��vw_z,�?�����s����V��Uj>�7|r:�u���_?xol�o�|Z;�z�3E���ob�^T�����J\�w�|���JKܙ����
�{eR6MA"�c�@��uA42.]�b2^�sY�sC-%K��A��Ϣa��"Vv?Y�*�WMN�t�<=�R�b��P(�1,��]fd���P����X��H����������w#r��u��k���V�d'ݧ�.D����E�h)ִ�������'�D2��Xm�q�s�}Y	�>���k�N����@fr�a�ȿ,���!/�{���c��<�\�{FDc�b�ZB �dx9Bp:qDh���%��:c����w49� B����p��X��SE�hɐ����̳ך��?��&���˦r�3�X���OC�(u���V��YO��M��Ey�9V"���=�ݫ��SM��F�!�J_ �u���zs��O����թ9���]�ƠJ�6�Kk2_��^t�yDM��b�Ú�*����ށ!�1��ǣdW�`:�K�bw��!S)��d|��Z54���U%�"ܪ��xNj7N%;U�b b���L�e7)�� b�1p��-z8�Nն���>.8�!�\*'�r��(,-�i�'!tB�LD!�1NK�����ڕ��	?w~�^Qp���Z/ע�{���C���c��Ze}�L\��w75q���Ҝ�ӇҦm蒟�ޠme�i.w�@F� �;����dFk%&��?��5��#���PQ�-��<ۊ?��~��`�K ��	�@?�`�.�7=Td���.�Ŧ�w�Q�S�z�"7�(�oʵ�T�݈�,�_�H�"<�H�,Q��v��(�G�Y���*Z� �|�[ѯp�D`��X'[��n���:n�#����b��iN�F����W�79ĚN���,%�u��9�s���=N6p�wvp7���	ݕ��&4���8VB�-��ϣd3b1j�KJ�N��B�$�~�������~W�aV�t�7H%v�a*���N��w������� <4�R!����V�6n�}��X�$6���83U9��4LԱ؝�ٷ���Lu��9z�*0����ɮ�e��Ank���Pk"����*�wI���T�Se�R���j��=_�0�WܶrZ	��]����!�Sd�ο4�q�߽�NO'5�H��/u���,ꠚq�����HU�ٙ��,���<y�j���d�n��0�q��^\����ޒ��td��S� ��W���=[K���B��}�ޓ���Ԏ��]�<����5�L)E�b-�]�Gz���m�8�X�W���.�leL1�SB=�`�7��,�l�v���Ip�U�i,l�>TOn��B�O�m�h�1U�/eB~
�JW��D%�u�_,u��#2i��1����6�*�J/?��!�����@��qu^m)ȉ������E�E$CX:jl�q¾���W�\�'/vO��s�y�wJ7��ky!�$�(�2Өj�*E������c�O�襃V-�F� e���!��A�Xռ/��&/)2�^��O�o��z���]HwD�g�p&�|)�Ayu�����df�"�0z�hr�U]��!���~GU��H ����>�;�(c�dq�GR ��χ�s���ꁚR����ڔ�>\�gP�p�-ʣt��
��=�ES����b�[x���K���~3��3X�_�����7'�&����K0Za	S�X��58t1w,_�Û.��N�cy2|$�[Z�w-#��{p��v��R�0 �۾�ٻL����J�֕R��	,ID �:�7"�B��ux��9�2]�$=+>��������b c��JM&C>�!QU�:ZXT`f��JA��U);����̌c�F�ڣ7���K\�<�3�Bz=��Aj!������{7��[��$��#~:m���ޡ���j�g�Rʙt��>��2񺞠B�)$q;�uۻ��	r�=e�*i�uPY��G��l�������ޯ�dN�W�[܌n�q'�DkvorN���J"��ם��t��9χ�!Xs�b���=ό�z��G b4#t�tk�)\)+�q���<F.;��� >9���,�Ώ̠;���z
0�n��K�%ꉥg[�D��5u��V6�'�tx3�P��yM��>�̌d���bdwp�7�(|��	ts���1�Y��D��f���6$�!�!�,/�r�S��}���4�|���u��Ǿ[q8�E�ւ$��# 1� `HS(mV�1"nJ���F�y��jN9 ᙘ1AS�'� F�N,�*����v�Dxqf'�o�ݤ���N�w�ȑ(Í�����	����S;w�jƈ������Mqx��ԤMN`t�LX�Z�Ҷ����p� �o+?��� �?b�����^(�3Z6]`;~��p�m���w(s�|�:���h����xl��-v�D�$�n���rAk5���S�`�l��?@  �u�9 2e�[��=ػ�57��}G�2L��v�ò#Q{:�cW�C��
u;{~ɕ6Ч�~�Ux͝�!�X��f�};'�y��[���sJ�l~-eɑ��FG���Y�Ra�m=��� G��ɨ�ˁ��o;,����������캅��޼<�/���1g��v����j��ItQ�<�q�CǗ����~�;oZ�U�,yS�W��������_ͼGؼ\~� ���Un^��_D�&�!��R7�J���>��lh���X�j	�m�6��
,l��\i4X=��"ޢI��
���Q$�b�����ރ�`@!!�7;�h���U<#�AL���<Ԅ�q�����wwu����PM�H�����Ȼ$�w'l���~���BO=V�ɩ�-�����8@ v�?����o�cJ�[���� ��	9����g��?������WGe���;ĸ�*P��F��Ep�kh�g�JJޱ��ti���W6�䈶�� �Q\� �#+9�%�T�;`#�=>v#�a�� �I�l�%P�B�&�:��`8�u�*3�1�:`�e�U(h>��c
߸�ƃQ���ڍ�����e.TU��ÚJ'�=�1���#0��Y8	��_�����L�1�������$�@i��AN�Eq����!�*��0#KO���ʹ.�0)� ����Y9 �9.�P��r�oɏ����i��-��g�
���0�ʳ��{���;\
�@�l��>W��}w�@D�x�>��M���.\�7��͑�ȇu�|3uٷ 
�P�_˭d�?%>�l+��(��C���d^4ɀ:�X�M)nza�X������D�HS�NC��{a�	v*V�'5=1l�p�nh�(�]x�/TO���9�r��E�D�
�&�u�t��ɳ�`Tw����L��v2z:T�$�L�0�bi<��M��?��OD�.��z�)C�ʹ<I�A�G���xGҿ7��B{*^�t2f�T�Ug}r�67��z�!�4��5�-m�(7������yX�<�5]?�67�u�ۙB�q���0��rx��
��-!­AC�<�z��&/��9��[���q������'��.7�
z�[[OU����PM#��JI�~'�(�`��4�WI��j�/U�>�EzS�$�ݸ��$�)�D?6o!�"C#	�`[��@� >���o�V�E�o��d:x^�j�<��:6�񲚯zU��hM��Y���8�ʷ����}Y�򴮰B���i���'Ԭ>�?�$��P+��aۣ�x&_���Q��0�d��C����)�����9ǵ�Æ��`ս��Ȅ��ܾ3 u�:�	J▰Y�O%��)G�}������D�1�\��`����p1vpG���Y�)�.�'s�.��
�T^$i�m7�>����(�������eB��0�Q/�̀�R���5��Yq��1<Ը�SoT�#���l���3�󯧐&��#�V���2~��0�~5po�M�S��h��6bc���}��s�Z��=vxJ��/P=~�ir�C���Y�^!w/����9L��g��B�����Z>���FK-���c���,L�cI���߭r��{/ܚ t���q��X{b��g��
�)���f��g�m��O�F\��8yG���]��!����T@�?�
�Eh��	����q�}o��c=ı��J�J�[���u�:*!�����@�����L)��D�l�T{٩��T!:V�&�p��E�'`E�^8�3���c
k�b>�wYL�n��k��R�ߩ�*
�H��v�|].�c�����1C6w,�:�7��m�8��^����-����ք����l������I� ��u`�����0-�d�Lu��Ao} �O�V�񶬍�� .1ZYh,�N����t'�Gɵ��W��q�\�E%����������� ��):�\�5գ��/�^�v����-.%�%b+��޳�n'�W*�?�-
������KL+|��l��Noy(	Lk�Qm]�����A�7���Hژ�I����9Fn�U�J�M�ipL�^-:�1E2��Ȏ�G�?�߿[!�HmjYO�k����[��~<5d:��<�-K�����&06+�?��-��@��e�[���4��9����9س��l��N[+|�WX�r��%M��r!�R!��SR�kp�L��uW޽����߰���i�	���9��F�w��m�N�]ܩ���:��ǻ�0�|��?�w*`E_N��1�O|��2�!�جU�3��͙.X��%oq�,P����x���*���Q�h��J4�_�i���
�Cui��b��� �ml|6��D�MI��T�AtrYev��Σ��0m��� n���Pܕ�X�G���dt�Ր��o�D|�=��L���_-!=���̿�[e��P���B�~��}mZ�V-7�ObǮSiR�	���q��b"��/�@��x�$���e�5�<�0�yV[��y?P��C��ê<]�?�{ԃw9��Y�J�i�Z����M^2�E�b��=�1�v�V���јz��=s lD�`�Zr�:@ok���ZF�`g�&u�,g�+,\j��������bvV\c�Ϣ>�[e�|�/ʙ��������J�1Yp�bvqz�歡 ��e�T�+I�m^fЩ�7�W�Q�3�Bd���>�Fӵ-�u'Ntz��׉�5������`���`"萁ݏ��'�5�>#��Vb�Տ�3s�z�9X�W/c�!��O���L*���!ُ�i����'��'�-�ak���^A3$QQ��ξ�]�w��Fs�.@�sd+s3�Vp����Z�TA@�P���.0f�K�ҿlP~�_P�+=�>�y3��	���E�6ґ'f��R�^ ��b0CE������L�9h����C�>]�Y2�i��'�\��;��)�R���7浛f�;�Q���RQ?��T���|���7�:Q*
ph U�,@!Y;���,4<�܅<���*�x��}Ye�P�pނ�ڱ�h�ޓr�&s�M���T�<����&1؃�-xe7;���aj����s\d��x&Ėvۃک/q�IP�*$[,�kPT�H�ED�i�uh�Q�H���VY2
�U"i3�b=~=�ݚ���0|�!h�ߜp�{���?��p�Xn1_|��ù�,�My��bV߃���>A�����ը\�˓)#+��3w�h�fH�̭{��1Z}�P��0T��|M����5h6Ĝ��s9�D�p���X�Nq�Z�ډִAQ�]NX�L�����^�(8��G��\G��������4���bpyf�,9D�s����d��F�*�+�����_��o[$��[��12*�GS����|�*E󸿊�3��B�+,�Z%���&C|�ߥ\��&��#�nU_����H
��
�� ���X`}�TWg'~K*zo/�Zi�������;hKg�u�%(�a���C��Sn�ز�N�a�7�����-�3l�Kz�Q�a��r�vi-��L8ǜ_hv��,�m.uIx���~�������C�O3����	|.�pk��Io�6ċ��}*��
�t!~:����y�p2�,�� ��~u��zC� xЅO�XNcL��{�I4�D��ʹ������ ��Ć:&I�HY�)]���境P��\�����_<��+�q�u?�x-U��ϯ�a�}���v�M�_���ZI]EEJ�[B4��=�Y�cSL$Wv���]F��ƚTF�B�wn���NDAJ,A���f-��cw%�Ί����}�8+}�*d�#�l�c���X����n`�&gx S�8_��h�b�^o����eMU0/{i�fA�f�S}~�4@��Za2a�<5n΅��Gv4��i
e���LU7�~����tSO�<��ٱ��#9�3j�N�'��Tƣ��AI4����=%�j��k��j�����z��,
����2��x!P[�#�����m )��S�U�ڰz�>���}/�S�E��]rF��6u����%�Ա3�d+KPL���g�����'��oQQ� ��T]%0f�ҧUl%�r����
�sy�rn'�*
�Lܬ����w��r`e6�A$- γK���pT#��Y4H����L>���_��]a��"�K����O�>KMzZp{$��p2����l��:\�I�^��f��M��L�բ昨���F��� c����4H_�~<*{�*~w�#.���we�4�RȚ���̝A�M�Ƭ��R��O��(���Ԓ���i1�Ϙ���b�N��^<�UAc�)����q�ٛ���r�]�=}@q����3��F�&�]В������%�0�C
K��z5����A�6(������Cn�b�$��V�
���4���&XC �ęܢ�c���Gw���5���l�����w]������r>���7�7P��ޜ��\�!�W�$�¶	&����H�>�8 �2��)�^_ǡ�6��"}M�`�$�B�eJ�4��#H�D�߁ַ� �����\��g� $��t�Rnc�d��$
Ӽ�a*&�i������d�"��#�:C�`��zdnީ�r@7Eg��)b�]��-��^����W���[��aU4��C���� ��u��'L)�l���\6�����q8��d���#�/r0���8o�����a֋Hl�^2y٠ɹ��;�DΓS�J�\u�ʵZ�@_�e y��BQ���C[P�-�ENuk�HZ�Wn`//V94WA?s�n��+D�B=�����4y�6 �;D25����9a�3�T<������7���`�[�[#��-���'B�p\���a�L��s�����KW���מd���+ Q�5�Lm����.��L+l��B��,��_�E�uLk߹,&?H`v���h�� z"TF7\����U�����\�M�<D���L�w�d��\��Py��nѾ5
ZJ����>~�״F��|99�L��!�Ǹ�o�n��?ʗN�S��N�s÷�P���3��^�=�8����q��ޭ3�SӄP�̵�8�ϵ:6�|����7=�O�I�44�K4Ў�N�o� V�������*�TSK�ق"X"��	���kTK�k���uƔ��}-�[D�������?�S.L�3�i���s�O�q_�3>1K%�D��]!Ҟ��C�����@�GM�c�Q"�b��̨Y�#MQ�2[<srj���9���O#�ͮ�J�ٜ�~������ȏ�*$��Bb�-��]
Ɍ�g�}���m$B"SIX��k�zSj�۷��q��0���(��)����9t؋q=�9�`ߙ|��<;�`�>�KLX|M�^ل��*{S�G}욳��t�_Wҥ�gQV���ߪ���֍��o(����P��EF�u�0�q$�8� 2������t�sJu@��*E)�:�t�Z��.��������2L �D����l=F�^e���g�j���CmD�G����7�]�����Ƀ�?V÷���+�]�Ok���c��%�Ҁ%<f+"U����O� �U	B�0BXL����o���Ehrb_���<y�\<��0�v����{�I�e��t��~��F;�!�*e����k�ܯ6^�8�'.�]����DC�cޗp�_�諶�WETn��*���*7�{��g�1|��omǖ���}��;gfٔ��kܨ
KW���נ��C�������� p����s?�ig�2�����Ҹ�����������HrR� ��p���8*�,�
��D�@'�FkG�s�n)���4t�y�G*	����d����� �%#ٷn�('~����io}%�(�EP
9^xщ<0���vl��th���	�4u܅S�뿕t9���8��7�Pː��r�g���@AR>_�c�4E�u3).��������1鐮�^�b��a/����8[u��N-�b?�
&��W�-R�*j�"$�z�9'�I%����V&��xi����m
E����)��r�-�Gr����|I;[�F�V�w���\�b� �2��	�#��q����LK��0/�W)=������)a��.��6M<�F1�Y�p�;j��[g'���90��9��Z*} u-$0Aַ
!����`�'�8E�2©��Twi�ZkQ��ű�@Q�Z-����Mvd�f<|���D�V��V�0��h��Pv�l�I�*<q(&43��=+��O��Nc�U	���Nvc"(�;���M6�y�s��4^ء�����o�O���)F�&	�F���G�%4 ���:S���J��Lgq%���
�A̡��PK?���֟LH�_('����O>�Ԏ�BM�|$j�
.O&�g�֪uf\�� 4yy�ϽgT�ؘ�RZS�e�dK��hd���b�O3�7b$ϑ��
wB^���7J��Y����ȷdIL�y�O\Ō��&4N�|3�3/���dê���5�,�}�Y�,�W�A������gdca�WF��ȃV�]��(���n������+ˢ� �m�}p
��Y4��;���-Z���rʦ�H>?1��[?a�ϥ\#��qc��U��|�����ݫ ����Y��;���_�WrP���1(�%0��?t�_|�Yh���xJ�@$5X��֟kqOi8�$��Xp��I	nX���V���n��y�-�pK��c�ʏ�2X����d��b�}ճ7M���Z�֓����x��`��Gs_M��=%�敫�_�(��L��i�'~�}{�op0��ܜ� �w��Q���e���mt�f;v���L�GOW��֟z�T�J�p��SW�0�����+
=�qC����a6�O��:s�������?���x�x��A���h�Z)�-up�f��8]¹�mZ���7���v�CY+��#�������� ��/c�s�CT����j�u��
@l31�%�i�dA�C�@�1��%N�UJ2Y&� S�������i������m}�RT��sЋ2���Fqkm�D6�A�*�DY
�f��<2�������WHv����l:Dc|�7fT[�nP���1�� >�0<�)0X���H�fe�[Cc<�}��6f�f��"W&����D�C�~M�#[�	�:�-J�Br".���v[�t��Akq�B�v�DmJ*������ܛ�:��C �鯍䇋-K��<��pM��2θ]�冀Z�_�s{0<�aXMqO$Y��wA�P�p�W���ѫ��J�oV1�,h]�7r9����Vj��U��kg�,m�^[3��_��^h���8^XT���u�+��8`	����c�}Z��Tj�I�ϼ�3�H�����!�|t�����b.�dI=ĝ�n9�������g.�`T����e���FT��H������z7C�B�5a�̳�o�8/~
rl�#���[7ʹ��E�28�"/�/��Aw=Z׆�ݳǗ��.�Yg�_��b�Y����MgX/c�>T����{Gr�v�1��i��$ ��5��ǂNJ��]_j�+ȭ~��̕�8	Z�N~��_�x]�g�Ms���������ڇ`�[/%3�`/hlY�7���=p.��&�@�+2Ĉͭ�plo��Q��� ��t�i��8ugz��yz*M�:��R��]��#J�����7^�W<;P���z�yX��N��h"�"4��~N���H�j���Ly�HT�� ��M(���{T��]lɗ���*g��@���4�DW�a+�#�����]� �<6}�/���pS|:c�#���|�C�����C=�|�N=%�|�׀���T���b��.#$�"�#p�����g8dtЏ��@�`��	�;���x;�W��z�|���T|Spt��o��^72?�m���� ��L&��%v��ɼ�6�3�ʘ�C��$�
��<��� Ғ�$��V��jk�<�_����5KwC��-=��<<2��� �#�Ty���_XgR�ܵ ���N�_q7��Hhk�D9��KS�T�B+���"��ö��Q>��{&��lj�a����(B��pQ����Z
'���yd;�%nN��͝!�ŭ�6���<"��we�Z/��3"o���褙7&"��+�&�LHA��rH�z$�bP�� _6�ȑ��h���oF+�S����L�+�<��@D��u]|��7G�2��;i���	q�'̻��i�N���]�~�����/�G�iIv��S�O���"�Cc1�
9M�x�^b��]6Y?a9P���v<|���1�_ĺ*�C�З\�h��!A�x�ȵ$����yN�~}�����x�x���y�Љ9�Pò+���?���+���pS����L,�(�x�
M"mh�g&:S:L�?͂��r��/L*ь]�P,y�ط�l��0Z�:����$�(�������4\B?!�tM�ݔ�2����7[��(�μ��+e)@�Y+��i�4��^H��B�OI
�f�x*Ɗ;�/Ol�9>{;���4���,����+���4U0�'0���0��7L r
��<��	��Y�ʑ�7�"R��	Sl�j�o+��y����0������v���c�ΤT�c�ԡ9Ѧ�hz%~fYX��� /�S�������%�N��!�C���'��^{@�W�fh���5���<��7�DK$���9:2׎��})�qt���
^>��)��`.9��T��0;;}���Sm:� ٭�C�P�;lجoteL�G.��>܃��X4��O>���k]�{O y�/�?��#�;��z9K���Vm!��J<�%���� ��0C�n���u螫kɤ��h�����}��W��Vh�(�D�K�_�����ւ)��|Sh2����H�;��1�Y�D���%F.Yܪn*�z|���8��.�*��я��?9���n�IK���}D��|�/�U�:#)m�e����e�1Ny+�>�d�L�����kT�����&�P���ڻ���-c�ä��2'Q8�n�E¬��~���V��&��>����	h��f�l�9*��E Z!7s��[)g4ʹ�@=��@�,�t:��8U<$�e�� a߶������=�Ɍ��"暿��@	�P��T��m]�A�]B�!-��n��ȇM�iKE5�|�5�"g� 3�-�m�5�_~"�6CL���9�C� ��T������7B"}D4��Í�[�Zc�o�۱�+����yRTw ��	����ʟ3������7tL{���j� ��~�ei��W`}��D	:h-¢<��<�$$q�M�E�.���>g���fB��8�j�z�k׀?	��LO��͝ @*wLw��l_wjH�]r��C��i9ޓj���{�z1C� ���;��A2�e]OG���@�ڗ�C��R��vC�V��x����q<�ӳ�D��W˝���C�	����դ&c�$'0~�'�L�jz��	c�TN�� B���,5m��gtP�pp��6��Y�)�k�G	�m �}*�@��W��g��`!S��ț�koX韨g�z�"4�1uث��rş�TD�*�<˧���{riC�7NE����<(϶�K����L�(d�.��4+�exy#|a�����<�A����ᕡ_��׍��V~�?8[��$��&�x/i���N��O��AyVUX�aB(\?d-�z@A2�<ԧ�r����r��U���^\�7���l���W�BN�n�F!���a��Ÿ��o�Qm�`dM���r	���?b0|{NѽĲ�~�3[ǍS��ް�=���-��r1�|��z���KBV����#�뭒�����zG��O��>��''b��nK)%�P9��b;�xg��Ӧ���6Y�
�Ȼ�Y�LD���ԏ�ωcg~��{"����-z�6B��Nŭq�d���_����hsM���f�tnO�'#�}y(d÷�Nu�b	o׮�i�kE��|�T���pEB�������ή��'N%�O��?��N��b&�,QD`̥W�Ü���E}J���2P�O\*[]�0͢6�K�J�3X�"�RC�.{�XHz�+����CՉ�q�C�5�Hm�޻1<�1��,g�3A��8� �ι�:���0O��'+�ޡ��D�Y���k'l|Q���c��'*��]$h�{j[����b���C{}.��Kvn�_%�ˣG���!���L��M��|�`���i]�}lc�#��]P�ل�c̄����������s���]���V�B�D�ӥ�����Ѷ��g,)֑HxE,�&cl��ר��Gs�#zhʯ����b@!��(�R>�9\Rq���ɕAgw^��5L��e!B�Ƹ�����ǯz������R���p�w��n:Ϧ&`G�>��ĸ�1��K�,�_ �$�b��L�*ň�a��8p��� �x���1� �g�lU�?�tA1Q8�Mw`4u@R�
���1�U �w�Qp?h��C�����rqx�Q��Bi�<ra���k�DJ����������q%�ׄ~:��g��ux,r����p���5�b30=?��aZmƺP(&i��#>�s4����D-6����	j�!,ŭn�{�0��-�|�2ˈ�oY~ei����B8�Wo�>�4��l8 ({	��C����fI�;��S�D�7kY�Ve����#���t@q5 �K�tp�L�Nx^0��!Q�OnP�շ��(V���X�����|�.��Z�cE�Q'�'wae���k�>�i"�+�5B������o������@������jh���b�2�)>ШK��r�R롩����љ�b&j�W�23F���G��ź����=T�x�C.���Z�i�;�����.�[+�+9Xex�:��������� b�φ�2���F�
r�ي� �nWHh<�2�Q֍����_�ը�\u���N ���W��N!������f�&p�j{��u����dT'��(�qGE�2Խ�1pVM;�ʝ�e����C���CE�r���_u]J�4�g�;=gj� �����H�N�8�RR"�D�X�2:�)�����>� /��v>l���m�T�\`R-�C<��{�"��c�bR�:&j�!-	�:ъ��F^����Y�7�.W�):�i�[�L1o~!������'��IՖ%�&d�*�b�rCŉ���uq��m��Ui�l��7����>{��j(LNT�5ݕ��<���t�.�)SG���/������k-�s	�F�^�$�5r*i*ᦱ����d4Y�g$R��}2-^��Jj3�Ens	!Q�����m�%'����ܿ4uW�K�H��[�mh�ӣ�ʾ|����lT۰O��NB瓉���.9`
��J{�����V v.����b��]�#G����./�u�VL{��"�M�
ի�1!15�Gy��z��|Ƣ� ���q����� �9Q�tGo����J{U�#� A�d�9�q.�8�sO�Jܮv�:�E�\%�]�}s5�KXl.t-�p�������@��Ϊ�������9ӭ�Xh��_ �V��D�n�:+1�X=K����1e�j�E���NQ�����ϳ>���"`�p�G��|�Gq�R�� 1|��*������ꡗ5���I������cv��\ڧ���i�e.�S��"ٖQKN���!mq�I=
�uZ�KVUq?���-�
���͡���}*%Z\=�8���^(��T��t�+���3A�����hA1����!j���������8����E��h�tb���{������O/�k�cB��������Ė����{��'��oT�#�S�Fb�-�l�\�AS��y���O"���dRjd>��_� =º&� ���#���HB�o�C�������D�LI
�:1~p�霴UxA&�[�� ���y�wgdݢ0���>e��!]Զ~����Q�xhwc��YW�mƸP�}�r8I>ki��H�[n�0�g���N0���G��CB}_vx0L�#�ZuGΞ.��dL5�����7��	�>��'2�[\l.ms�D���&N�ӫG�"�wm��9A>:�h�O<uf���u�1�c���eQ��xHn��F��Ga�AvA��;L\�̈́V��`��|.�>���m���i?xM�	��|nŬك?WW�����6oR�Ю�� F{���/v���}�|�^��}�bM4�K%���<DT����o�<�HY��1������~P�v����ST�t�p�}�c��VŮ(��!��[!Jt
$y�N3�����+e��q�DV(n���W�~W�+�<����q��K��Q/O!�L���Mz�m�sy�tC��f<Ȕjag��euRא����h*ۿ�tl%������6�ꅩK����β��i�+����L�Yra?˧��o�� ��!=�+����YL¥:e�9{��ۆy�Ｋ�r�5�� �+fHs-&�vb,��!!�Υ�lMm��;F�α��C��wQ�9;�דt����yj(�N�O��,h ��X�&C�x���%�AQ���-��S�m�K�8��E��Bs�zh��t��[?X�S�K���w���<?^'�ZH��	6�/�Ȅ�
D��!�E��E��'����n>����� A+>m<�k� 7o��z��j7 l,ߠ�~���W���O#��z�D��{FV.�KN�·5M۟a�4�3^K�?,�s[ܨ��Û�kL}#P���>�U����1'��64�#	�B�b�;݂�9\�^�����9z�W���=�֯�c��`s���g5�%%H��4HW�2!K3�<�����zh�����=^n�J���s@x�b�� ����j�"kFy���z��{��b�l�	������C'�CNJz6�i�`�����������~0I���g�M� �����,{�i����5��y���,��{.�J�Rt��tr��D�ݢ;�"��,��\@�������o�s�o�H�'z�Ѐ�(r��U{��Al?���%�<�"y�;��+,ϰ�ŻXq�� ���dߟ�^zW�6LX^�s3ձ��g�X(:H�-�֡����|m#�A@<*�S�^�8�ڡ�s������Q{N�]��.Mh�B�;g�I�[Z0���%��Ejt�����[g�(m���w;��MU��+�NgS:�6Kk�R�Ȃ��@�&N��'{���IW��[s�b*�@���u��2������G g�g>�p9�`v&ϋq��F��z��#��7a$�3"(ŭ��c����e��[�:�����A.��f��w��RELn�u�M5#Y�И�`"��$��E]Q�/��|"�m.Ppj�D���r.{BD�� ���=�e���תت(i]��*�rfR�o�,�'�d⏹S.����ö$�aѩ�z�r�ۆ����5�G�R�/��C�=	ІX��t�� ��վT��k�~����=���b6����y���J�X#�_�H���)k��Ɖ$2�)%��J��馎�t�w��U�.o#��+{�:���U��T�����rP�o��y�������Q��W��wx��I�ܜ4���3`���W@�Zkn
�'޻�7������^��D_π�˃x}�(��������z����6��ߜ��*K3x�7��
�E�p甖ڝ��q����i�H#��)�������3f��&�֌�0��k�7���2��ͨm-~/s;;'{�2I=����W��HġChD�������q��A\�kO�̛,��/j_F-�A��[�������}�j
Qrke��0$���ĥLd���w��D���[
AI�y��<��f�>)���>`C�^#�����p�F��oI*&L��ML��j�6���aQ/���S�!����s�^J5Tv���2o$&v>��v���ܐh���
ya��Un����:P�[�<�D�� ��f�U���BS��&�+~j�̉�S�� ���y�;��Z%��tAWa]�N����wG;�������o�+�]LÙ�>
�	�҂��S�����ײ�LJ�b"#���>P�)���I[s�'�pچ�o8�~]=���R����:B�>S9�_�rևT�Y�g��r�����G��<��ܾ�������^���U-��w������qK�x�p��C��[��ޓ���"�q[B:�H���vC��v�a/,�Ĭj|g�D���[����Yϑ�R�5�`$���PC�>��-�+;��׵���hΥG�r����d�i��H�Nv&o�`l^ħ���w<!�W3ܮ��}��)KM#	�*�N��KF�7{�w�U�ˠ̷.������Kzۍ[��Ǖ]n�1�bњ�1kɛ �t*9�nB�6�eՎ1��Qd�Ol|����a&�-���25F�v�=���ܮfg��5 �]��n�|K�L�G�*��@���ݠ`\2h5�����䏈PBl�������5l)JN#�}|o8����.���S���`R��>r��ɥ/2ELxÃ��G�d��ߵk�����r����ڀ�-l�Ю)%�3�e�,��܈:;_���@\K�"��`��}����r���%�_�/����%8*���a̕S�L�S�վ9�/��|��ȱ�6/F$�9�*qpL�[����ظ��@S�[t����~��CȬ��?�
�a�|�R!؜9f�C.�nA~�4ϭΚ�0�^���W<��K5$�^�_#��8a>^�����9�O�Va���>�q3�h�<���Hi�L���,2�T�*|��M��p�����>'#�`���'$2�]MR
�*Z�$x8������&X�uH��L���r#/wl���hs�)��U�cTp�o��K2�Z���@����N*Bڞ<EQk����lg��^�q!��RF���v�}�ż�.&�.�I�;۲�'�)�%ʭ���`�.v�k�.�^�͢<ާ�����:�צ�Х[��Ү��i:/�A�;KY���ot�\��|C�؄��iH�#�S.�����9"�syf�W&y���4@wzLcw��%���d}&��J�)6���~��u- ��Ǭ��`�+��;}z���Z��P��^���FD�j�`i�oO���Q4ӦHS���e�Ņy�r�l;�ܧi���74�����9S�#��Awu.R�d�p�M)���8�e��$\+�k��	yQ6�@p��/e��Ы[�ō����I!�#�2N4����R`) bƘ/{K.�vy���a�:ƹ­�n���-��T3�wّ[���E+ksܕ߽J���DZ6̫'�[�I��-��Ìp�ͣ��ZJ.�6�F��1u�u�kk��e�*B3A��_�"U���\�n�Q��K�4
������f����py����"	����Q�oޗ����O{r�WFP�O}���ADK�wq��#���i�g5��?��`�ճ�n��BǼdT���a,"����F3'�y��W��}��ٿ���]�_aDK-	5%��Ϩ$���H�\8����4�+���=������@n���}��Η�(�x����YVj��XK��;$ڭ�wTvg,����!47�R�qm��6^@(
F�G����ԙ�� �'�}�&Q����Λ�2$�m��p�q���Kdm0� H�{�< ��������%z�X�yrd߉�(�䲬����7B�z�z�U%g��H��%�k�M��cT ҆/)�������#��� ���ޱo����E���~jm6�Y�G�L,x���Wծ V����ŢSw�M�K����*�����A$]��9�����bD�A��b�HC��K�A�l��F6���9����� �j0���(�`6�����ũx�6SFJ���}Ɗu@%B��퟊�1���,F3��c�R�'�b5˝���C����;��EjS%�h;~�&U/�o~�qX�5�
M�5�K�)]C2�MG�xd �A�D��*>�Ϙ]\��@(�=}�H�z�'��UIw 醋1ZF�q@=j��ء�����5w��ɏ���@4.�Z����L���di�x�$��;����T��S긗˧�~)�q�uU	�R5�4�o�M��*��lx񄸵Bu����Kby�b􇳵�b9�P3v�-�ϒ(�޳�>�� �\x&c��+�܁� ̊�N�1\�b�@�[��A���~9{���p�;��i��´�NTS`|�
�n��u���u+��L��K��{z6$AcJ�YK����.n�ܪuJ  @�O��Εo��eNF�{W��KR�X��ߎ���Jf�
nȇ�f�����쨔ʯ<�
{M+����Kf�U��Imρ�M�#76���jo7�;��
������{Ͼ��|3'�]dɖ���]6vk�L�z*���Z�cN�S~(�̑��[��Y_�c��)���@�9�am��T�)sff� �f'���KZ�����_�UV����}�sx�MS��r�~?��6c� 1������c]lYN7�����R����eK�lؿ���j��Y)�$^}$Y0߉xѪm�e�4��Z��t_�<�^w��S��̞f��O]��	���8���
�ڶr�󒓀��Ds��U0���e�=ǌB����'t�V$��}Oo��V��F��N�K�[�<ӷO�"~�t$��������L�J�G
:c\�_�7��,c�PP˓(�sۿ-\�S8:�x7�R bߜ�_�7q#�(��*fM�7�|�\Æa_��2{/�z)�K3�
�	.2lt!v�r
��5&چ(����Ell�C��*�ùj�ly����쿅!�3w���C�gw˲�;�		���?�y�x,� ^��t���͞�l�;s���'��$���;��G)9m�Єq����G��9�^�uP#XD�t��=�a���>!	*F�S\M\�h�km���]��l;fBg�y��6���l��
����H�� ��C)n�.�5+z��$B���zL��	~x�]h2$z�v�`�7I�dX���� od�%y?�X4��LW�J(ꖍ�K�?��z5	�u����`laBB�N�d�b3�ӞF��T枊��l��z]�"M|��aPC����!�����.�(S��ꦊH�Hrұ�c�E��uA/g�u�O�J�5j��JP��r/�hH��v��s&��9���q� �Յ�3�Q�i�ѦET���/5H�ҔA�A6������u���E�#5�Z�Ѹ�4�\��S��0D�K�/��Z&jYe�ɑ�E"þ��m�N�יڳ�7�S����~�pHY7Ͻ{�Y�f�%�o��-�dk]�5�A��+N�L�w�e��݇Y����~�=f��6@N��7F����������������׼9�ٞg��b{y�θ�l�*ëw�N��[�)�d��]�ϗ���8����Ƥ"̇���a+�׸�(�٪�"����1>�!��M/Zⵌ�Kƚ�ٽ�&���_42��&�+�Z�8a�M�IfgYY �����?~��z돀GR��M4�\�?�j	��P��3�a�8yԅ�l!UB+�Al��]2{����
?�,�bA�x�-����+�*Xd@��z�W0q�;��<�-�h*N�����S'O�s��S-b3E�A��*�ٕ��\6�]����=#п��`.�1h��ii%�,�?�5�P���X�>���I���h��� ��E_���\9Sߪ�,M��pwjy���P��`?����(��#�EEo��5ZD��y>�
#�!*,����ZP��?�?��ī��o{k�td�t<>���]�#�y�0�,: �dϠ�&��yx�;=��;�5����8��b�s�Ȁqkܤ!n�P!���dR�s�����cZ�p88$D�0uݾ[����2�����[O/��KXR�+y�/f�����(�u�S�9A<%YU0��|��uY����C��<���i�8-0�c�����$tk4:�����0PX�b#}�ƞ.�GФ�n�N@��ws����+z�姐� �&S��`̲?@�h+"����3�����]�{Yc@��x�D�/!���l���G��\&��J�r�&J�k
YZ[t��4c@Ԍ-�`oU��`wQ��#f��V���*P�Znd$��AN���*#g�-)2!&넽M$�n����{L��&g�J�-�]D�ZSY���ga��#�߱�`%�5I%ā�2.���p���-F������r>����g��s&d\U�+b<TpG�z��73b�I]�0/l�MV��F�����)��a�K��E17vU�W�4���#�g�H��Ag��~���U1���xU�m�l�R";�@��"H�m�3�.Ї��[�R_��j�
�8���Dg#���SP�㐞�]��\I���}��H����K�')r���3��� ��)�1>�xˌ�1N����s{8�I "��T@�h�^��� �h�����
��My�%	�{�{�љ���j�v^ا��Ru: #N��%�� 3�,��	O�Þl�<�hWaꕤQ#������K�82�E�ED�"ѿ���	X��܏�n�GT���S\��Ѫ�䦃��H&� ���?�JD���v�g���N�g�#��N��P(�/3A��,�/M���I��9����)wH�� <�
� U#m
h�W��c~��̒V��bs���q�MK!20���9?M�����Ʈg�xsr&YL�w������*��rBb�s��Z\��"sT��,���������<a����.�sTt�tVn�4㎫ԜA��X",�0���c�v�7��ɢ]��X ?G釚��~���'�Wdm/ۣ`�W���*�@vr*&��{��i��B�H��{U��I�p}i"��}Ný�~���zp�h ��>n�kUk�J[0tݞ���-��gr��7P�wmv�d0���	��*�);��ێL���v̓�Y���E�(?��,����UG�q5h�:2mRh!I�tS����#��H��M���L^Q�6��Q�^���{[W���E�������\�)p̬�M�|Z�k���▚�����ڜ )����[�Ch�.����3��N��M������I�jko�d��?�x��xY�#b5�`-E�S;�_��Ĩ��:R��"I;Cf��@�~��*2��~c��=���a+jZ2A`$���3"E)��/.����0VMr�ҙ�8��$>1��m�[���ސxjf�G�vn�`E�o�ɓQ��h̅�������pZ~[���G#��M��-���9�
9�0�t���Q�9���͊�*�k���g2��JU���g!��E�k�T���xn�r�e��
N[d�sa�Y1$Y+<eo��*���|ȥ��r���`D�(|�B�<B��=��y�'�BL?�tr���L���a�a� 6���>L�/7+��ݚ���1�,-�WfJll��2k�杨="~�
N�8�뻦���3�iN��.��!�)A;�6uے���C����u�S4=�Oh�uD�-@�o �Khd��I�����P�ɞ�h��q"��/�U\��nr	>�7�܈���}&�Ma�r���!�*��Sb�?yVJ���B/��_'�DV�G�gfo>9�I�ܒ��r��.��Db|8�^Kd�f���&��T#�%Y�:����
�yK�v��W��i���J.��]�<�W�+���ɸ���$ �k���+!�	tD{7�jHn��@��E.R�੺nE#>�<,�K��65�>T� �!�!U.����1iS�t���!����w�ϸ���T�,u��#�X�
�ep��������mpY� &Y��ߓ�ֲjsi���EP�}Uᾖ)�-�����?�ޙǌ�x(�F��`SfꛪuW[%�m�!���n/��s���wN��Z}£8����T�<�*��;��6}�
7Ą(�M�h9�;#�~i�X����#����}yb>Ǔ1�T���[����o�`���8:����[�|�`��!L�^*�31Z?N(�����
an�(#�N�ca����w�#n'"�=��u�z�F�L�4��Cx��Y�v���_v3*���V���u�KK��Rl��g���V�v�E�KSX
l{�ڂ��*�-{c#oqu*�ګ U�G�������QJ�E|���X���ĸd
��xO�&f��A��v�y�؜4��!��b�cA~gp�\��0M�"J�s�%�����G�[���a�e��"���:����lTZ�۟�-���a�E�\��� %�.:r��Ҳ�΋��XMV+I�Mϡ�]b�<�_�{R�ݒa�˚u�-�Y@HOxCV~�|G�=��v�j��E��N�=�>,�2_x}EdhuR�F8l��-0p�vw�Q�/�6������H��R\E}6�^�����*�C���äxוy��|u��Fc�����q?����I	��C��^\$���W�O�sw62�-��+j��^-N,=Vd�h���}7yty����<��:�쁠.��� ��k�'�R��p������ ��3^���-v�h+]N}�����M�����j�W{��呦 *�6\�ğՏ�U��J�oO�$B�L�t{U�EḢ>�*���&2��p�ٖd}!��0"b��{�� ��[#��P��V����ٙC�HA�kkQ�2�a����WP��a��n����󀱂j`�Ȼ��D9�
r^6�W?K�ʽ}>�6z�g~<��68�Mm}��6�`�A��E�qV���Tm<�"��[Me
B� ��'�c�v�i��yC�%��Z�8��5�i���[d-$���� ��+Aw����|Z
���!n������^��p��g���6�d2�� I�k%��#����tA����B�%�{�k�������G�.Aa�כY���<���`��'>\*C6dd�^��'w� �p^ф��yl����i�q4�Jz�y'�֔�p�te�!D���_��Ы��7L��PV��!)�6_8u	F-I
��L�S��@D#�4(�Q[�B\�gRǾpv�1���RJ.g��~����H+���ċ���sІr+��c���'@�]�|ǔC�{/�R�f��ԛ�X<4 `Ld��ɋ1x�1F>������Ǌ�V��j�e�����Vɴ?����S�\,�G5��3g�r�C��~�e�+���|��\���'Sx�tSSv$)�zb�9s�Ӕk�5ѷ�U�$a��L�ߐQ9`ȍK�Zш�^��9[�������,x�HX%��ANl�T�/�wk���$Q�_��4&�fR�sg(X���nI�����v�g%M�:=��VV��sI��"�X����6H�T�#��)z��� �_�	�l{��v|"*�)��Ja�ܶ���^m��s.��xG9�|�DG�v�M+�&*g��e�O��t��C�c�_��D�J��|�{O�Nx�_ԟ�m��i;��)m�n�ͷDJ���O�/���,E�m�_7����C-�������\�ip�XX�Y����4f {����K�.�����m�ʐ�_{�;	�t���D�`r�QX�.0D4$����Iι��Cfg��������^K�ϗ_��^�����%O�ӂ�����%�w*,�ZĴ@m���x��5ty1�8�aʘ �-�j���⒩�������<�<��_;������zF����{(CӉ�ŊW��|.����\P9e��dZ�[H*�(foR�LD�`Wꮮ7�P�˻�j$��@~�a�}�V�>��QV��L!I���\DBu�&픩�~j�k�t�U��#�ǘK֪*���4��Mp�����=�s�C���{O���}�6>���5��S$��u;�k�g��J��B�F��p�Y�ks�*���7T�r��/�[�]��{�O��[��X���Ņp%��J�B+}g�3��;�	%I�{Q�%(%2#3^f���k����=�uV�p|oo�������lW��S���f�H��G[)���ʳ�-���c'��!��}��8 ��*���A0��'��Z�s,|��VɅFBjBm��uvA���Q@�%"���n!�a��0���)�ڌ���S��d��?�'P��̫�:��k�*��m��9qVv��Q�̀jTCS͡V
�^����Im9˧��;��xt��eN@��SZ���KS�T�$�ݵ�	WF�=H\p�g�O,$���,�os��+�©g�e���8�j�Ί!i>���lox�<�G�.ܹ�vTℼf���;Y9��n�:���<އ2y�&�lj!��*C���Pic҃P/�0�d�r7(�� oA*�b����Hz���������ϔ�+M�aQ�>;k	k���:Bh�'J�hZ*�u
	a��A�9&C���?����!јW3��z�C[I��ƼT���Wyi{���T�2�%C�`� ��r|J����)�F���J�-&kH�1��e�s.^E+�z��%r�<�Q�@�H�_P�V����ՠD#txʰ��􎿗S+������}#�c��piQ�߇����R)|^�L�؈�A�Ґ����g��}/���<�69�ɫ������b^�ŉ(�Ĵ��9�t��|0\����F�[�1�GEBs{
't�x'����bV�~Jr��EƁ�<���É���T�I�N�^dP�b �Վ�Ҹ�F;�.���r���򍰣�U��ʅ�T�1Hn��5���g {l&L���߸<}U��!V���0�+�VR��/��LQBp�����Мd����1t�㈒U�0��-`n�*�:*�H؉��5�]O��E�ߚ�ؾ��F&\�|d�	��-;�w���ȱ>�� m�1��!�� �#���,$����1���UP�ʕTI��P9��ߡ�-��k�S���#���w+:"�������o�m��5�U�MZ�M��$����eRJ;6�-�+��_t��a�$�j�N{NG�ݗ� �tx���A$ k�i{r���iC0`4��ZL�*-��8
(������:�ݕhLz!��i��\��܅#�5([�+����}�SL�a�<aWh7��S�]�>�AE�z/oD7Ӹ�v�<^��Ab�-⨛�-hY3ڳo.����}��[�� �e���'����������Q6�K��5�8�d�
+��Y�M��{P(2jy	��P��Zk:��T_���_��J@�Trx7�o�m�dE��p�ԬMs�5^k��ƚ���4������"3��!��X�6��tc�Ř�s9S3�+��<r�Z"#�S-a>1�$���L�[�'׺��x�:�8=�Uz�-G�asde
�&ŷZ�����3�R�����Fb^��=^�ߒZ-��3&�h���6I�<9�Z��@!����F�Ą��ޯ0�`Mtk��HoytƩ2T��ԉg�b���:_	ZC(�`�E�o֐CGhጇ��O����Jɽ\�q�9cY��P�U�� � �'�cn���:2⨺Zy[|�E8	��rf�شJ�%)ZK�Y�"_ LV��2��%qQ+~����.Щ��ʤy;�H�Љm���Y�p��CN�����z���cc�~����S7�k�V��x�mIB�fºN_�y�<�������o=�[I�Z��
p�54�Q���Uy���z�J{����l�\|�Z�[R?I��G�Q�K�V�,��7�kz���h�g�\�	J���;7m�)����@��g���^�3��Ƙ䭲�1�=�V��1D^�}OM���W~���v�e/H�9�Ϯ����,v^�]$�ځ�F�"<��bvg�V�#�v?cLnhb�ϢAؠ�|&�&[��w;�2��D��>���.xL�}��Ei&;;5�ܴ�'�	D���z�C�`�xO{s�M��=!�&pQ�M��#�S٤��Y���
w��$If��#�����Lx�T�I^���i[c(˶d.ӂ���\�L</f�2���<p�b�X�{��"6%y�D9`�9��^Ux�D���BC�qBd�u�H
��"�ht8����6��h 	��+�b����fA�cS��n�	x�w6O��U�{��г��Y���񁛤 ԥ�J�dQp��`���mY���UƈE�6��d�jI��8���r�-��Þd�c�uX~�� �֑<���D��h`�	p1��~���IK�f��BO�yaߢ��(Zu>�|�/O	B-3KԽ����ж݄?�|��ðRL�'��7�"�_kE)�OHܰ=��K	ӡ�Ѫ�$�G���󨔓��L�"ar�����'7�^5���1Dc>�,����*z,��[`���:#�ك �Z-���ϭ�1\�)f)�OR���)$�N-x!͗p�M�h8:�{}*6��`P�_�q��D��	��Ī�cr�j�|����8EafVL��#��@��qV�)����%��˔�uv�YaX2��g�Y�G_P~��uS#P{VF�g���_����wq��8U�i�+��g�?9�(dUq��z<�RjD��t�Ik����U^�1�������AӤEP
���a}Vô�5�Q&E�.�B�ךC�c���޺Kd�S��4� ��;<�z�א�l�ڶ�oʌHٶ`C驏g$Fp*��x��=��;ߟ��ekr-�bv�F��^��K�L�M3jMeu-��2�`O�B�
&9d%���@�
ɷb�H���(�����m�+FB�g+�>��I�9h��D_���+ ���'1['(n����Rt�g�Y!�i����P��Ҹ�	�U#��3��f�1���)a w�ժw�K7|�wc�*{��7�Z�k�H�S��������u��H��W6��f�1��ţU���{]ݑ�IG�ByJᢵ4�^V��R��Ё�p�I�r��ި�b�A�Y�.I��-�$?�v`K��Ӻ=XB�^;���>��l��	Ԙi�����<���ᘘ�[��0�
KN���
��>����3}r�¬r����Z�c���khP����'�і���iy��I����䌝f�<�7��<
l���%�BR�2@��V�UyFg�x�����Kx���o=J�8���_IAt�b%�}��~~4#L`0���H;�FK��u��P�|�D�!xS�P�Μ�R�_��S��%{�� ��9_;�U���џ{a�/L�6AΥ1���O�R�5;:S��Za��.�mBbu~���}@�<���Ut[N~���6M�h�O

s��O�	� J�)+��=��>> ٦`[�;���� <d/��;���{mf���XN{ �ۡI��L�)����|c��@|�X�%-���]��?��X�6ci�M���K����"Z,��N�P���������
��:��1��_�ƑH�W����w��X��ԙ�n"���_@doi�"$�&h1S-��T60J�$��3�-O-��f?�MJ��؉�Y�p���Q�]$ )����M�3�KI�� ����)��R������q
&zNz?=[�&�\������9WB(��ٔ��)��ր��;���k� �W�5�F�9����C���N��b�=).�<��w��n>SY���i�*�U�J>EG�퓯,���pkDC���nI���OV%����|s��[ǉΤ��mzC�IR�w�K��ʯ$I��mb� "���4��;g�r�{v�*c��@u��I������h�3A���(;�L��O;�&�gA�>3���}q#�2z^Z��8/�Vo&��ɰ�� �kEXIC��T̎����qk��BYO���7��ܶ�o�q��X �zA�頂�	?��v����{��C '��T��],�a�:�#h���/գ;�(��o��4y��솠18a�V{�o�\ⷄP�m��1[Ċ~�Z0C�B�[G^�)�,F�\$�w>���4T��Λ��̏m��7������k�w ����aP2<����g�M���d�NA:e[���8��V]�'��V�H�kM��:Uʉ��{{�@'�O��Y-�Rf����C���k���I;��]Y4��� +1�`�'wC&�;� ̶x�*n���gm}���N�]v�Z�e�>I����~�w5��1�h�����&���n~���9H��͇~�Uw���f�|�I���J��tU�b_<E'Hm�6��a/�N��4vO�Kq#i�f�x8�J��GsYk�㹠� vR�"HLQ �4@|�o�[���MTY`oe�����M�Kߓ�Ǭ�7?t_�
�2�V��Fmdx��'4�	�#�i+�U $QB8{����I��~i&*�(����JHPϕh�h����H	��	�]DT�Je,*�����e��#0I�eӃF�*V8�5���Jh��c����Y���	�9�IZ�c�b�h�Fڱ򤃔>!�>��¡�@}�y�����n�2�R� ��crl�~t��r�Őj��%$�䞶x�2�m�*j��Im��0wc�v���:A��P����Z>;t��3�O6�� 7b1�l�w7XZ�(��P�\;� La��]+�$�/�,� z�����Е9�0q�����L���L�����&}Ѝ��B�� �����vzi�t��/�n2��YWGVLF*�4n4$֒h�؇�kA�:\�C��ɶp���4~��m�g̪�=�E��:�]���(��L��%����i�6ͮAC��GC��KM���ePH,�5m^��ÆA�,�j�X��7�!D	�����F��y�b{�[i@|���8�3$�6 C���d�P] V�� w�����1���m�8Z5�L�����sM	E�=�*?����vPC9��l��1�-�^f���+�L�!�X�2��U�e��ْ�/���&iߜ�Bo���?�g�-��oI���=��}=���~�H�.6�o!�A/�͆7?efE�V��R�y�]bX�H3Gk�M%�yy`�C�Ϙ`�횯vV�l=&f}����q��ռ�����d(g~,UHfu���]l�P���4%R�������۬:��Pb-f��M�޳~=RaDC���F��Y�_u*{K`�n6n/� ��&}1�NVsI7T��Ѩ�tV�*�e����F���=y/��
��_�$i�2�g���ٮL��I>�43�\�#�����n�u�R�V�%�����}��[��EƤ���
h��Gz�@kG�����[\�h"Ɇ8٣�1m�b�� ���܌���og�4�2�{&C{�0q�2��a�����\�(���Di�UJhE�l��u��xW&�e���4�q�lyZ��ꌘd:��	E]YG�U�ŅNJW�, .�a jL�E���bfSw������i:>�:���wX,�#x���@Ni7a�9������FQ;<��A��op�-b�SE�ւ������Z���7ڹ,�!��K
a3w�F]����}`#h@.u�KN�{]�(@�V�, �?��s��jW���օ��=����rl��W�o%�z�夯�������-�O�_�'Y�W�۾X�PJ>����ra`��X3m�?����I�mh%a��7
 ټ�
�a8������ي��8�$왕�_���x���J��C\%��[TƲ"~A���G=�A(�4d����%�$��T�����"TiRBk��lO뽰����DG�(VR�^i�G�
�DOI$�Us�)�>�<����=b��f�_�3�������C�Ï�ũ����c"��c/���DD�oF���޽%A�0͵x��$i{ ����w~�Q���f��Rs�ggJl0�D�$��,��p��w�ի4���}�v�6T�+:��:�ˌ �����f�.�+M���:������F�5˼R�j�rS�����$���*)��^-����]�����7��T����fh7#��O�5�s%����	�Bs?�=~�8ZD��N�%5m��0��I�{x���^ i@h=|�b��iI�����b��8u���P����m��P��&I���G$l	� Q*���[���֑e����Zb�A�ب6�����^ĕ40��t���G�逴d4�rcN�<��2qRt�D
���gk���ܑ�?�kؒ�s�9l"� nK<�$wt�´�����<�w2^x��UL�` �C�*J'w�J(u��'��H>d������ԛYP�����Ij�|
��^G��ĊO�+w��V��^�i`�FN�����p#�+x������M-�,�Ç_��B6vS�0r��u�vvB��7���#N8%Y1	�G�:{o$���� �p��1��O[�lK��72��~��,�*���j7��u�����v����?'t��dў�	�O%O�^!�t%pt�6�_f�|��7�~U�!^�����5[ps�FXRf5���D�W!�IX ��Gtm�{��p��1�]P䳵�]�v��Ը�v��Qu�������>��dv&,,��7�l��CS��G9S�Ʈ<�l�Q��S�%��A�W0Y�!��@�3f
�,1ӣ�)d�>��B�hŋd�?����X��z�����aV�ja���
�]j�x��M=v�4)�տ���6�)*�n4<�E���wx���_l�NQ��߽��*��n׍�Zh�=c�"6���*�л �#��'�����C�&Y�-�v��ӌ�Iu����)�?v�,�ߊo
�<�>�i��V��R�Չ �;�M�?�Q�r}�����`��w������S*.��A��A����pN�����"�B�|Q脨��e�)��}z]���g �rЦ�ƺ|� K��]{6N��'t�ڡ!���;���&�rVS����X��*���?B��̯��uVs�3!3�Q�$�>z��D �n���m"* �0s��LD+�w����������ǵ�s1���DVS�K��J�( �N�j+���^Q�f"_����p\�f�������Ď�3Վɧ��:o?�#�U���/��-��$PB��ྕ,5�fr!�R���mC�����O-A���y��>�=�~F]�[s-�����zz���t3�DW_�A�@&Y������k3�37�pJ�&�u�3�惻��~Q�u���5���α�ɔ����Ȏ�V��]E�ñ���yBn���$@�K�2KndIÂq���_.����1TLb�uu�$:�	:%�>��w���I��R�k�dn��`��=�O��q���4s�V��f����q�c�]�G����Ppv-�e��� W�*ޣ�l=��8��L��:��JPS}�Ǆ�51~,}c��iH�FJuꁱʢ�y�4��ʿ�,r��I+�&�>kv���?3%�lr��f{��^���?���IrC&	�XZܮ2$�6
Z�ҥ|��$۪j�������LB4,_vnH�]�$�U}|"s�U;M[�8���iϮ]{�_���W�ͷ�6��-�n�b�YR���ӾR�h>E�M�M�a&�cJ�y>1���f̿�뎾�����������:� "̢(�Rſ;�C+��q�nT'����w�s��1�5���:����T�Y�;�[p!C�J�+)i��F��>W+j�R4Z0EٹѦ+��X��2%�� 5�(e��-����t�#�U�w��@��ׇMէg�ҷb�[g,���r!�wfT+��0������Ɲ��8��u�X�p��F�@݁�.@^�+��E��s^͎4��pB��m��M��&��kFo
��nn�f�M��"��Dd�&;���b��ccQ4�P��7
�����-�#�fp��TYL���
�(�,�|�41<�8t뺋�c�Da
��eg:��=���<W�A������:m�H��6E��K�N�ƪ���FZG{��,ܿ����r����`r����V� g0�Y�]���B�i�vV��9���W��H��-	B܎����]Y �l���R����ȧ��ݬ�m#���U��6�8��V�,\������a����Nƿ���O2��D��������M���r��*Z�÷�v�	һ�͋���K� =��v�+��+������w�`گ_`�g/s�b..Rɮ.6_����	�����io�d�� |��v6��V�A���4�ń!�a�/�NF�����p�B�_!����6W����Q�'�)�v��#�qF�:�޲��!�ov�`�fjb/R@ cáOđ������I�CMkW�jb�P�����z�BO�ޘ���x�"�u
|��zc�z�ԁ�Q�oC"����<��>Yw�"`QT�<4|U�\�]=ip����>�އ7�Ә"��'���7 j87C������Ta�l��Ȱ��3�n�4Od�9�FP�ھY�ݒB|��p����$h0^��v���nn�G�����|,r��h�Offf5�W�[\Ա�v1��X�?w'p���X�N-й�9�����D�?��s�Ͼ3D�ͷ\�;�̀x�cz����#3�����q����o�3\މ��J��M��e��?*��%��s���2�/� Y��Ȉb�`iȊ�����q�WA�����˹T�����$�bf�҂��,rWŪ7[�g*-F��\�tZ��4r��m�g2dy:5)")X=��e�gݹu�nF�b�%Mfh)�=< IO_��	���Y:8xԎr��`�}�]��43�o�ѩ2jI����3��X�O��K<��SV0��.7Q�Ť{x*A���$�&�%}��L��%��[��u��lZ�[�#���Q6�F2:��tl ���OYX�v�mDB��d8F4,+V��yA-6�`�5O��-&-lp�Z�}��tS��,�!�`+��A�Ϡ������%4���}Ua���P	/q�_�Lm�B��������7"��L]r����[P����5�g�a'�}��)0-%H�kg�����@��E�ŉH��Z���u��:qDbT~F&����ycJ�tp���v���Z[!%�K�D�m__o�5�H#��,�ֳ5�p
][/QN����ݣn݄�8.�;�e�1��(5Ĵ-Lc!���@�H='un��G ����v5B�6a��&��M�7*�����~�
�r��RA �ݝ�푖d�\ԕ��i/We�/�,=�t���e��JA"*�����#�����&�OͼИ^/�����xz��5��k�՟������ʿ��'`л�� �d���8hf^��;3�a/�&߰aZ2���R�Xɭ��5�S�"���*g._�z]̄Z�	m�w<��$ ~ʏf=#�WaD�Wb1��Y�����pcr�֓΃Eu�4�h�~z^�Ģg9*v{GbH�Su����q�lG9�__T�	d���9��%h|&���S24�����5�����g:i�@狼�((ś �,A�Ġ�T�%��c�jfp5�M=ni��~�ɉm{�(�U����R :ނ�AJ`ͺ�q�[�T�߇�i@-�����Gہ������ZOo��4͒�����}2�@C�� E�y'g(�-�|]Ѝ��(BǻO%��;�t�����#!Z�,;���'w[we� �O���=�X�zN����gDA�g�����\h"�5]����{�g�H��p��M5����;��bi��Ll����"܈��1{�Y�`\`��mR����:�)�@jO?.D�X�Ħ��6?�q�3k��-�יo	��$HȾL�8"�p�L�|;��A�Tm3rk��5������@�sa�"�ㆍ�!5:�/�����J�</�Kݗ�S�<ZE�4�]��� �o�Q>�a�36X�b�Z���������5��ï�/� Z!��'�����F5�
1�Q��Ð\ٶP.�,�`�.�����[�����a�IC're�EB��X�,0!D�)����Y$�2���Ѳ�D��0 ^ .8|ņTm-��9L�k٩�����O�`f�#4�R�S�6�Y%>}��՜�o=,k�S���.��P�U;��STsn�w���$����V�Q���$P�#-~�G��t�ڻ�E����0�j����DR��c{]��Y�9AG��!S'By9����K��MHR�hƂBm�,NZ��RC�q��DM3~�'ߧ%�$�Y\q���R��9L�*�g� Bū���Hm�j�0��'W��j� �(��,]o(�{��x�7�Ƥ�V	2���]\����{�|��s~q�C�Mrޔ$�
֫`i�2Emz�R�`��K2N�Lg����jR��U&/n�
��c�
�(&�l.�֦��b	e���R���߾��&W�]0h��� "\��T~`�_": T�؎�k-�(��9x�0�=�ej hq�N^�Y�r	W� �C�K��	t��	{���z{��-H�q'��.#�"��b�] �T�NJ�@�/-��O?�O
[S�O!��m~"��j����y�|C�Azޗ�+�˪��}8�����Ʉ>�\h�?3�k7Hɂ��?ow��dGv�[�H��^�Ħ���1��K9��"}����芾�i�(^|��p���I_�K�+�;�(p���d��`=u�/y�`�700O;6�3���h�r�%��˲�=1r�㷞k[ѽ����&��O�K*q�2��Y~��L�#����dŘ�Y�Ҫ�=77�O*M:����I�O��Ƿ;�P��r��4x���v���s��⤖�8�qs(�w�5�� ƗZ���yn�7�P��AW�4�̩�:�|��4)� ��� ����̰��S�J�<=xj��k!9���A���:��e��3X42b"�(��6��HJ�v?�X�]�Q	��J���7�Gu~�Qj0��_��1#�5�����ߓ�DJh��t��x�� B�����\����<��+���C�=)���x)����R�@j/� U�)1C�.Mț�^vrL*5q� ;EsL5g���"S�Y��������k��2��-t$�mCFޅ�,�Y?��gۥE[ >�����)��k�O�X֗q؋���Gx>2��iq��gg#����2у^$�d���p����c�+Ϫ�C�gw�`B�Ǧr�wgX+J��lh-VxC�ڬ�pq-ZU\N'��!Ֆ5_��d3��B&�[�"ǩ�.)��ED�5�<l�_�z�K5����x_�ؗ�П�@��BN�X�J��q����@���(c��3�)��ʟ���.Ƕ �.����}�T�ǷN���(�_��,[�E7�+0�[b- �������}�$�>gXƀ�jc����^Lӂ U�yW���s���$F��>�����2�u*U����;q�f�5���D"�3`�Є�>��;K�dx���Y$j�Z��8CA����������X�fL��j���E"`�5q4��G-�eģ����B+�*~�(>��7�.���+��@����ʷV��ڣ��?��9�h���R}g��/O�o΃e����RtT��?���uhC�'�����p����m�H$m�A��)U�"�"�.Θ���&�������Y-ŴQ|;��d_�
v�̞ϙ���}bO+�){[%����� $+��
;㍄���˷�������|n~��W��\��ڄ�q��K�Ɩ��#{"�5�.����1]Lbk
	҄R�|�[�5��#:���>G:���t��C���/�_�Qx>�Mݼ]�Qe���!8O�#WHD��ןQcm.ȼ���}�dzk�	��˚�}Y_+R��rrg��FǤ��y��U4��Q����ߡ��$�kUP��V�\\���LR�>�C�#B�������8���XZ4�B'�C�$Dyh~�q�mU�F�)�I
��p��c�[V��g1(,��_�J�@+�{'���hhz�#!���5[8���	ҧ���_���c`;���D1k�u��n�
�8^��������9�I�_/ˁ��m� ���t�b�I�%��_3�}�a�%���jɇ)��2K?�z{�3�빃8��S��G��R�*��V�7i5	�/y�2<"��
�U�<~Lj�%k7S����a9��7F�X�(���t�WZ���a���%����à�:^��֚^Z6q|�������2`�H	2vb*NgR�W��X���f4En����m<�����ut ϵ�4o������_��՚X?� �eխ�z�ʗ��)��/���S�*=���$t��̟1�0��c�so`�{4�U���ހ��p>���k]lǦ�n5�8ܤ��v�}HI�ZWC��� S�eDm�Ί
+9ڡ�W%Xr�^������Ҟ$���+���@�$�\�<Qv1���qٖ|;�)�a)�ҏ�y�N̸ۭ��k��	ԍT|�xކ9�ڈ�}t���n�.�M����	!O�ǉ��}��;��w����n^_�̚x_������9)T43�^N4�κ��:�1b�{[�,�=�&��� 	��qGa1�lQ����Hq�,޲P.���!�0F�w���� �Հx�]ilt�[�Gɺk�CAU��������+��V��8��J`B���z5���i}a;$4�4������9�{��m�$t��JvV��^���(���3�>3�:�|�yɝ��UA�~���:s���!b�����b�O->��I��i���T#	^�
(��`�Աx
~�%�p���\zC�,h����x}H�p��K�ѶX׫�~oK�����ݾa�w"�16�d8ȵUR�r'�u�v���=���s����4̈́��z����$W�������0�YQ�`��.�p4�!�Ϟ���y,h�>`5kh�����@�[N��"���Ww(pȝfK��&��"�ض��;��ȅ�+�^V�*H�G���4��~ǻ!���	
���
�)3#���FC0��S��L>��3��ܱGy�.�}xX��NX)j�ǽU�L�0N�@��2`ny����]D�˖Q)��M"ѕ�l���l���	���P8(�g.2���TES�R�i2:!Q`���zwQ��+�r����{���7O��mcgh�E��Kq�er�J��I�����Ucx����z�x��)�����@}�1<�T��O�� CN��9��+͛�F=l��l=�H��9kI���;ƃd	/(�|Y�ܸm�2������<��L����ոKāxP�j��
�F�P�]>	*��z5u���4���?aD��Y����k�HL�6�{l� �,���϶��1���g�>���t⭠J�#��<ߋd��%���n���D�&����(Kewha�F(�5�f�kM)�l�춸W�NFԈ9���;(\oa� ��hn!��nN;%�F�)�������˿ �r�Q����u�{�h�����
n@g8d�:R������r��TKJ�-�����PVm(rfs������'�	E��//^J��,@g��2FF=��T����5�<2��n�#ߩ�X�j8zn�keMe�KY"��/�C��"J�>s��C\C{��6�t��c��p���������on{'|%����J:�;O��=\1ݠ�ݵ}H��X+�ֶ����yV�y,z+B_;��)����I_�4Sr����\ޅǾ�S�QTy�O�D�A9�=ktWs�9�D���/R�%���K�`t~��z��w��۾v�Z�A
��me��M%��Ewc�+�y�D��me�\i �j�|�j���]�"d����̑��OY����Ľ�� ���
��/6h���6�^���`�p�,8[����W�G|�mI��/g��,�TM~���Y�����au�	Y��V��Y�wš]r���������� �?Ӿ^nC�0t�`���Y���T�m��F�2�s�NZV�ϹQM�>�u���%�X-��s{DQ�q��̈�@�F�ԍɲ�6�&�����������N���!�a���L*��b�zQ�Ns0���#zH���%9�,���{rI���yZI] �pդ(b�� K�G����o�j�)'d�D�Ck�,�G�3�@��)�Ո"
m]-��=��F�^����&�Zo:���!и���e��+�·:�v0}���F����LF)���Y�ଣ/ B��5X��X���}:R5�"B�p䱌��*���S]dNb�HŵqD��G��
���b((��!�.,�u���E׆�4D	]y"�/��;�;&�������+�l���F-P�-I/5����@ӵ�5�>�/�����LF�\����e�+S���Q6˵���]�������6�6���N�~�2�s3wo��A+v�h7��C;�W'7��z��K���4*�'�L��� A�O����1��h]�]�1/��*n�^"4eΆ}8x�@结Fv��69�sH�=�V��Q�0����U���^���dԤ6%��BT6�A�F�� �g�y[��A���IsI��c��9��<���p�H}�֕���;�
պy���6�}ۤ��䧋�~''@5�Ѹ��oh�&�Lh����0���a�H𹭭������8I�uK�(�dV���13|>d�5+�$��ș�V(��5��\�??�)}$�����sN0��:	�$`�Dt�
:�dkt
��.BÜ���B'g,�4��>���Rg��
BE�W�%'#a����}���wF��+i������R�h���>�����qm}&fD7�nZ�N�4�1�Z<��Ɣɣ=U\-Sc�DЂ���Ƈ�6Mtt���ؠ��q#�Һx���edc"Q8k�s�zM���M��jd�N�s�Q  ���W����NE5 !�.q�z��!�|���M��15DcG�2�0�_��9�IG�eK���3��|��Y�ұ��Z�1aûo�$��h�����U��K
��Tg��
����u_�;�t��(��M%�����;R���{M��pr��{N]bڃ��n�0�7JX�l���q�+(ѥ��~L�k�dQr�!��z8�/ �b+DV��pAЍ&Am�HД�3l%�Z�h�l��o��z�WQ�n]��>��[�lҘ��F�CG�i��G�6���?�zƜ���h��%#��zn x����jeZ��ժ
��/!�������@��#�y51�:�V��_����&qk��΀84�/��D�x���N���
U"%�(���a�N--�2��$����V���ҋ�14����U��A
y��N%T����d���s@Z)t�;8�"~���0!�*�.�,YdIn.��m��C����L+��J{�>�^����� {U�Kӫ�;��y^*4�/���%��hKG��AX��=t��B���m���]M�T7�#a�`��+З��{l� 9@ő>�f.BGw<i*H�/�U�kG�i�������̈́Z�o��O��P^%F��L�Ck\_Zw0Y>�҂1���I���W�	��3��B�3�$��}�ʤ9KZnK������3r��N�*2�q���`\nΖ��/�������������[��c�س��F ��P�*mc�X�)K�Dv&�V E�z�sq	9�z�:v�@���L	�>��o?�0�F *ha��P&�"ˈ#��swL\��{֯oO2d.�C=yX�����I���A�4@~��j�-#B5�I8L���ۯ?���0C��1xf�Pݎ�6�0��>��O݋|!�(�G��j��nA�0j<�t�R�@H8�n�妫P��dA���}52��.Pp�;!�K� X����[�,
h��[�L0r�����̼HI�V�8{�`����U?�h���H�fH�>#]�z=�l�V3���af7U���w~|�#W����1�Q F�@s�������	��~(��*Au���D�5�k��˜	���.=����8����;�*��u�p�*�&b���|D�܍nB�X�L���������@�o_� ��C�H��k;ۑ8�z��K�n*�1������֯x����g	��PC�@�v-i�iB�����hcRS ��r��f��O�H����c�^(��@�����P���ѐj���t4����Q^�+���"LY�p�y�xrU_�o�+%�]z�<x��fmxpg��r�a��1)�i��=�,h�*����?�A}�DTL���n�o:3���+#��zI�ޅ�����T��4�0��E��>��Jd�]-߰o��K�5����̀����K�S���|(����uV��dQE��r"���fO����|��/��$M!R�I�΃n�!tO2
���'7i���`b)�g�骲j�ӱ�� Ck�\ȟ)m���HӷhS��,r�O�K6*�Tl�B�n��aȨ틵�`����$8��z�C�"�༛7zi�!���.�<V珱��� p\y&���8e7��v�a��@�����ΐL�f��I��VUMVj���s/L��׾nhƬ�kM��(W���y$�n^ת�gc
B;v
�[�`�7���������X����=����G+������Ծ��u�:���;�0y�3k���������,J���
����t��n.�/N��6��F�Z�`[�������Ir�e$e�����J�Ju9#���3Z��7ڂ$D[d}�"�.'c �g�vH����1x�m�A���Tr��#�#���)I��-��8ʦ����3��=.*%�n�\�	��X>�M��c��UکU���-�TM�{��W��4�������@�7�i�Dvz��Kk�� uR){x�<�+aM�D#?7���`z�$�RO'�G� �� ���ߴ�}��회�!�L�+˟�2'앪���A��n���#�n�e�	���I��8��6�4+�*BÜ1�,۝��-Ğ�#s����i-_�D�Wu�"������2�Hy�v�P��i,�)��5;������rC�����[�(a���j8�M�ֵ$�"���i�c��`ޕ�6�e�T�Zl+�9q2�s�໇
���a���Г�D�^12 ŗ�ymt>��O\|�F�y����x�iα��/:��ʖ�ކ��B��jJ��R"w��'������2SK$%-�N��m���Qk�e��q�p�_�����X=,��e�1������$��t�JyG�Ru�$�OY�Nܘ� \��!���rmk/��i�E�׶vKG��Y�$�E>��A�}��O���z,4/xd︢/6��|�b��uºnA��l�>���\R��˚�]$Vbi�Ɛ�	��Γ	| �#��?�LO|הyA -S���eT��eG��YY�驞��m	z�p�X�V1/��Ǘ	�G$��l��$��XX���ރ��á"�x��|��7�SE�3K������K��ǻ�u�o�o��VįD<tخSB8$�Cc��������
�g[� M?��;�'&���B��
3�[��j�<�Q��t��˯������YT�|.qy���\19�[0�����K4��	ZH3�*�l�'��T)�����$����.���Z�L4��(pe��&'EV�����,aAM���2
V�� �����$C�r�V:7�q�{�\� ��L�)��	�9l��"/�Ě�s}�c�"�5��̆/k)~J��qU�r��f�~Iʛ	��`>��Rںl�	���K��|\�*R�P΢��ZŦ�JiL-����4Ͳ.����%l�=]k�9����,~�'-����!@B g�k��d��1_��v��	d�����@����C?��T&�����WHu����D��E\]���B�xP���n5jN�F��6�.�n$��^�m��˖b&GٌՊ��KZY�¨�y���j�,h��Y	$�++�0VQiDP6���׌�<I�B�{�a
@�?�hZϬp�Qc�C�|4�a}/��4F�o( �6]�u�Ds���k�\+�.�26�o�w�bb�x�?'���]�l��`g5?��k��\�{k9Ԛ���D"�l�#ї�LG �i��������WM��Fj���D�;M�b9�������\;���3A��e��N��*�D
Tu
��.�9�AV�Y�x'㷁WzO8V|�\�w�����_;���P4\���-/>ϻ�y�6��P����1jC̥���)Eǔp8���eF�6�T�{zyMO�K�p����xN}�KJ��MOV>���3𡃲1�:r���+�RRq#ѕD�����j�O+�n	O�wX$4�ί�ߔtX������~��/Z��#YL��u�� e�rͰV���E�M������,��lSL�kLc��&󹥷�/�&��u�5}�x>�`V�
����_{0qM]���o���v���1��%�U���2I��D2uK1}1���j��z��&�M��>�ᷬ1rQ������W汚��5yx^�|�#�� �?��q�8�hk~})&l�ˣ�=L��?�J{�Z`e���j㼯��-�N�@�c�n�I #u3?J_�{w�mu֥[�`XӇ(�N'z�D��>���|p����<�.~++�s"��*�Q͒n�J�k1�)���E�B@�q��W�z����5_VDLr/���KN�L=��bgݜF_���sK���5[,*�aJ����ai�k�2<��q]��\�6lM�xDN�פ��Z�s���p�S�d+Q����M@u�4E��n�n<ԑ����b�bϤ�Z��?�n60��G	�% .Ȣ�+�~�}�������IX����XHd��Kq~��4����_S_ed�J6蜾(PB��/���~���!��̩��q�()��,���"@ ��~f�1���D�^J@Q�a��V�p��Ӥ�2 ����TY����{A�ϲ�9X>�:����?�xy�h_�&�F�h��[�����(� 縵���G��%+/S�3���'~���� /�d;�ς8�C���X����)X@�,��V�'�!F/�y|
B�
I϶�־b� �K�I�q��_;��[��Z�S�4�p>֥y��8í?���K`F��F�)��$u	�D�I�)��4}��9����RO��)ڧ�p/�/N(�r�OX%� �{��w�^ }�.�a�����Ϙ�����"�pⶺUu�x�����ݽ�Y�I�
ӱ]G�����kȥ&���;�.Wu�!e�1HF!�ݰ��
�q|ڝ�85Q��
asˣ���\6�2�ʨ��Pg!��A9���-(�.Ńy��Es`�S�~A��=ʻ��NИ���/#��v�*��G64��ҹ�fl{C}�&���i�����ϰZ��$h�}�ޭ�._�8ڬ�"��2�!�=��9��-�Bd*C�����O����c��HX^�ث�O��2z&����v�R�(s�)PjS�	�j+x-&�?�ݯ���>�1L>��+L�X؟�e�hT���[�S��p�TJ��QՍ�h�ø"f�RDn��-�c1�����oJ\��K��	,s�h�#_Nit8+�B�-�N?c<�x���$5�{	JW<øzE	�;�ri���O�Ie�C�x����
v,y)��f�&�Cy$��H���xf^���8�bP�*��ˍl��ZNw�4��;�Z!F�N���h����v���z�8��V��D��N��+rx�����})0m����|$Vv�1����uAy_��	�f��b�g8�TY���%�~/��q����؄N�sN�'ǚ-t�Y�.n�	�?�L�������d����x��Kޭ/¨ik��f=�v���I���l�/��6u$Ё;����Z��0��b�ߍ��f^צ܇�߯PTe��Yoy|����B#���$������s=o=-���=$eޮh�@�E|��i�p����(/�2�d$���
�Y�g��Ԣ#�&���� ����<� �XSt^�:� ���ýB�h �4y��?H��ć}�f�[6,d��fjB����0  �����z&�R\>���\��mb�*��B��y���*�y�5,�-fz����r���o���|O���ۭ��}}y�@d�5qm\�����n_�¨7�܉�a�E�6Vg�Ϝ�dH�s�Z��-H.�H��dZ(��V��t���ΰ�pJ�����%�����y��2ֺ�x|L	�e7�{���l�񩺺)~�����}�!ܴ~0v�J�kn�A�Q� 8ʒ|Qw�M�x�8�
шD����y���@Q��5�J���Ch+]㵋ȵ�I����P��`���}
$���H��
��?�����K���T�UV�t�E��N�9i��B:i�s�+��̃�6&����n�^ H�z)Jˀ4�k��
��'	�<vgQw�����q�ws8����
EϣS��f�F����׹���5 ���C��A�n��?ĩ��`·���R6�r݂`�N/_�������ԋ��b"� c3��l���|��H�k+x!�=u`���W\�]s��ǸW��l�w��^;�Vo�/�z�C���w'h���1�'��ҝ��������}����-��QE.'/�?��=��h��
mX�U�Ê��X�\p�7�r6��<�9'����T_��2�5\��M�1������
YTt$��!r��a0�{V��ڊj���2��d��L�n�&;
���J��]Q��2y���J���l&s=Ɋq�T��7��9���J۴m�oqb�N�Hp�[(~4|����;2��[�ǃŉq�ݰ�m���m��{��;P_ZE���R�D-����t�t���T�C�bxR7��S����o�W������t�(K�c>�}(�g��\{ 7���ӡ}�S�9���n:ҹnI��N�dԫ��4�ۚ�ה'e�2��Y�G���z-�=��+����y1_�3V�/��e�H��i�*]ԃ��{H���X��t�B$�w�T�>2����9p�q���g�B��r�g��Ac�j��� ����h�<�����r��N+;���bNz�2ʙh�8[?	Q/�a|�����J����������� I5���}X��,��M'��~�p��U݊A�u�P5��4^%"e�F����RV�e��Y�3���E�!"�Vp#���t����'n�����;��*���ˆ� � Zo(�)��J� +�Y@�Z�t%mų/�]��)% ��I#U`l�w�Φ��ߕ=�8�H�G��f>K�ڰ+A�^�mM���`D�d��R�<,5���΁��rE1Ǳ`��4�M��I?�B�1D)P.�!��������V��B����΢S#S�������HM%�A�6���=�c�8�d�Z���rIm�od�R�C���Hlb$��FXP9�U[ >�i=? �q���Z��I0vWU�;���f���iBGGc�qٽ*,��>�s=t�2�>�:�(��:���3��U�c��!I�4��%��xe8C|	Ar_�@�Ś\���͙�WTб�";ut|'�X��pE�	��Vy��F�� ���]v%�;����S�᳐*��-x��jo���W	$!F�p$�,Q8��f�i�t�^f�C_9U;�W�˦Sl%n�l�h/��L�Y�1�RmH 1�o>�MnHpr���Q�h<����ؔ[��>m+��5Hɴ���	~5����X\�ZILb��, �A�f��@�ܳ��2d{6$#��t�P$��LS��*t�|4Q�Mtqop�˻G:��l���g�g�O��ѭ�v�rG!�\x��x?�[vIЖJs^�[:�
�Ͻ�a�ۡ�y>��T&��Wc�g�Ǵ��{�Gm/6��`�]�e� O,6�ϣe5���!QCtte�h��T�
�GH���=�Ȟ?f^mq��ƀ�3\�^yH�� ����9 �-:�Fo��E��*���R��@7�uPb���

��i��6�=�
��G�x�!�S����_sq�'@Q@�	��Mj�ua�����q�(�!FkE���M�^�VƐ�ץgʸ=��[)��5����b����� Vp?[[OI���H���όؗh���ۭ�؞��ɽm�������&�'��B�#�0�D�
\2b͇�"��XrE��_^�{s�Q�e�������G��0�
1 D�!|��Y�F?�0e���{��ް£L�r�IU��d+Оt! g��!�dO7$?E>��-e689f�+��G%R�4*�`���N�W�~��f�%�?�&�Ǆ�f�u������Y��@)v#.�fB���J�X?*��{����X�ɢQ뙼	�����źK{�(/�P��{#�=�6H�����:�"�Q����KJiKc�6��So侳��m�u�ڰ,-԰硲��_����۳fY��3�p � ���Տ��
m����_�*V��.f�Т�`m�N�d���n)z='���h�R�l[���5�T�K�p�Z��R�V�XDV��ny� s���l*�?]L����Ѹo]d�i���HY�ky[�5�8�"�kv��L�=9zy%'�V���-[�S��r�[� ��PA�Lկ%�Y��;%0��`�!�r���8�Ka���T��)�lI:�����$�?	!�NZ`�,S54����>*o��S�� �o!��O�w[l�6�OD<�ޙ�,��u5��Kh� S��������LN��vw)#V&�dU����"�bP����w����m��&��/���;�x���4�8�Uc��y��^�5�@������<����%�.��@̉�	Oc�sr�K���7�z�/���"|��y#��5�
۴��CS���1������A�t��6qO�K����B8wX�v��u���M:����*x�Cы*�n��!�s��Z��Y���2�ى��2�Xr�O��8Q����Tf� �N�B0^qu8�a�Zf&K�}2c,�Cl����Z�9��۸7�MU4��}??������(҆�Ow��W�]m�C��f�(�/aZJ���<�VD�ħM,{���=�:&�(���CS�	���p��K�̚�0N���J��#'�
�3I��L���m�T�ڔc�`�a7��@JD����D�蠸pq�mL�:B ���A��QB[k�xSøA��z�bg��LPqt�r��6:�K����_���F���Ѩ |i���m�Gn�PY�o��Y܁^ܒ���Y$V�dzk�[��_P�&�a��D�5A�ۧ�b=� ���ٔBs&�NO�?�Dn���yw'�D���{R|�[,"�#�s�]��`KE����t��7��=b��b�>�dւ����2ZN�}�Xİ����¼8�ⵏ���w(�`���5W{�<�HЮj�i֍�>�q���1��V��x�$`��!AbW_A�O�����Ȯ$� �p����:�J(3��&�g#�7����Qy�O��韙6���s��1M�[�ٔ� ~�6�Ӽn4�V����W��/�#��yq~n�P2߆�54�`M�V���x��n� k�Y�̘��Y��XN]Q��;ܩ��J��4J��Z��5���t����<�$���@�\��<���y�u���Fn_��jh��UB&��g�UG^�X�3��{�|��Fs���m���۞.��	A�ΐP8+�K����d;�`@\����
¯C:��62�~�>UwF)�C,fY�d+��v�?(|����x}�am��}-�o΂W���.�aG(Ҥ͖�ŉ�O�}(��i�}�7)!����#����N��1�����C��1�w*���o.��[�,v�����2QO���}��*�B,y�H{/�L�1}���|��>��6-��w��mG���z�칝��.[l=�~�
��U3�v�ZWIKj��u�L>'�i����l�0�g��+
}o<���<9]�Nˑt��R�����B#$)wÜԺ1�(b󿊥��_4Rѵ�0~�ѻ=b���)�W�L������,K^��J ��; VV�������`�J~����Fx�m��|'Ѱ$�N�S���_MLb
l�2��
��G�">-��s3VH+W��w��ߐ��>JPډi�"ꊰ��ˠh�}^g'�w�y�u�h�o�{TU�<]�����[�U�ѰX(�;�I��LV忢�zE4��~a-?.Ĥ��VW+��S�';����ɚ����ծ2;��U� ;��g��ąv����:��{�l�>���ՙ��]-�#��ӗ�*�\b���;�Djiظ�2{X&��5W&��K��><|m��U=yY�3Ƌ<���N��Ϭ1�ο��v?\��P�ΰ�j��a�-�%����{ԗ!]Ls��3�0��.�|�W�����zBq(��>��ݡ��"wq��"���c�['���%���KD)1(0%a�]�p�犵l�vY�$\����{­,����ÂZ���-`�����R�^�j����ڟy�iﵫ����_/����se�8LuwW���t�'&��RH�O5#��*��Y<��y�"�IZ�*)Q�(����T��8��w���"�:�Q`Uީ�=L�G�� �����
�!�^^��V;`�D���Un�g�����5�Jk�EK�J��-"k+���7�&�� m���K)�! P�~R>��]4}a��^�B��$LE:��[��z[�|b�A;� �a���&c3ח"�BWX}�>ӉT�SCU�e�K���w~v1�68��kSs%�$(P:�����ѥ0};4qC���(���7�ۓW����EoY���E�\�#:�%n
8₱�h�nԓ5�}�ln�`�X#K��0�0D�n TP���a�gȂS���� ��������\i1����byH,8���ԫ�%;�p��:+(����к����)��y�P��Vj*��`0jo�(F�a�¤���?�O�� Q�o�@����%���Ӽ��i՚�ږ@���GƲ�>W���,���7��i� !g���Y��O/��mF��W��QU���L�r"�>�u��%���wXj�����gi.���r �5�4"mF�B�	���9�ū�(����6g3�gܒ�68��	.TF��`1����V���/2}���Le��hT�u��
(���ܼ0���:�L���TW6*��(
k�ՙ{�����ܩ�rHisW����h�g�����v��g��/�:�)u��;)���Yޜr7��ˬ���1���"&�0������+ܙ�Ö�w�b��q-Wɠ�rA���3(�m��0�Grgݴբ>�A�1�@��� ��p�z�1�6b�Tx�k�벜���5g�;���U��A@j�p�4�Ql�^��7�I���)8���T�!�=����
'zÃx��?�-6�a�⽀S����O�iY��7�][l�ؘ!'KYE������UߵA�3�s����L�~M�bF,dj���ײ�b,��f/:���9�#Q��K�G���Kp�*<@
��J�����y:��u1�x]Q��#g*ؔ�� 2�"g<Y[A���SJn�LLsF��QT.���%s�RJv�O1��pYt-�t�N!���YT�����E��l�9nf\�:P�������7-z�"������<�0���t;�[����s�?�����<��O4K\��E��(�^W����M�]�Fx,���k���9$��j�3>�Q?�gl׍�;^J�рc��^(����ѣc��ꐳ�鷄�)���?3ƒ�u��xj�� ��A�ukD2V�r�fWf��F��v�C~ �`�"�I<٢��F/i���]���c-�$���iؤ����ۂ/6ޯ���\˺I�� ��:O����Q3��|e��k&91<���˕�`��iE��2�����a��<� `�tL=�q�-=��ũ�L��3g��}�~�h,�b�w7W��7%o3�2r��
t�-�?G�� 6�-�[��}��e=FoOSe�����@y����ۑrJ-Re%6��n��fg��%���e�]�����*�\F��w����׳	�޻/b���������J�랗ʹ�����h�|���Z�yg��4E��1�Q��*��t�dK��޶��1~u��'!�-FV���`Ta���&�����s(�17�\^/І��� ����K^�g.rGTOD�> G��xh;�A/y->&�x��:�R��~	�lr��3���v/�b�A ��d-UX�9� d#ܥ�Ϙ$�:i�� ��;R8��g�w�M��Y�ec�)GA�IB���#N����3��r�OK��Ǒ���r^��ơT0β~hLڒ֔���U�U�*�#��!ǀ��Gz �`��Z[��7�l] ���Jo��\��eo���8��Н��Ś/vq�CKaͶ�vf���1m&�]O�c�7�x�7˹�WAu� ܜr:�=�}ߙ�8<�-�:����B�-i9*��%�>ˆpƇ���Ү�mQ�i�L�:w�"��V&PU,�V ���p������ 9)������-
[���j-'���	�-����DM����`C��j�r/�q-��"�Gl�QM��ZZZ}#�URY�J6�Y����8���qIU���)�Hi���9���=g&�C�>0z%�u�R1�ĳq�}?�WE�ˠ�����|���mk��
�~�w����'��#'�{���X<,3Εp)ZBC7}�^X�EC�����%�Z�U�������.3��z7��K7�!7�a�~2�s�a9��������*m��R�N��ӱ;t��Kזe鑿����Ցe�6�塸`ԨP����	t��}�iLU��U,ԍ�����f�7��>�Δ���/	�l(�x:{��R��C�y{�|��D��ns=z�Ɯ.���ɑ�4|�UP�e}@w�#[p�.�����\ �e�
c�R�j�����{�L�j�
�۲<��K@�n~��xM&��Cg+��ڶ������(�j��vm���t%e��U�(S��=c�BU"�Bl*(Y�����GV��4Q"�:�<6���]�#�BAwŨim�4XӾd<7����(�K�uq&hR�ej��A����\�j��gbw;K�>�gs��ӌ�o!��vaZ�W�>�\t�з[���[񥔗@r&fu��L �Z�{����d��M��XcӨP�- ^��������)7H/�$=<f���@��h 7k��k�	��U�0���.��ٟҪ�8�E�5r_�����b�[��kwk{,�≧�]��g�3��t�v�2�#���$|�q.al�iF&"G�[,�C1�2�U��U<L`͉ω�ý�����2z'�E�nV��L�Zee�q���8>B1At�������[z���t�p:*���C��\�k���z#r<"��ǘw����<�WP4$^|\��{V�a�@�K/�Ox�(�J��;VwfmCZ����z�K�{�V�P�ܯq���Xvr�����_c���&3®S������C��W�3]B��YJ
H��l腡��?=��X�ٚ��5��o�gpl� ���C?��l˫��̈́s�N��:��u��ތ/�V��&Wʫo��Mu����
��1�c�1`�ީ�8��|��w���y����:��mv{�� Μn�St¼e*F�Aǀ��=��;w��@��lU�
BL_4�|c����^|�󊚃��%{�
d�no�/��QcQtW���P��ʘ�9��^���`OM@����{��b�Í��0j�xb���*�������|��c���I�eG� �r{{�u �l9G�3���܌6���o�n��r���� 8uo6T �vk��ttWLA��8��LtC�pJ����R���y:4�7t!e���n�x[�Z^��u�,����ť%U������#�̕��	:N�K�;��MN�]jRu�W����҈|Q��֚�̴��$)�Q�`"��+~���{�"�����Z�$�,�2�M�.�h[���l���Z+��y,��3���WA�[��;Ķ��鱁5��C����N�^!K}���$�S�+$d	@�v�$p��7L�b�Q�������.L�v�6�J�%�N
z*؝�4)�XI[�~��3�i��e�J<:��f�t�h�.R?�^�,�Wy_�aZ���ݲcᆶ�HU+���s����0My#Msz���2H�u7�A5K�㭵o鴦b��ds
:�"~eo$�n�#�hh��.b��E��G��º\���8y��8�
��{mdwg��j���.g��v�$��`��] 5G��Q6�x� .�b
�!�d�~ݧ»�!L9,�N$�M�2�L	�:���QƟ0��ɬ��z	ģqd�^�R�B���>G-9V##�\�1�g֓�4�'�;Õ6�5̄��=�[S@��Y+��yJ#C4@L��K�{��dW��ŉ�����;�"5=�*���J�[���Q�XT�x��jG����#̓�HL��}�� �*�l`��Z��GgƋ��ح�{���<`��u�nb�-�$��~�lɲ���C�Ĥ��DI.�G��
�1�gNH���j�.au�~a�S���W�iY�b6�5�}(Y�������*6���E��.ٰ�.���0yK�*H����n��+gI
�ͧF���3���j2�Q��yô4�=���&F��m�UVk�~M���r����4�t����ɋv��&ƅ-kb b��$q�V�<� 7�ZQ�_1���ʳ���BOed�Z�5=�Y28�묫���t-�~Wg�m7��-'�w���zX�O���HڽJ�'3�����8��m���o~k.�	:��X%�&����̎8�nh�/���`��@nS9�S�|�]>�)��j,�͛��8o`�7���ILM$z��1��"`櫗�4�_=�es���y����R�ՐrV�m��1P�oRh�=`د�B���1����~�֨�����z��ǩ�|L�R8V5XY�[�/�㥏@�g\w LwmA���[[3������54��6�2%�
�Cm��d�/^>��+�۷�!O�Bf~�:D#yy��.�=6����%e�������`�za�oZu�)$/8Y�mn�=���Qp/UK�@W>!9��t����
�W��x.��w?�Y�'t�%|�X�F �����]�s,�;:�2rv������1E�ؐ�Vq�?�ԲA�n n�qق��vy�bl�Uz�}��H�C����\	�U��p[:C���Y)
��j��}��i�²+KW�P�I��MJ���u�B�E3FD-7=�7K8���r�O�M��5[��e�Xb�s�7��ؗ�m"��tM�n���2�ѣ��B��^�_��|�cO�cS�m�-�&ZbSʵ�#��fAmj��61���?2nȄ��M^���t���.]z�vş&K��ںd`Zs�d�&�?��6܅҉L���/4|eJ�FU�6����`հ���d�3�ʣKO
Θ�Ș�y$�@_�"�.<'�u �X (z�#̏�<���Q��|�9�-� �H�o�-��C��������0鵓Rh��7?[7�'�2b$W���Q*��i��
Uu.��{��|0L�����Y��0��H�f�5�$<-в��4	�ͪ����n��c5��Z��T�}'���A�T�[����y
�N4����FhB��S�^�
� wu흐 �by���NX�W��Tܚk��r�\$q~�7���V�����aSKAe~a�} �3�rE��.5�) S��ۦ���0�q��G�5���#o���'Vs�i���78\���D��6>8�
1��_a ����W2
��`�6�Sp�ʪcf�g��`p�M6+����&���2ʟ.dl'>0!fH���f߼\G�}����:���݈��C�'K�N����S�jNs���7�&�џhˊ�T��dK]e�f�L�:�9ַ\��*k�I�Sj~�ⲧt�>�A�/T��31!ԋ�nF^Y�0�NC����9v\��]��(9��urOL<߆Zͅ��^ZHMBz
ˀ�'l�B�0�����$[��,���R�^���W	I����v�,�̏,'�z���ݓ7lǕ@qɁ��B��ǈpC���u�1w!����_��2g-	��������܌rlÎ0;��l��Pv
T�5��_Xu�+�W4��&=[h��߯v��N��؈�8s���9P�Js i����}ͳ�޳Zِ%��fm�˽�o�!�vh#M�t(����������1�>%p��y8��4��2�O���JiE_���K�[�>��,�/����n/Tm��,o?�{�b0�'�(%�͏������7r)��Q�iТ��	�$<Nn��eæX�}�y|�:C1F5*�+������d�kW[`t�+Xe������U�3
oF.�0�> �f��M�k�+iz��A����=�<��ɐ+��iW�����{l����:�AQ~N�J
4� b�?��I^�5k~�i[�� ��ZPfNJ`v)<GXWQk��\��˴�,�e�I��+0Oc���4��=kgr���¨�
��C,����|��F�>ω�y"��/�X�!V�!�c3C���t);-�7��6K9�������k��?��w��_�^��紦�lh���Q��d������F`d��@�>2SdKpNJL��_�}�1�v�23������5�.�#Z��@�yz&�uxV�2����(;�r�	*D�U�wt ���+��=e; h�$��@��ׁ�c�fq�
�!|��[zRh�'E�+O�;���y�b�U����|���?�����S8o�SYE��<1��,��r�,C,� �sH.	V�%��e4y|tQ�S��_��n���Y���UKy��zl���Y���r׷��[��tp�s�m��6y�O�^�4D �����Ю�zNѩ�;Ǥ"=���9V��>Dژ{�?]r�צebKKbV�����k_����֯XK�=�]�������$`N�@��iV6�X�������vjq��&���B�+�<+��o��I��ցY;���][Һ��Cq�_�ʻ0iN�p<\�����g*|V�� 1�'�%��\*AA��J�����!�w�"7�Ģ�����4�ק%%�j��< ��̦sqR��9+��d؋kM3�!J-=(<Y�e9�������체�����/ق�x�KVF�U������Ǒ��cz��gO��KG*�h�}8�w�ǑRi�EVwQ��t���jƻ�	[�O�.��mn ?�kxî?�|0q}�)˳�W�Y����ďJM�+`�<t$��J��� ��?���ѰQ�Q38x�Ws:0&.+�}�8X�	'��	�����KD#Wo1F�sy�GD{[����tu͑+0?��|�� ��L]�ܝ���kE�^��d���R�����;N<�!��A���}+�@�V�Iӂ`���byİ�٪���/_��5���.X�����l������p��Q�$���e��u5��Zyú+\Add�C�ڊI�F��#���v��4sL� ���`+�'u�m�����OV�O8����	Ń)��ˡO��ړ��V] z+p&���27z�,�A��G�d�d=@�*�F�
dY
�f�����-��&�)r}�vD�����ݟ���+�����L0Rw�q�M�!� ��h�֬�x<t��ɐ_z%A�b�k;��\�|s��M�+Md-�1�] ����� �З����A��&�I�2��A��i��8��S^;Ͼ�`��byq��8�4�]-���"enQzm����`Z_	�in�֛E?��vg��ަ]��M>U�S�2,0����ji��L�-;9��!9���Z5�|`.�j�H�Ft0��~�`A�J�}�ߵ�ǯ������I��OG^OM�s�]@ �UR����p���iX�0K��	���FQ"�1I1$����5D]��m�vD��)_��VY��g����| �^J�x|�Bȟ��+pz��3B9/�{_�|[��o.8Ŵtɤ-`g ��WZ��X�a�����Q�^˃�o�j���� ��J�[�VB .eF��R���d����ޣ����r+���i��5U��a��~�W��
Vk?(�LR�i[�2�l���95�>�o9�г�>�o��&�a�mt�pM5jo��Cqt7�$:��[�\˴�����E��#��j~�$�R_Ջ����eǤZ����9��X�5�l�Z��^u��*FS�^Wm9�6�C����@�~S����D%$�~�1�p�������9�} ��9L�{�bX��?T�Y������k�@P����?;��n���7㺬��L��V�o?p?R���0�s���gٽܨV�24�{ �<�I㢼��ο�Ŵ!���M�$Eŏ�Y������94a�G���G-h߄8�2ծ� c�C��)��	��)�a}zD<��2�_Ħi�gљ���6O�í)+�T�H�q�uA��<��!�����և�
��;����%r	����m�$25�^�a�+��@�KS�P�eKv�L�@X 8[�/RH���4���v�e;TUd�������,tfP+�אS�2�cE�b7����]���xϔvQ��7��0���W�i�BH��(Ab=�H���1�)qᤵ��_�pUQ����g0}~)��G}��AhE�J�|3�^@6?�1Nq8D��Kȧ�ӿxh@����K�y̞<F+�I�:j�g@���*㓤�B��v�臹��@�]��!+џ@�q1����}ƙ\��:�K$�1�B�̏�4/Vn�}��n���%��(�-��=��9�lBn���d�pD�2d�"֨�;�	����&�3ڔ� ���5�.p�
и�	�̽2c�ݖ��Pw=���X9����הB��J�� ɧϜ�P��4���%��BJ�u��7�_F�YB7W�/h=�mmՑ�[�����\*Zϣ�Wd�\ùe^���6�������t�6e�նKfQ��TUGFߖ����^�Q��a��������g�<��F����a���0�*�ĸ����V��;�L�5l�t�� �\Zָ���|�����'ƙVa�_��wH!��li�����x�'�/cJ9� �����ԩ�:,C��o��u�&M�{����6�
��!Fu�.Љ�
2��H��ؾ��M�%���;����X��X��z�L#����k����u[}$�pKe��oIv�C=f�&�c���ǨR N����y�������f2ܳ?�����a��~�>�ڶ���bQv� ���3�����_2z[��4c|�ʐ�qԀd�Y��1͸�)sI6�5�2V,�j�4��[	�6����Rɠ�A��h����`'d��jg/�N��ja� ���dD�4~#����|�������b���A�~�b�ci�6OԺs�4
 T�KT���PHq�3\��Zhĕ��x7����ezl6e����sT�Z�xߋe��"�ڈs� I�T�����gZ�� �"�^	�q��e{3������W��Z��^��v��`��(}{�ufRN�e���$�?��t�Lg������m�p.�&�0�e���m�C���?w �2�>����`�4)y9M�F�ꆏ���	[^Py����D4Ҍ��hn4�m��1�G�k�!��Hp�V�af�h=!w/�t�����\��g���/%�V}��z��O�ƻ����p�,���4+��;��|v�ծa�E��P\s�����Z�͉�t��[?��,w�j��<T�<<+]I�) ��@�;��Ƹ��n?��(
�,aE!�������GKb=�V.���.yB�ӳۜc��%�?|��0s���7M��&�7E�8Kr �T�ʹ�4���0,�[�"9�I�Z��'�G�$�;z<�!��8]Di�HN�q*�q���P��e����^��b9������R��
I4p������TE$�����-`z�J����[J"J�@v���WA��0?I�xf�f]�Du�������N��`� GںMk�Ԧ{9@����QD�px�顲���k;y��6���3�e���+$SA���J��t����Z�c3�G�=�{�"��e��ԓm!�nQ�#��u�������p֊�����^��� 9��W;�/�bj`��0g��}��<��ml9`����,wE~VS�\�"	�I�ʆ��]�]4�cRy�b�)uE�5�z��p҆2��8|�SD4�z饥ߍ�mߒ8��n�̹���ǐҎ��vm��zeA�._��ߟ^\f'�MG&�ܪ]�����0B^��Mާ0u$5�%t�1v�8�_$\+{�8Dwt�C���	 ����?!���C*�n!�W�7�m�F�ՙ�T�E�7�1��5����T��,�+���R��#Q}f��<��K
k���vʭܞU��Gt�:xJ��{|�L�9i�+��6"�y5�WӼ@�X� ���"����L̓�s/FL�:A��R���D��_�^z�'�d���S|���pw]�0�au�uTC"O߶춢|��{ע$����˓Z�}�j8吿?�w����詄��gƣàtm�&b~d�ɓK�9�) ��5	P��������������@�Ye䋑7���r-<uF��8��y�W|��1�^G����Ʉf��=@�����eD+e�+�g�-��/-,�$�ר�90�O�[��;�f\8�0�׀Z��c1��ެ��cY�fS���������	@ZԵM\?)��� �������<����,�"��Ϊ2C��eh]z��wOCȜ��΋f��]>���Л��(������OeL���$�ݱ5lQ��w�KR~��&fɘ�����\EaG(uV$E��JLfe�?.q�R"$-�����g��ab��� <8E:��U��ѣ;0�ĵK� �K�a8\ì�Q�������t?Q�s`D+��F�C���h�gaD$8_���tѭk?ى����G4�	[��w�6~;,H��'>�)c�xd�d:�]��
�;+k���|YA� �_%4�!U?�2
�z5^��#R�=���ܰk1�.�wz먧%�*�*͓���#k������&��K*Z/�7m�o�*�D�k(�nge���5�CA?��"�P�Ų>���ܺ��$�d�|H%P���
&�����R���zhSB��}-Buٔ�u�f�˓�m 0�ʏö�M!UN�K�%/T>d��J�!(�ht��g4��n�ǔn�0Kqq(x�D���n��o?��&e�� �nlM�+
r;��O���x��X�֯dUP�,#��6��^i�}�Wڷ��ϵ�2w%�X~�\�K䏥�x��Cx�޻D1��/B��v��	��+`h�����gR�; ��6�`i�����(�c���.�ԅlg;TiMV��7«�]q��|�]Zm��H�3�1ԋ��.B�\��JO��?n�6ߎ]�qP��#.s��̾�Ğ7g|�2i����e�����M!}L�&!�D=C����7�t�\,��n CW2XTo��i:���Xg�bK��餼u�u����
2�N�s=�;�gƺ�P�r*�٥#�����2gT0����dYם<J�\�QL�0�%�q,���\T��8��R��vD����y�~2�1苂��:#z\�r�:�Ol%�t�uB���m�mZ�S^G��������M�)�Ϊ�2q�Yk�-���F�g����g�U%�ß���)���:�;��T��GҢ)���\�ϩQ5N�O9�r6��M,�	�*�����d�dd�(�?����f
u:&Z�w���43^�K�q�r3rn��Ïm �.����p�y��� )�~dz�:����<�߱/��쑜p��`�}Z���u�pu�x�(����/e9#�������������ml<:p!�P:�&�gg�C�'L�M%��e$����ڟ�w�0.6I�|�,"��Q��������*j1ZzJi��0t�"����>�K�B����ލ���^)~pl�Lyg����ᗿ��)�Ĳ�lud|Qܚ��RT�u,wɀ� -��|��8�-�dH��톿e^�? -H�$�j�`�E�N��@���� �ө�f�B��g�s���Z>��ѽ>OG�j��ŭ��?O�쇪�]�Kbsv?)�o����*�c�屍�?`��毒;w��v���'��y���~�1�(1WX����f��(s3@ދ�� �U�Ǝ�G).�D^6?�GLF�yڨ��3���rIݘ'5��"u~߶D���`�E����Mr�V T>Qsry��Ru�������Ott�����ٸ��*;H[����1��u���8�����nbQ{Ԝװ��4�2��.�OI�۰�,L����T�ذ������л�[<��h��2�^�z2<T��Is��P����Nկj$e�{�H8^������qB݂��K5��ir>��2J��5�;������@��T���pe4VE�U������Rh�V��=.�Βo�۠� �*t�ة n-�T;r����$��!����s�|Ћ��d��z�:UH�F�vlU��_���t1�)��X^�q�hȢ�>�)�)և�2H��[m��Hx�
OH��z�a��N����@�j?�,�֦�.�n���vv�T�l?#�8��P\~��R�<�����wO�ws7\�#8�P/�=i�ǭ�F+�BI �Z`�wG� %�V�Mj1���-Ӽftnǘټo�R��\h&�>i�d�Nc���E�O� ep���C��{�6��[�E��&�ԕ��٧�Y�,h��asd%d��u��B����;ZªH0���R�����aE�B��E��+���l�ƫ������Gz��p�e�m�V�f{.%	x��;���.[���:��,4!��k�H}�$��l���;��F-Yk�t�<���xH��Tს�q4�89��ؽ��#<:xt�3�^h$!Z6�,�c�Ł��^BKbӒ�q��d9����G�IGe�%V�2܆��H6�M���+��x�-��-����+$d��F�86B�O�ջ�j����o�9巃9�틁	��xP�.9����._��8
jr��p7 ���^��T�"{9?+���=���͟�M�G�<�����KS4m��t+_g��-W��	�%�~�O�&*�Χ;���?�t\&��z�0[}c�Na,/���/��"s��uP~�3�������������(Zdo��I�7,�߇��}��>�ۻ�(
ogJ��k<�>a�g�p�lP�sJ�� �՟��3���c���Q��Զ���80��R�'��Uջ&(�����������dD��WT������00����HC`��S���;�s!Caj�.��'Т8"�Fڗ�7l��c�qM�1� 9B��~��%���WK������']�w�A��W�hӯB��Ϡ�'�&��?lA����9��a��$��7�kCA��;�k/[���A��[�w>û��Z�;��/,�y�C%�I	v ��������gw*��ệ�n��=(�*���r4���;�d��<�7)��Go�\�l�ؑ}i��/���7`�cM��E���!�cb^�Ǩ�:�b3%�4^S.V4Q7�y��lW.A����{�eĤ#��=��DlC�a�I�0�~oN\ЖKn�ټ+j����&``��S�Iz�X�;S��'�8�>�!O�=P���FV��A��]�9L��z�k���ݳg�:�|]wD|+�������e�R\�������ԸD�K�,0�n���:�2�.��y�aؓ%ps�a�P�
^�ơY��?�TQ@0�9�ش�@7:�SMhV�[N���u�3H.�8d�u=9�]�P���<�1�AjZ��G���x��@��ɵ�)���|�O�:�PY�)�X��7���4�~C���v���ͩI~H�%5��D�-���c�©+�"�$�R��J[�--s1P�Y+fk�w��='=�/2ڜ��iوn��Qy^��Ut�
V�p%Ux���9���g���Z��?b��e��U��
��JD��H���˥Ηvk�<� e ޏ�;�K���5�O^����k�n�+>&Xow�R$ZSRb�D��b�*V@�V����o\Z7��E�^�_���G�l��#L���p�hL�{�9\�#ן?Mw����*0��Ϫ(�9i������}�%��O˙�{���i��aW�ՓX!vи�g`��F�}�8�k&���$X�;��ݖ:S�B4�/��[���;!���=�g���8ZI�v�w��F��;'�GY[��s@L���2_����+��@�n��<��6WTBJ��;!����"N~�Տ(�z��Àd�n�n�vp��ǅ
�&K,Rj�[:��Sh���3�jtI��+�V]!6�jː�`C��'T�n+��rHqWJ�⤷�R[JځGp�Kc%DL4L�H^[�+���z��"8�p�2���..x�|[�/9�b�:�_G�RXm����>�J;�b�e��[�����P*��5�8Yɏ�0=ݑh��)����<�v�w36��X��w1��܂��oS��x/�H�U
��&�nx�R��$��n#����o��ͣ�P��L�J��[/�,d�R�Rq���Ң�`�=3��9�)��F^��v0���J��F�RW��3�p�����|.г~��5�O�pƈ6G$�X�^$#�t�D����X��$�-���@�_'�{�E^�Y�����-�"̗�)���uf�b38E�V��h�O�,S�����`�8��UE����/@�i&��`:F�]�h�Z6Q��X�����B�����+D�z\}���M䓶MLNI�}��,&^�o�n����Od�ރ�]�H����T�)�!S�E��,x�Yjg>R�ȃ����'P^"ċ��B.�յ�/����h�Dq�%�5���OC��Nx����6��-H��]�K�F{ݠ�Q"�J-V]Ӱ)�#.UwC�y��<���i�c�Ya�Rѭ���� ��"3Ms���\��U�?�)�SQˑ��ͨ~� �}���١-��ð�5	��:o��x}NoE��v�k�*��㟜$��q��D@r�\��-����Sd$ �r	U����Y�����Uh��iPtVv`ab��w��y������ѧ�)i�\�3Vf<����l�����b��KW�g�@p	�	%������� ��Y�"܅���+��sf��5�����j|�s�����}�Rש�t�i�PVү|s9aS���N�]AS�9�v�a99je�W��1����������n���>d������A܇��؈+̜����� �m��K�Ǩ5����� �8T���U1؃3�������):����$��0�Mӟ�z�_rB\��{
�ˇ��(��1]�v��w��(�yY�m�C�츎�/\HԗO���!!G���P<䅊ڶ`�� @(�翭�@�#HoM?��	�����{&��<Lq�W�Y��r-��b(�$"a��U��~��'����\���%�Mڭ�?C�N���d;�j�)<:(����O��e<���n�K,��O�ޏg����ڍ�wFn�ī��<9�ܶf4N�
��U�rc�k0�]���p!�/�S�}�!������~�� X�d��O��K�*+0���vxշyf�+��1.� �b�Y��9��Z��K��bO�p!/����:�O�S^c�%^.;�s�� K[��|K_��B�Zt�[��$����r[�D@{�::�A#(g��&�JnO�wh�C�{�k�,I��\�;~��p�ڛo�ř����t|��喥t�����rZ3?ҬH���ϫ�e�?�	oI�U��D�ݛ�5�5�b��;�����n��̾I���1�H!������t���&t�qzOy�,kb|�ԡ�dp��ad f3�V��k�,�Kv����IzD�n�0 �IB��\!�RP]�
����FeK�S��ľ����>�d���F��J�����@����%��Mf)*iPy��(C�I�0wͼ�Q>Z�޴���6,%��:Zܿ�i[��o��������&����~5̎\}���8t6CH��]i����| ��䧬�*�K}�ڀ5\�(��<�迍��� H{o0�X�윉�n�b#�+�r�!l@#�L�)^�p%��k@�2Q�]���,r8C�<�tw\�����m%���L?<��4/N���\�
���D!�R��
�0��㺬K��!��a�v@e�n�!��OG��+��@�a�#8�F�a��t���޻P���h
�M���Q�S�_�k�)�d��O�;0�n	w�0�F燘�[7�%�H��8ĠmM ��B�-iL2��Q�d����C����5_��VhX�|�w�Wu���Q�N�S���+�=�`W8�w���)��g���D	���͐d�mW��Z�N�I��u����(����w����qΓ�fN�} <.}����m�%�R,�$�ȑO�̠���}e\����la�K	�������e�6{xlaAR��̉�M��NE� ��P�F��l�,ـܙ�d�"�a��%2T��@�t�t���[�v!~,�*q��B�����;� ,��+!x�[�0F�~^w�..	-wB9����LT����r��!�dl�*zpk�mPVLńo��o�fZ��S1&@�|�h�DX�ӒG �-��r�DpbIjX{@���P�vA�d�{K��/á����Q-h��W��1]�3� HJ�~�T�T`��~�:�An1	@s��vo��"�И�x$��H�a*���bIu�v4 ��-��ȁ��� U�E��~l�g�)��'�K�w���,��N�tcKWb魙���]I{|�0PJ��_J��ҊԊW�;^3�*}4 U�_ƈD}�dv7ދ����+a���U�����������h�f�G�oC�k��J=Gxx�.��/z�g�B��� �=�,"1�/�=�+�c��)�B�|~���҅{%s,�,}#�@��[���N��C���x[1���z|b��a)�:�X�0�r�ƭ��#r��+�.�]#0��;��Ca7��
�x-�}y�X2W�����K��I� �W�r-<X�!{�_��ԼTܳ�����-r�wS�/�ft�ucӫN^�{����ܚ�]�+|4�}��kײC�IǛ�"xD�s�uQ&]��s�th��к�g>@��G��A�w�����N!!i��:�o����oZ8߂I��u�B4}�*�jl�]\�������6ؙ������RU(na=|L�С=�\��-8]UK8=)^��'F�S���aD��XV�i�Yҏ�Sk�$���W�]h=�h�~��K�@�(+�����&��׍Z[C���=��RY���/pfk#W�$߶,ӤUZo9GF� ��I�ϕ��H<=�Z?�d��� ��l��ɾ���{��B|1�{�0�g�����!ݚ`n��)��ѵB�UZ��ȋ�����su��yۼ�Xy��Q�3���'�]�����d3#��X.�u�e���H���Q�W��~���>�xs2[� d3S�2"�V��_�4^ͽ1X��?U��}���J��;-
���u��E&�B4��7^�ŕ'^:eՍ
�� �f-���2��>���G��@ەZՆ��jB-RR�1�!�^����upҘP�[�!�L��>�^�sI���I׏ǘ#����X2�* ;c������U�/���x���i�2�Kp|a�(Sl��ܩQ{��S�RИ�`��Ԃ�y�at�� �� ��f_`d�"��ed���@ik/��.�z!8������&�Έ@�RGҽ�(���+-Q�������{.M�R�ddq���~u�A�b�U&v�
���A桹3�6�``^з�%��g���Q�􉍿�D(~>��-FI$d�H�u���誷^ycĚ��d��39�����,Y�-�.q
��Mi���vX�@;�J�_@��F"��c������K�M);Y�<�nv+��X���+�([�\���� ����hQ����\���d�������<��¥k����'{�1��K�D�~i��#�Jd�$���c����^2����iƺ_�ʽ��J�yX(�Z���b32O�Qq��;��q�D�2+4�I8��zxSmCtj8����/��TCfa؂@���M�Q��K�-v����}��y�fc�=:E�{	Ѐj�8ST���S��{ϯ�) ��4��s���ʲ�CrCqmX��P�7r�K^Mj�o^����0э�^H�s@��]�{���:�Ŭ�hL��T�`��59�t"�� ��O�pp%�j��c}[}t��{@�	���.y�-�&�p�y�P#�!�4O�~t�EJb44��jNaD�O|SlI�u�q5�:��cҝ��e��a�I4�$bHZ��d@�V����J���Ժݖ�V%߃l��K�#��K�c����������9W����vQtӚv�]��*�68���)�NNc��ߤ@���֧
��\� �g�"��T���]���*��E9d�� ��~������:r�H����c�8N�İ��0ڠ	Ftq�dGG��q���Y�k�h\��n}!�i@�9�e��w��[r���W�~c�fB&�`ڴf�sъ����@���ڊ�i�CyPS(�u4ŷ;�~��]�H��;�Y�YgP�^ ��ΦD�� ��<��eU�t!���Cƹ��}	8�=�~��|;Z��u8�30ɶ��k�ؙ�Ra��w�}�M������Ͼ��u��Uٸ�X�V���F������#�t>���Г0�Y�9UQ{V�gp�660ڧ_�Ȩ	����^���Y�@y~Ȯ ��	�z�!��shA孑��;]enW�ܼ<�Mͩ�i}�����OAC����	�&_����ҕ�E+�A��%}�,��'�f��_�i掋$cұQD�`�����kNC��Ŵ<V�����FD�[�VI��|�5�$.(�2�%CY�W�mZ
e���R�UPDסq��eK�M!�4��\�:]l����į�}k�Z�b�=wqKb-�XQ�Z!�|�l���:>%/� Gy4��Ս.�@����E��6��OҹF������c�[]����Ds�U!�}��(58ף�ȹh+M.�߭��|9W�H�����
�3���T�$���ɞ�G	�!_p�����R9M�	�azU�x���ޘ�'2^���|gJ����T�uu�r׭�N�f�,��/�+Il&�j�����ɑN5�܇����j9��;���(^�^�07̝1�_Z[��Z#���g`��R��eK�}�#F !��b��%K�,�.g����;n��S�-fJW��g����v��#�����;�����k64U�A�l}���9騸�����AYS�sY#�=�S�e9Ԏi�;z��}'P5�6fsZ*�d��z ����^b]�]C/��Vc�PRP�8�V�U>�D9���=��+J}�[Ԙ��~F,�T��B��ۼR���e9�[�T�E��<����)��H�7!H��bPݏ{��,ߏ���}>�D�[��]�^=�W��r����Np�	�i>'^C��|�Ϭ��ܯ�Y~�υ�8��+���j�I����W�:g��F����&�7�u���fi�eKݼ*o�4�H�6�K�̌&j��-�q&%7}���n�l���ڽVzN[��"~uc�ʲ4�p���⑼Z��@�b|)l���N�Pi6V�s�����R�̘���c���r��7��8<��G��O���IQY@O)�žY"_�k�˸q}�-��6D_A%��!�&�ΌO�H+�l�	�hK�fx�� 60}��M���@b���_O��.�'i5�c��F�K2 ;��4{#�k%�đ���ҩ��&��5���0Qǥ�μhe�#%U���R\�Y��hҹ0 ez��K�D%��� V�,�)�ɛf[E��Z�H�)�Sz�V�i+B���5��,��{ ��wC�oDp�,�b�`�(��� �)|��bF|W)���Wz�пE�_��՚�)��>?�mH�59���q; ��!���h/�$�/b�-Ԫ�h�x�l1;aO���C��i��.c�B(�И�Y�ov�A��F"ap�����&iѨ��ŵ�%�f4�Yz���2�_��t�AC��R��	�ӒM�Z�8o�[�=��\��j68{Xj��Z�0P�<��Q� %��-�GSBJ��Q,p�ՠ�~��Y6)'�c�O��I�<��������.�*��<����;�&h��a6��ăݸ���E>g��^�E�7�`�C���(��lz$NR����H,qx-���ߗ��$@*�)�ۍc5��YY𶂩�\!�Q2>��8PjN��!s��:�D\vC>�&�U���!A28mx!8&����vя;�K��:��O䢍��ew���\�$�*�M0 �6�2��ȀRe�_�|��c�(%���Xn#`���ބ��'�$Y�1� �e�I��B�u�6�Ĵp]2E�>R���*���fݴ�l>�oY��_��"D�M�A�쁘9�a�%��V����V<}q6S[2�2mO}�DO�-d[;�g�G���#�� ��Ҫd~`�q3L:��ϯ���ΝL�=��w*��909�䤮}�_���` �^����f�G�%���紏C�?w~��N�)6f��5?��3�k�Z�&+ַU��"$��6�]�����q`�"���G�6��C;��Hڐ�_��
��P����	�C�h��6�	��e��[C�=�`U����L)�J�S����ͬb�<A�Bl�jd��b���n��ʽ���!T2�|��O�T[�pfL���81���E�PMv�*c����=i���z�@lQ%�ױ�JJ��4��0u���T���bu{��Ӷ��;)[U���h���<-��c��C� W;��@��Ġ������9
݌���J���8��h���]�tbO��8��a��4y�g���B_i�d�С��6����'#�iC�cr�n<{���pF�/F�S�5 Jb���# ۵�3����y���l9_ta��0s���h�hi�F�F$w��xj�4�vG�8����Wܮ������0�H����3aS���9�c�R/g�6 ��D繊"y�c�[�����~���:�U`F�C��7��Wp�5���3�����@�~a��LI��g�{�1a��:6�Ԁ�o��;�~#?��q���_���F�[��wsˊu�:�e_��!��*����������T0��/De{���I�A��Ϡ �a
7��ԟ����J2Z�Y���[m{}GE��S�C�䳁0'�b�V�!d��\�aC���ey�L��7Xb�0"�zǁuU�e����$��u�N�%$N\�P�j�w���"qخ
��"�����3_�@��!�"�w!0�r:�7宊�ì5�Z[���L�m�b*
ݿ�:�}-a�A����4�G��S3�83x��H9�cE�%��N�rL���3B7��"	��)�IC��D#u�������kjC�)��⎻#~2��P��8`PA�O��"��S]K��<��4�"��EA�����g[WB���\rbX4L.=L+%zfKiQd�K�P2L�E�6��YQh7.4f��R��a�b��q�������D��!� �>_^X� ]��D<�����~܄x����H�)R�@�>��f��r#����]ROݼwdf�ϳ����K�nAڙ��q'j�����q��\��Fn�N�hM�z{g9�_,�K;�V��e$�R}}T��uFkE�	HV�`E�ٮ�� ���E�i$����z� �����DG�"oc�d�lX�����܂�%ל˪�'Gq>���s��/��^Z�"3p5J���J�#�=�=���x�A��׍gȟ������G�K��5��fA��G78�p�)n(�!��o8�*g㈚<�j�`e�3s=˓�c�'�~Ѩ�#5�әwV[BF|i���v���Mꆮ�RY���C6��Z��IK^0.ր0֕,$�4�D W���ȹ�p���А����.�cZBo�:�ſ�N-��q������Ϯ��M�<D��/8��`��Ƌe*��FP��1��?��(��;�g�;����1��1�ix�e��K-Ϲ������[o���Ш����:k�`��W7Ѝ+�UAT��"�A�yHr�۠��ƒG��w�G�0B<��`���V7�����?<�}S#��F�~2�j_ŗ&*دnCc�����Z��x�dE��m�i	a<���|����\{���~>䠇\UigE"9��`��Ŧu�8�3p�� Т9���֝2yVi�VfG�7��3�W�7�A�|׫YVn�������([��}�]Y5��E�����s�
O�t����[��j)þ�����>6:��B�F& �+"�@[:�hDI��B���7�I������b�p��LG<�P��K2�J���`����ɑ${�����˴��t�^$�o�B�ݏ�#uf�ӎ��y��#�}��:i��_�pf���y��� ��$�B��2Lx"E���o���$V�?*�cn_T�L�DG����W�|�
���/֭ "G�y���oJ��X�RB�f65��HJ�3��fqd���t������ok��R��s%Cp̯�s��1@T ����]�ek�Hm�'�k�:U��V�Y�+Q2�����:
�h>����_�|��
�Ɠ���l.tGq��>l���a��R�rÌ��Z9�>vxv]��)�ɭKG��$+p��V�^|	�9)��aF3>F�wy4�z^�����{Ű(�ۖ�#S��f`�4���^���V#��b��)l��LvG�ȓ7�����<Dj���^{:W��(�m{�wڰ�+�Z��_�·�{�TGD�S�|#z#�8O��7,�,��6]�Q׬	On�ܦ|�)��!|}�����j�˶� X~x!�#��_2?��ц��׿�����倉~������ĉ�0�[2���Mc��/������|�Q���B%Z�MԈH=e�*m{v��A�ә��e
�X�J�G�>Z��M�?4�Ra�R�˳ρ��ʔ��Dl��8�`����2�꨽�WU�P�NY��,e:D8p7�7��c�?��w�v��|��fD���y�Q�_�E�{+��NW<���(Ђ9��k��~@2@п��b�O���t�T|�x"OFf�S�#x�C��c'�Z�d��FBC��:dj��p�e7�go:x\ȝ���)��_ۊ�W�iOt�( 50ރ���%���|D��7�ba^�������%����W��}F��N�-9A0��
;S-êF�;.���a��x���Ծ�)%l'D郂�9��3�Y�Պ��;��(�?8@��j󥛑uIu���	�[4�)�l�Ud\t��?�N]��R���kn'���~���w3l��9q�{@]�0G�hHw�aF���z�i��U��%�z��B��X�VMCl�$Hw!@�������Vh�T�!	]h�`۱��g���A+�AD�@�������G�� �A���K �۽����׿�_i�wM�ݕ����(��ds���Z�Q� �OB*������\9�[�b��D�.��ɚ����� ��)��v�2�dˁJ��Y�ѻh���@��~X��Bw.x���k٨�,��X">���gٱ��7�
�P�w�[x�a�Z��vW���/ڜ��3З�:p�u��x�Sx�ͥ�m�J��M��k�y���+�~��י�'�Z1���6���2ͪ���-�Y3���,D�	���3v$� ���g�V c���׷tX�Ϡv���Te0g�:R]G��R�MG�AE!��54I�l>O�kTcUR�"�'� �������I��m�*���i��6yl�Vѧ�k)�;>�=�wP���d����Vc�p[}GE���nT�HЊ'�i7Zre!wH�wi�Iu2d����~Z��!��&K�`F�l�����\A䵥:�B�����0,�,�5#/�Y,g�8<��%tL&%���,�[Ͻ�v)Ggw�D&Vg�4�9$^��;!ƚr��zB��P|񧜨7t�$�UT�[�t0��؆�V��0}ߴ���5��*�����.��W^g'@�(%����c��[XY�g�r���M\v��.Ù���++�:���)���'��6��u<ǎ��UVU5���cC��zt#�$���h��=��s����<��%����mB�>�v�޿�1���r�LN���<N�{ܘ�I?,�|��r�2%	�[�╮�@Đ�嫜�t!��7�e�_�<+ʬ��B(=��QR��Ȅ��4��(�X��$�۔�8kH�J_p�.X�"H]�Q����O5�<^�U��Ed�G3T�8��,Br��X}gF_|����N�fi�١v;��r�l�. �$�j��*k=
l�+Ư9<���:�*��&1i�!"���+E+ÎX��� �bS,p�v�BS@J����9���������*���j�p��)��6�Z��y~���aՖt-�m��=�b�𭲒�R��s�W ���Hb���������<������Âh�qP�
�R���+�� �[POX!���Z8MX��wf>kZ�,�6z���(����X�m��<�O�r�k'�G�M=C.Tioi�r�%Ѷl��
�E8����/�\e_����݉�d���|TP�:�sI��2��WwuX���W��>Y�T�b}�~r휞��ˤi^�봑a�ik�h%��A���=����~/�[mN*
����W�8 ���a*������׸������c�ps%�̞�+Q-?�[�S6�s�@�"�;��kTt������?a�-p�#Mm�.ڂ�������;�2���L,~�7/_~��×���.����	g'�CΐZBS�a�P��0􁺓�	�6���;��u�v��гRH8���>�+|�D��/`
�����K��6�햪�����P�����
0l�,�ȜD���z��?��Mx�Vy5*��(��X�t̀�o�KJB�R������$p�SD�'�_�ڇK�+�W� �t7�8�mJ����T)����=�9�����G82�G^�Շqc��}>�3�K���ɬ3Ʒ���ԍɨ����J��K>��􁶲��Z50(���! �CP�S^~j�d5Ny���ʟ>~��՝��(Lր�����n���@�#� v�R�ג�̺�i`��%��_)w4!̹�̹Z$P1��>�$(� ��bu�:��p9m~�/��Յ}��Y����Za�k���%]3�j$#j�
SȣP9H��O����Iʩh
K0�|�)�Ή����q8�@b�5�j�]�J^�)w���D��+!+�kj�9yG^��
��'o����S�m&���ms��;���un,d���Í�^t�D�Ņ&I���`��r[=�r���r=��,�ωLmP1�q3D�sQ��ฬp=��:~o��Q:_R��II<��a��c�jzw�a�(ƌ�8̕��Į
�»�I��*~L���\|r�[�!�a�HՃ;���Q*X�7�(�zl���]�&�	F��ƿ�
�r�&��\U�����Ȁ�K�� �"Dg�bY4���Y�\T*��7��t�h�~�#R�'ۮg��#��6�{v�tz#��cb�� z�B�	��iRy|�ˬ��/�C����f���N�4��xRn��,T3a�B,���]B�{i�����$�r�XPCG�x���7臥��52Yr��F*��b�����N��_���V�Z��g�Q��i����6U�wu�
Gy����$"ʆ0�y�u�/���;���x�i�u��a�yv_0z�N?u�D4W��'�Ԃ�aM�_�Ҽ���F57h!��WG^\��&qV	;��&�-0[	Q�yT⧤�f�H�m+�ql��6�
)��X��%�+�`<��eVq2����-�2��Nl̩�f� �^�)�����C*v�ׂY�w���@�CQ����Fj�I�cu�̱&�?��T��	 'D�\���������(�$�Q��Q���x����dO3X�ƮP6<�%���<]�-�C�.���EG:�.!})Vj�N�$�̕jg�Jl��j���=�u��q�ճ������o�Bk��>��フ:	w�
�_n��`��u��I �� �Jh>�Ӯ���}�����+,;i%Ewe�5G����}��6F�� ��H
�RW��uσO�nB(�&�$b�����y�����J�	�K����]�����)=r���[B��J���5��XE"�H�T ��uv�J6͒�?��n'Nn�G�c��JY�o���U]f8��g�PWټ3r?�.�����Y�V��n�:R%_���P;a���OX��r��L@ǲ�`^�j�+OP�Ў\�k�mU-�6�	�)�0g��0U��wg�|#��B=�s������ �E-���*6#!�����F*	l����cAu4���ɵ'�&�a�_�9X��w�~ �����-���|�˂ �؆�k��W�Ϩ�ς�,��d�R.����Xu��Z6�$�[��%�Q҃@�� ���}B	�V�BMI��(���c�8��U>Ш�
�R��U!Rp��g���å�U�����җU�9�5�J�9د����J�=�K���o)��\������價I�;%R��FSkQy})�`�K&����U�wˌ�p�Lt�qؼ㥓��Z&���+Ю�
'Z�+����5��E��ImD��Hd^K)ʘ�W��V�T�}ڴw��1r��� 6��1̃�XM�;�d�A�U{z��P���%RP��e�����@���B�c�uFs�id��)p\�Fuq�m�ꍀ����p<�\���R_7ҭ'�lEI��^gT\�0��y��%���`�T�9��B��� <+�Y~=�ay�o&D
�I�C7M��?����$X��,8 �`����c�c�.�{�G�R{o���~*� ��a�E�3_Y���1������@Iwg��+O�Ǘ���|����I	��~� B�B����X�!�ޏ{�"�Ƒ!I�A�Y��ͭf�*��PX(Z6�(�zX��+���#���[�)1�|�KPf���@����x��ĕO{%/�m�^�r�����x��~gK{٢��|��V`R����M�� ���`6U?�./�Dh�F����S�$�e��k�0\$���?�"R��{��V:�}Zd{^A����9 ��!�#O۞Y��q9�������&1�0+�!l~�l��FG��\��0���O"e�Q	4�S�)�c����n��?#�#Br&sr8SN��h�Ŝ�˦�	L��������-���*P�)z��s7ɬ}�O�޷�O	�2n���Mw��~̈��A�^'ޅ�]Z:3΄��,��较���FLUl��5J[���EC�cÄ��Vm�����PJÐZ[�Q��)d��*!��d[�+��R�
؄Z�rwϗH�ݍv��Y�tk��Z�ױ�~p��r�5@���]=853C��}t���E}�����t8�����q͈�K�f�Qy�]���f�$Ɂ ^in���Iż*)��IZ;��l���"N� �q&i�0-}P50"�.���N0�K6�e)A��2  ���Xy�T���O�w&�GhyQO��ÞΌ�k���#�L��
���^Q��̄
���ghF4��B�OW�Y/��RJ���f��E��p��Ί}���R<����>�g���@�J�(����ͪz�9�rD��MV��R�
�v6A��T<T�і���P�I-*5�����׌�@�/\����ɹ:���)�8���>��/N�C�~����M���/n��D��S.����<�1I�'Z��Eƽ���2���,��.�>;���8�l��&�2�Ȏx,�z��3��FXHzKG�̢�꤄�2�۬%��?�����?��ׁI����y�j�1�G��`����5�f�.��\��M������|�C�;l��'��8��ɔҺD#�Q�v#9!U�q�x�|�K�ȇ�˱p�����s"A��*]"��(Ud��%��-�z�t�;�$��"n��È��İ�$"�G}
�z,�RP-�W�Z#G����Y�?��;;��o�#aw1�Ak�/񟃞6L_�Yo�J://��z�KbiqR�|�9T2>v=D���tF�وS�����wQ�+��TӘg�#�±!*ئT�.�
g�V�o>�GB�DQ:WHT�Üw����WS��g�u����I��KD0�D����0�+�#έ`����f���0f�-�?{�Ct��C<�i����h@jQ_DU��sT�����q'�c��|�r�k���Q�	]��~�H��!�xEay�T�+x���R�ǻo�$�qm��� �k\��_O@��uU%��"�b�JE_Ҟ�B�̋5�(���`fŨ�p}[o�,�n�6��s=��e��աЩ-cLH�R�U�AQ���"<�!�\@��9>����[���N��ƕB̎�rt�#+\��V����X�US/L���P6��-*>}�`X��*R�w�ݭ+��L����Ι|�� 5� �bIYc��d�>mB�fJnQf�	08��4�CJh��O�y�r������톮����B��Խ9�x�ɀS���,�~�[殹�F��iy�=*��a��l���mp
H'D�ٞ�I�rk%k�~�����F�����m]�����;j�N#j(H<M��>}5	�n�]���UY�C�|�(�]�$�V#�Ξ�5+�ߧ��RL�\X�g]]c"�Qc�4Q������QPvj��q\��E�Bh��˲ק���R9�FXeN֝9/G��v=�
c�.S?ד��*���8ՙ���稲���7�8�[ �^�'	S�~9��]���GZݥ9��W�o����y�o��0�0�iq|�c
��D!<	i�p�ǓM��\���t��}�#�)V�m�!ۮ/�b�m�_�J�Y<��Y1��	20q��C��.[NyREHl���a�z�qd ��`��<���{�	n\e;BRҊ�眮�zÓ��j��	ֺ�l7���� s���_��E��ę8]'�Ǆ���4#}�ib�x^��.������0�h������m��W�LP8�X\%�|G���"����Hm_i���0��7��LS����9�p�Z��;��U�����&`N�B陂|v�e�7>+��8fs0��B�6��7�b��l�|��(8�n}��
�?5�K$��3�z�<ʇZ��eW,�k�bό��R1����)3;V�g.}f�-G�{z������q�Tb@9���L�3�}����������ଣp���/��sV�p�<{g:������6��>�����n'�l�z�)� ?�w��OrXڟy�o��w
�Y�i�Bv>�?C�S��uB�/��6/�.*�A�Uj	1�Ti3��·3q5��YI3L)�J���2�z(#��1M�,5D%��緗�fٽj�sr�ԯ���@/���:����|�-Qp�r����R.�G�Ly�}�ޣ����{���A0a�$�>�Y¹�7���W�ܕ�Z��?���N&�]��5B�4e�y��G��Vw�����s�R��P��	'��-*�I箸����|8��݀%?��.�5#�m.V��^ʯ�:��N����KV��?-/��z����g�	�y��ߩeT>�hU)��=���E˶�+,��Ő{����6��WQ����[�g�v�{�.9�`S� �+�����>$�'�����5"���;�W3Ӑڱg��)F=�h�HO���_��=�����ҽ����R؊[�t'���jr]���2<$j_��mdL���y6��Ŝ笜�K#��F��J�I�V��v��ͳ��%N@�յO"dT����D�j_|�0՗�.beޛ�(�<yG����2�����>��dG����qp#;<?�Jg�{�Xua�÷�79�{r��dXN�B2�Z ����1d	y��������v!���uo�<��+����{'� M��)����tTn_	~/�!�����	��iY�~�^ G2���J��dUٹ~�*4Y�:W�"%+�i>�F&|���a���a~W����m���EE���-S�1�䠶�V��u��z{�C&���O'�e��T�V~�@e�	�P3���H� ��� �?�����-��As�j+E=2��ܚ�K�H繌�LO~f�&`�Y�rKKV݄�I!��,<<�UJT�Gyo�ܒ��~M�NlS!>|�0��P|p���;�'aȏ���WE�����a���ծ�S�E)�5ƭͬ�����ל���@��o*�߯��T�ʵe��c�T�s{k]���f�B{�c�a���p8gL��C@��r�,���Nw���q�����p+��/�A�F���P՟�E����^�6�V2_I`��E�ɷٷ���ͰE@k�I(P�1�g�3�-$0|�� ߆���=��m�g�䲁GCp�p����6J	U#@���mQ�ѕ5e�i%Z�f��@��OL� ����bq��t@�Fk�MR���y4x�Vy�@�꘍)�8V��C����y3\���{���g7w*��j�d�<�w�_e��ѝG���ܙeQ����?-��z��)AO{�K�>&hK��p������F�-��W3��ي7Q䲒J>7V~��g��'c_d��&A��+0L��c�oF�W�wORY�/Hbp�zn��G�������*wLn��*�����dn0��4h-���Mµ�9��hIƱ�)�Fi����!.���d���7�]Q�k�����B��k<U�ԃ�^I��� �QU,|c�pv٫o���(,�p7���r�����x���2\I���g+�i��]M���HR������%z:b%�v} 5*K��7	w���8E�>�3ˬ��9�M�j�_�=k��c���s��K�e���%$�W��3iYqrf�]�	j_i�ULGW�Mv���Ni9�"�Y�\A���`��? �F2���o99+!��LD�G��S��T6
?j�zN� �z!��÷���4�2���S8�$N�:�;$�V���K�,8<#��}>:�ծ��p��5gP*�,�3M�m-�-�æ��D7<
� <��՜M��`	j2�Q���(�v���"!<������KX��f����2Ԛ?/p��4E6��kD��.\�A��g����0�X�7�~˩�)�a���_�0���/|�r��}|���Z���&��2�~n��]�z|�p�)�¶�M ��m�� |qi���,l#�Ë*;�����%�_,���`V���F�<Tx�x��يhA��N����Ê:��-8���紟��٩�����_�P\�&?g2F���p��? ����G� z�r�tT��mҺZP�U����R�>�vT@oPn*Z���OW�]h�zMJ�s�-y�}�����lVm�7�	� ,-e($�9�/:���@ QԬ�4}Wm���<�:7��W��h1�����p��PP\���U��	e�Z7�ז>���>f[*,��N~�@�GCut�}!����U`J�ZSUtӌ�h�Z6�����Z��%�j UN��z����EZ�k� ;�|��ݞ֤E�:���@�h����Y @>S�i�\�g}M���o��"�?�c_Փ�������w�ۤ���zKH[���e#���͈���1�A+��˽f��. ��'
�V�zKx�@dX�H�i��7��)��a^͟�
�"n��)�c��?���o�� ��Ϝc�U�� �.��-dS�2`������ڣ�i�u�p�f6)��B2�1�U ��D�ǍG4#�k��-�Y��ը��]�ց؝�>�͑YF�HD�oCׂ�%:�?}Tґ�L��+����[�C-N��}姘#�
۔"��6�&\庻�u���L��A�����e!��"��w3�e�y�Ax�Z�^�F�Ƚ<�㻓ƻ��8����.����p�4���@a�}�GӋ-���	Ƹ|�`��x�qwG�D}0=�Jk��x��(�-t��O(?t&��,���N��WB7�
bs�^IlnUcT��������X[���_WT���x���f�d�8�A�D�\��z�7�rȩq��{2��h��3ZMgU.>��:L���r,��}��G�a����;��|6�с��c����띔�y�F�pS��{Q3i�x�|F@�Z.�.�.�X\���`���o�MU�o+�.���b5Έ��Wy|���
�$Z�Z�K�?���;'O�zf%B�q�ΓQz�	�}�c���TRˎHYF�����m���P��쒔�g������v镾��
ה���Ƿ��D������
�W<�Ő��OޘN�_�^���@^��^�҂;�U*�_��X
ٵ+�v���7R[� `�&�܂ܝ�x���+�O�=DL�A�ܹ��*�����_���v^����yO�?4d�S%�۷��ץ���8o+�d�Є���H�T�:LOH�Z
�����mCj��I�S{$A�hP��@l(��Xk �yB-�����^78�R>b:��'2m�q1^�Um�im��o���F�v���/��<��[��t��=�J�7l��L\������{HJhz�_L�f ��9�s�T���2z+�_Ø��e��t���ȫ�:�|��N��*�C&?$40Z�JE��b*(�1�&
�u����ƅL�	��0�H�%؈�sr�*]]���#���;������l��%E�p|Et��Ę�X�|逽6Cv��`O���I��/O8E`q-�3���<�q�U�j��.4L�"I=�nθ5�Ο،(U9�3�q �5��D�_ ��IȦY�5��0�&�Y��:])���q�8��S�J���%[�j}@��~¸x�- Rh��	1�T!���t���!o��g�'HL�6��d�8bh1�%�����H�(�zpS��W��F���f��ok_��Oe�6Ʒ�
���_[�}�#�}�J�/����t7���C�6�R�<�f���� ���+8��J�3=���H�	՛^�I�i���K=�`hZv�6�ο�yVN1G_��HX��gz+�b��$� �Yq�IH.�E�^޸�I�n��Y%Nخ}�\a�"􈏠עk.pS��#AtvA���Z�����/�S��[*^"��̨��Ҁ��R3�����Y�'���hF�h&�������2��.�Њ��ns��0�A>Y"2�0zߞ��`�B�y0�Z�"����A���l#�������u�M,l��yp&T!w��H� F
3����dУ^,'!%J[^@L)6?'�u�r�B~}^�O�����he�:��_=��e�����gF[\���^%�z�	�Pr��"�ƣ{�y����w�����a�M��;�����m��o��Ǩ"+dz{�YjQ�;���}���Ŀ�H_i�{AY�ٻ�ceX
t]��[C���,�N:�V/�GM`nPQ���e����ڄ��V{���g����j_̇�k-���̶�>��cU%��"�|��EBk�v�gM��,��i@͆V.��t��B�� �ha����u(Ҕ:^��Ȫa&���6�
c#QC��zt�=��t6��-2S��O�+�gU�,��)��(��zm�J�n��c`��%CyO�p=PSE^\��X��2Cx}�#�o�g�(ƃ|�l-�F7篧&G�:ԓ-p}�� �����nc��o�z^Fr4��\��f4�?AT��l�ʘ�����)j7O���/O��RH�J��5�}h*?�5h����N"=��{-�L�����|ܑ>4�xi�$38�����J�F��oalԳj��{��/��G"�Cp���N��(ݫ'R;*�`��.bnf��֚�b3Q��]��j�龈A�)I=�����D�񱷿�MΰI�hW���o�
3�,Ո����A�+)􅰨�@���F�ċP��z$bH�{)�.� �����Ht�`�I������������)��q���B��E�3멩���x4M�K�lYA�����6<mQa`�lԷ@7*Qaq!�o~(����<m��"H"�l�K���,8�Ӥ���Yd3��G��QKJ�h21JO<�ƎQ�an(8ힺ�%��@x?�dn=�l�O�}ȚP�d��YO3�~�Y����xH�=3�D��Z�������!-U���4�FH1��.�i��}�fE��Z ǈ�Ez>�r�������qZ1�a�e����FV�%�0 �b@XA�!��d�	�F�j����M�������'�*����D4�t\W��~H��`��R�ʒ�q&݈!�j���=V�[艆0�ע���ޙ1v� �X�z\����B��M���߆?�m�8�wW�2���X������oqs�;��*E^"��$^]�v�o���u��]�B	K;`��g����#�~%-%f�F�CZ/TL��1�;�@���2���7y���/+�i�b��hhᇢ�s����Zl ��%��ظ�l�'cf�䧺Vu(��WT�������ͽ�@��13��ěSl�'��k$���QH�6Ʋ>\W~Z4�)�m� eH����w�b����GB}�a&�x��8��~5�Մ��#%���<U�����w�a����[���%HW�RQ����x�\w�I%=_˄��_dn�D�l7���:VJB�/`5_\�ˡU-�W�u�4+��v�^6ĈFt�
�J���ک�����Po>�@��\fd�=�����(<�]�6���+���M2�Ҵ)/r�R�c�9*�R�r�{����	|\ʿ��P1ނr۱:ڧ쁤]즙a�^vcS�͖��RM�^�I��N�z�3n��l _˕o��	����纬֌;��%���/F0�"�ėQ�5�o7~��&>���];� ��iGl��n��Zq_��٧��JLx6F�~I�.k�U�ӡ{�aCu }������X4�*	��ߤ�lM.�� ��X�EXP@�-��=>)�j|��]xU �I��LҾx?�*Y�U��/]za���]�� }ˊ+�V�ݷwp��%�Cב�O؄-�H���|�t��o;&�@����}@���8�"jwao�U�5Ծ#��Qh�O/P��A�K>��	�ho���;�T0�E��v92`�0�.4�I�Ba�$e�Q[�:RtG���/�SN��$I�)0���]�D�x�1·���(�=�wm�kot���X_�Z/�0?�����np��&�@�x`�ЯCkp&#�Bx��[k�/�1
&<Z������Ɦ�qm��"�ĥ�lm��]e�А�]�!\�Ln�Ճ�RE�xZ�_�huI�)�N��F٧�aL��
�ɛ����$h�U��)��·gZ�y��������Z`_~�[J�?~-�/�Z��,H����Ԇ�����U��gDZD}"�458G��9.>�%J���H���r�mL�3t�UG?)� ����A,�9[b��C��Y(Ξ4�T��[P5u�w@"Rh�Z���ND�Ρ+{����.
�1�K#��	&[�]:�:1vcy}P��@���e@E�k��W���CхF�)/���v�U|�����-��5��sj��z��y)��r���w�?��w�������^.�I_A��("fe�Ck%ɤ�����ݐ.;�B��c�6�  ���_T� �	���� &�h��^ٮ�)�q���R$���'��ī�x{�G|n��)UNc;z�#w��������Ys��1V���Ffט)u�3���*�5�5k��Q� �9������2�dJC�G���32WۋJ�|����?�'�ޝ��i��t�Z!n 9Uy���w�乖ю���ɑtG��}�6.$4��#���m;=�،57��~�i�S��xe���O��Dz��*,��Tgn"{u�B0BY w����(�#�F�f����ݕ��]n���AFX
?C��k�:��7�D��ǂ6�v���RK�o�
��/�����_��2���Q"�� ���3v�$�`F~�<���ژ�W�u��Lv��t*1L���'�?��2fg�ˁ�v����x]��N��q�(�Z��~TN[��,�n4~A�Lc/��i��u�K ��9��|>�b/׫�1��ܸ�͖rq\E	"�,�0�v!��?�P�3�X}Q�휻����%��<��86��7�k��p{�% :�$� ��.�hH����u�21!��AX0��7���N$��y���,ȳNb��]'�u���Q���� \�n��Q����ăBs(��?ۖ^}�"RUŁ9}�w}{�KRB$1 ��per����:Ȅ�����8o�{Pf��8���,�]��A0mu�<!������\�������5kR��Y�� ��O�j,��,��+n��d�,1 d��gn�~�;ǹ$E�����Z|d�}K�u��t��,�M��5$<�˘���"&����vޒ�6�aS�q5����ďΜ�:�n2d�6}EC�{� ��놁�Ox��'�(�PO�q�:&m�֠��"o�y���d3 '�!	��v�OT�Ԕ��`��B�qܨ5�?uש`���%�����Ф K;���1��ݰiQ�3^���J��*	��ٳ"������M��bZ�/q���w}T?��ݠ�g\��@$-��e�۞q��S�W�%�X'۸gH��M�"7�.���y�0X��ּ��+��y{!�+n�i�����[Cn!h>�Us�rP}���8i����4 ����"�����a���b6ЁFb���c-Y˹�IM��`[K��,�=����>a��Y.t�;@�j�U29�\�9�\��$��iC�t1��&MB��w[�i|0��pM���eG\Ih��k
����W����������~�R�	X�2}yO�ɋ9�CO��r�]�ӝ�;j���K���thJ��;"���BeZ�So�l�֒j�:+��ˇE��<fOρ1�N	��\y0��_(w
׻���C���`�՟û_nT�[���l�jb���n~
`�T|�oN7���>-�m�6EiD_j.���M�ب��Q��?��P�����&o���3�
�b�7�5�o,ڍ�h!����O��"J��~,)m �T��c�r�S%�� %5��,��E�ì� ��;u���o���hz��R!�����}�~��>[d�T�R��~),�+��^C0s/�*��ɖ2B��ʥ��<�=Q>ɡ�ݑO�������{M[�*%��8v0U�/��z�K`#�1��{��뷥pR���X��U��l&�����6/X�����F�൶j��B�&P9u��Q��m?�PV��Z4a'���W�҇+���/`�I��(5��Ҏo�1Io"�e�'���)G���[+8NmqsMʈ[��'�T�����C;��v��d��}��S9�:�V2�'�P�	�l� f������(���ج�'�&E�#��� 	��c����k�=4{�	01�h�x#�߽�s�_��a�p>�CO��k"Q����*ә�M����5����B�P�y�E�x1��8Ğc�·#�]�0@�C������M݀�QL��{����84Ap�"���i�s?�D]i�y��c�r'��30���#�����n��r��"��A�(p�7!V�O���6�T[��o({	y�M�֦��"�L5�7�+��Dc�P�F� ̥�c(J�1|�X?��$5�id� 0��^G�Cp��6��@0;�QKf��z�� �Y�l�h���m���&�7���iA�efQ�`Rh�G��<^o���� ֳ�/���P9)�H�~.ʛ�^�
� �]�;<q�3�o�Sw��̛	+��Y�1˨��C��*ސ{���.��'IY�_�"��O���x�'C=P��*A�J�q�'�%f�"�̀�*ƺ��S��y*`2�ݫī��,I�cX����u)~&L��f]�u�m�TDz��"�v	o�����+��Yd��q�r�2<�2榐���\��������e�ՙ��.+����l?�F�W}��(��*�\i������@�$�?$&�'"���߁O�!����7-N#c�C쵱d�������gb��<)w�^<��1���L��H�d��D�-CB�w�\���VD�����]��e��A�gx�H�[���F����:�$᡽�X����9�ŧ��R��5�Cq�~�xOR���^͓����	�G�����Pu�-7�^b��  �%՘��m!H�A�-8���ą�]�@L�|���\gV(DH�>~�.��֯Ơ[@a*�P{��j�;t��M����q׻MR�6�|n�?��.��� �J��_�#��t&���o+	f�) ��z�2.9���p!#�oc��o�d�����[,�����2��C=��|��м�.NID����7y��t��b�i�,Z�c��s�d{z�{�N�=A������:-���LG�q���=��@9Y]5?zڙ�RhVq\��5\{Ih�2���i���$���'e~P�w�r�gp�ǰ!�8��F�u������=H�j�M�� 
�_ew͝� G����1�<����ӵsu'�'�8d{�2�̲D�M������]��=�t4�4~C[`���E�ȣ �pkh�`�0�q��s��׹W� XD6MB	m*��zBC��]m�B�}M�}��Kk<�Y[">s[�:�bEv҉�7�|IJ�BSq}Z�M����&�!Ʀ�S��H�9�
�pMal,�V����0j1X~lޘ��(H����<7g�6�&ro�d�`��e��N��萂���n�HQ����~�8Y��4�{�)D�k)�������m�H�|�Y���������mc��6�|F��v���#:jg�Jr{YN����Ř}��K~�!�oA���`��.2-��u�p�cEA����EZA}�_d@���3:��sc$n(�o�%-64ۘ����+z��r��m��;�W���3ǂN�2�~{�����bh�b�����6�C	���t�#���C�$��T�U��\o����A�2߹/
o�x���/��=u0�ghB>�^�bE�� e4�C$�e-�{�䪣�,"GG��2����Ty"��eR���6��mu}�:曙)� kBq��(���j�r�V�a��+[�������F4V���R���K�l�8��QoW�gy�����8���g��`�2\h�3�`}��i�:����P}6z��{�\A�Ȍ�DF�?~�[��U�"^'u�0�\5'\��V���x
�~����,���C�8�ݺear��A����-\˴�[��3g/�ҌA'���Wǔ�_1bhpU�,�& ���U!7�^��n�{O�Js ���J#�l��$7�m6fXju�TY�';sh:��E��0Dĺ� ·I�"*��5����>�җV|���ɠ~��"b>]ż$6A~��\��e��nX'.�I��`wQ�Kb ڧ� �؃[J��2�{.ѻ�[��M L��� ��I��
%��宝�V�i��H���ê��K��	�	�$y[�#l�˃���Kd�� ����gڼ�L<�z�9����1u�)�����
֚#J�)?z����@vR�S4.6j��>��0,ѯS	iI�: �TD]��s�Ā3�z��C���O4�dцq[�~x2��w����{�;5���4z&��-_�PX* dX�� �S/���0ޯ����m}F�ڞ��䱗��,��wnE;d<�0E+
���A1��������O�Ϲ�I	�ҷ��o�Ct�9_�yDpSgH��W	�"�\3\U�l�ތ'�`p �izwY������1�H�{����mI�����re��+�]��K�M���sC�D8I%:U�P)�b#ݮ���Թ��@��9'U��ڋ�� ��4K��CM�P�u%��ˊ@�ί	��y�� �$S��4C���$������q����-Jѳ9@퓖;m�L��i����:�*�Y��aqlU����3��K�xq>��'�f�-s�ݚƂ�N�1����l<R�Qm�B{�!�S&ؒ{G2E�.��p[1�����>+�͋`#�FeN�>���1D�4R�=��:�'O�t��m

2h_� {0�|�rJ�:d��f�G�F��*��\�Pen2ȏA ��4�] 884>y`..�t,���b������	#��Hw�f%e$��n&!4��Q��lΈg�?�7���$�]�$7wX?$��Ü��O�܂tt��i�ƹha+�H�$Z��>B[`@�+CU�K[�T��Bbʻ�����U�=݄j'v�>�L:���/�B-f�_��2p γ|n蔥!_]�:���S�x7����vbeD�@�=�j�*�H�X@Q��P�k����?�ҦL6C���ݾ�*���ƶԔ�Wq֚�@m�ߢ���l��G�/�jm�ф�!�ɮ���Eܑno#-bL���s��uF�v��*M�&Q=usN�M�L&ph���S����o!�i���f<�R���2[���H��&G�I���n	ٟ [ ���ٍ�����U�Z����n��T�׭�GZ����Pjx���%z���j$Ӂ*�n��K�?�����'�["[�A�EW��I
����w��t���`K��� ��"oB��E�>�b�.�GJ�ke��C��Yڸ����!]�f�~��9����tw6�f���NQ��ie��f�܍�$���yxp|�5�`��K��xQq���m��f�$��jE+/4Ց֎���V$D�MN�vz���X��4��j'���*{]�R�D��z�=��2��z��׭{9�S~��2Kl�%�J@Ҟ���W�D����7)fX���퟼���W?̚��ʞYJ�:��Vi�5G�H[�h~�o0}���,�]]�F��@rJ�Is��R�M K3�����&�5M;� ��OA���~�;��x���jW�a\av��m%h����
�՜����N�(^L�0�&$�����&�)$t��|"Dq�c:��Wuf"���)U&�w�q���ᖔ�>�LU��y��:���,ÃG�Z)Goe��T֊����@B!\���lKr�J�z4ڟ�K8C=�Kn��!a�3 Ǐ��lRD��'�<`V�ħ�6�X�j�Zgt�}�md�y�3莜�ggfU�Z�J����;� ��b�.�F�?��TO�1�2B��쌻F~�hsR���&+}M!4w��o�ц���8E�h��'�mx��Q�|/�+�J��x p��'��z�ACU��2�g�Ӝ�?ęL>�&1�+��z��mu�����M�Kp��F;��ФQ�3,� =Q]C�TFk���5��� �gU�7�ʾ��Ä�l���I��G���s��8����FT��� ��?�ۯc�4[�7|��Ɯ[��K��)w�;e-(=���J:Tmq��>���o԰Av��Ϳ�����^R^����6���ң��g��]�֋U��v�?�^�-c�Xj	VJ\����T��p���@*�I�I��rdD�
��WW�x�Z�<,���r��V���,��9��)+Ng���Zɷ�?!V�_�i
��=�2ݬM����RC�X��i���ݜB��*��φ_.��L �&p��}8�ꍦ��_�J�8Ň_����(m�C��ǡ�]i��$�h�G�`�1��.�qp�.�L[��F�b�U�H��lY���������*٣���y<#�~�,����x����3�<O(�=�8����&*쳌���>�%��Vx��Ŏװ�p��+B;H2��:�ٹe+m��ٟ�d�9٫�� ��/9_xV��|�_�h�{�kRyB�V:I#��#��<t��X¯8,$�4�L(���&�"`$n�C
���M�ma.��$�������8�����������4{���R]Yp��!�榺F���QNKa�4�A���SP��J���v�"���ϸµ�UA<�aF:'��|�}N_�Iwđ��\�U��8Ҕi�K�F�T߆�W#�0�Z��#�Z��Йp�S5��<9>�3����E�R�{��'s(��ƉQT����p��v�����3�j�*Ҹ�މRc�	u�XCƏn#�l������s/�֬+q����:�ç��<�jn~�4�-/����G�%�=ù������K��k�����̩����="��)Хd<��M��Nz� �g��|��-����B�Wc�/��6n��n8��1�X0���1z%���V%��`�MYk�q"f��V��l�.%��X����󽎒L����:VmYm��r������Ӻ��&�<�ťȑɛ������P{������fg֪�Fc����2
4�Ao`Xc��Br��>K�7������١U>��9Hh�XH*�?5�|���V�,?}o0
�������gT����&�u~�x�ݝ�n�wQ�H���a�@��h6���O��N��|i/�����
�'D���Y[3	�G!7B5�fd�*;���Z�E�zd��b�C��MbJ�����7o�B9z3�I�)�ʩZ�A+�5�v����'_����.g�~ ���DkƱ�?��c5b\�������֓$�A8w0j����y̅����~��V�	�1U�m>\|���
@7��ZU��?35��|���m?:)�~��z�N����ψ�ҾB�)��� K�=*�+�%��_!�!oZm�#��bT�L��D�C_ ���ls��M�eD|�aK[ʲ+��ķFk��A6�'s>�u������dE��$V��:tA�%+�9BNp���b!��Q�F��,b�dd����I�%�z`�+�`�F{\N���}��;� ��.(F�	E����^����^�>
hi�i��X:���ZG�%��ں��#0�����E�W�a���������c�}��bj(�g)٣<��(۸���&D,y�C������Be��`��f.��X*���?�E@��3��Ce�~H]��!%`�O�cW��S|+B˧���T�^;��E�5.��I^�%/2=��]|'��Iܑ���PqA����+���*�Pb��x��`�N��@�C���ve�m��P��%�,@
���EH2�%�E�w}�r����h4R(w���_�Q59��|�%֦��Ճ}9)afܣ�fX�}�`&enu<2yb��DZqv��?Bw�{e��n�הƣ����X���I:棇�dz�)�������_�4�䜮ߢ�\�X49�v;����״�+E� �\~z�:�H�]ĸ�Ϩ�T�@���1�=>��S�� Y�$��k��N ��HgiKV������$����9s9���5�Y�ݎ]z�$"}$^����O�h��h�.	�l���1����h����8���?��fh�_�{"c.�K���:��n�``�Ґw��F�S�y�1��r��_���m��8A��SiXҘ\x�cǀ��"�F[��(F��dV�R�:�ۓcvd�Qu�j�9Y�����O�ȿ��3��#HMI<�M�[�D�rX�fD�����t�j�7���hy�`9��u�~hܠ�ٻ�.��&�zoy#ɉ�SA)4N.w��=ؾ���怜�M78G� ܲ,A̘A<�A�uvxP��gs�%��F�$�j=_�yf��ߡv�k�{}h�1�$��5+[L�*c�׫H.�x��
�z��S���w���үUYPm�y����d�^��������^�4@t����|���*t� [�Yv�22v��\��J]R�?�W�|��D'�jx�3߫	V^>�L��=6a<$��	�}A'4Q��� ~WΗhVR�_�˼٣��]gh8�CH	���N=�k5�a..·�,��M��\�n�$�I����l~gV�{8�� t|Iñ/>=�;p׶j`��]���d�6<��?E�nü��]z��}X�2���r�\�T� ��ə��@Y�5eww���k|��kR�wC����Ս"b:l6CM:�X*���*oQI�.�V'�F4����P��`�<�J�XeDh���0G
����i����Z+w��,Wq�f��_`�ep��eC�r �.G~���z�7�Bv��M� �n{x��_�4�Z���fG:�O�]���4�]�Q8�4���>�+6�_��KS��
_g�3!�H"hX&��E9�)3&��xT��8#������O(#_,�h"k�M�l3ѵ�4�
���YQ�8}��\�q��e���h�=�ɸo^-]HM��.1
�ֲ�>��{ V�:�J��ڵ�	�'zii���Zy��E�s��s�G�dT��^����H�4g����;+����_����;~���g��9�@���=�%�4�����	�Qɧ��n�Ro$̏��6Ҋjq�==�m�˃�[����~�i8y/P �OE-�t��ll�����L7NOoВʧC�\v� 521y���x'���rvڣD���~l��᷒Zs/3{�_
�0˿��,F.�#�k�c��[!gK�]A*%�y^ ^IyI�%Т"L�W�ly�	�r�6�-�$t��d��P<	��*x46��F��P�G����@�u4���}�[
ï4pU��<Kd�[��9����	�Qѷ�����!����P��U���u\)/��]�`��\�P$h�O0w`X���f�˶1��T�*�&�V�϶Ef������N>��f̕��c��x�߼�㑵���p�m�x2�@����A�h	���T�:�'F��YS�R.U��򄀒"�T{ǔ�<H�J��^<�����#����~>�HG�آ?��J]��m�:	��dJuȢBZwt,`娴������_U"��\�'�7/���O�g͈V. l�N����I��i_�wޗ��W��)�,�4[�q�+Q��V$�X[Qa��΂\���p������?2Ҕq�����M�x�¢ok��⿘�~<�����*ʝ�45�ti�O�<��P�}{i����Y�z��j2:��2l����#�kޛ���tF�sutq8�'��A�A7)�Li�CG��JLh�}ݒ�����h���Y��1&���z��gb$%�����*��8xi�����R�liw%ֽ'��[�;Up��e-����~L��8�8h���7(>�gϕ����I��*��?r��)*kF�OuLTc%m�xR-T۾�.��"������=�ױ��J�	�B�lܑ�/[IMPU�����f�3J1.�� X�$�S�������_���=)��8���ς��CH	���/��5̀L0�~��A���;�����&rx�p�k��$�N���b{\D�����#l֤2[�s)�|>�f�5ۅiq�`���z�Y�p�([�M4�_�*o5X����?����3pj>��4򻘪�'m*lR��o�`��ic�bxM��w����s�뱜�"q�}��J)5o��S��)�
��Ⱥ�����/�u� ΗM��끛��~�u�z)6W�O?G�W=����*y!�}�~�#��*5�둀^OgE��kt����Qy�����$e_�zJm���C���V?��
��0��6{�:TF�U����89V@�%P��N�ڬ/ƴ�r048�*���Δ+V���]Nd�Z�U-����{��$p���>��C4�1{L�����õ��c��66�|6�=#5�l��޿����.�(9V�������(�c}�ƬH�^�:�簠ڹE㷖Y�L9#H���{��(ݎ�rr2#����z��9o��c� ���'�s�vw:n
�o\��C�𜭑~Z_I����B� @)�hI~i�ANj�:�]�%^�w ��_�pf9�ً��G6��~��aT��i�0?̎��Z}�$'R��ǀD�`��s쳆����w��w�㎽ʉ��bߍ,����^Z������[�e��+��O��j����p�n�R�A�?�~`�:�hR8n��=p��lm�YP��@�]��'��;����E��7eѾ>�vέ�H<@�=MnnG���y�sX������69�VȚ�hE���7i��y;z"�h0�?��]�r�����i�)��
���38�H�<�߫��M��u��t��Q��+��TL���U��{���:nw��+�w1���Tt�Q�J�`��\�	a�+�"&%�	b���G�[� �Q�+�㿯�C���������dc�r:F7,FT@��f�f��
�sghek�ra���9:��^�oe�qz�Tm���L���ʙ����E��C_��/V��@i]W}z��0�r��R�``ץ������q��AZ�c<�x� E@!8��߅rf�]���m㊊o�a'旻<=C1Ϸ���0���6�Yi`�>��YC���2��2�w�K�{u��Ć��B��D�l�J����ͱ��OE�{����wI�^�ĵ��(ݜ��n%��b�N�Րu��Bu�����+��b�G��U��U��i���&�e"��x��ez��L���OF�Z���`8
R�߾ِ����Y�,WP�s"���	/�1�rX�M�"�zO �˛�&=D[n��X��vV�6�kq�T�^g4Z�0���ԙ�c^CR��F|��3.}����:���#DO��8�������YmN��@� K�7�>k��� U�V�Gg+��������8��8"������E:� �"�z���ObPg@���:�$����
���ͣ��B���>ʸ��<�oV�
��U�n.��(v)s���@p33B��--�>c��G�*�Z���̩���b�-�P��>��К��}�v�;ҿ�8꺀����O�)��K�8
4�5K�T)�:�jz�s:�g�>���RYܙgT�6v&UM�k�������L��`#S�/�7���"ҕ�)B�⫭��Y-��[+�^�¬ ��O �kz�1���F>3�q	h6��0�j��3�4���IKe	Uͯ��?���l�.�:��|c�i�ڽV��gS�'|�iu^��bWV���##���ݖ�_7������蝏��a^�s���,�0e�*~v� :�ۯPN��M�x#�y��)jD4>�8��q�Rc�J�v0��1w���S6����G�f��g����m\�.|����N�o�ɿt[X$Ã9~�R���$[��m��zj���C�{֥�o^_�d_\����O	:���q�����=]V;+O�o�iu���)<���Ł7��֌�ƣz�@
�������`��Ud�.O�����ά��nL�
,�Nlr�Ӻ�,��$kq�6�ݶ 4��.�ʻ����eؚ�|�i�Ħ�hܚ-W�&uf
��A�3�(��%vQ��e��Հ���鯜V�Z2�z�%1QC�v:�V{a���I*�2,���;ᥚ�|�0�B��lYe�hF�<`	�.4���6n�vC�I���G����5��`�%�vۀ:o�!u���&��MfoH)1'p����>���D�yI�ёNV!���5�GI&�M���#P��2 ���ݓ�OB	��SG�b~i&Y����,´�$�~��l�f�~ X��6�~~�-�a ���S���b��U��:~ǥ,�#��.�T��m������ƽ�������j`t��D�i��} X��/��sS�|z�'<W�d���:�9���mW��$d������S���i�[�[=6c�e�[�#��I9����yZ�[o��ع�0ۄڕ�(���^߇eρ��z�%
����W�%(�.�w�ئF���6>�|���_�/π3�]Qv���ߩ]\���
�8"�8c	p�,H_�68b�Z*LDo��U���՞;������ZR�^�����_�����{�nK/)$�ƀ5�LxM�&k�\@r�����xE�G$
��	�y-��ޅ��pp�u߄��z�s��va[D��r�� v�g�m��I����1y=��)|���YΖ�w{�kG]�	^� ��m�Hs��g��KC%�y��)�\��?��K~K/�\�`K����@�A|ι��{�c���|8ا���ꔝ"�JJd
O��[��m΁��֡e�p%�N��C#�1���'l�r�d�f��T�$�>0} 
c֋ː��~F�w�W�O���UA���q� ���p\L�����${W���3?LMe-��8�[�ꦙ"#�VGP[5v�C��)a{T{�#��e|�h�6g�w��������\�;�����r�qڝ��k���w���\'ϲ۞�Vj;�K�U.�~��w���/��{�$���h���"B3�9���vqC�6�5=�S!��l��e��? �J��;�x���4
���'#j D��ױ�³Ւ�h��عd�gxƶ���.CP�@�l��j���n?��p�*(�0@d�מ�V�,&�$�����Q�2b[��F�Ɯ��q�1$&s9����z@��wm�s<��t�(�^�!r�R(�����S��	�O0E��B�ᡖ���GU��>}��C��{�ಕ/�[���a�Zr���+q����W.������v��?��$�&@�mUb5���R9��n�ިS�%Qv��jH��+�g��?"�6i������:�%\�0��,��Y�v�۩���G� 'I|�N��1x�R����[��`�$�h^�p��D�t�$���7W5�Ƣ�*~%`~��i�@k/E��2&C���~�tU�w�����^�Ė'%�YSH�
6�Ă3���*��R� rL�r3��j�rb�U)�H��%�z���NS
Nl �]�NV�Z�]Ё����6t9�[�ܧ `��*DC�(_y�Z�����h��o���\�	���L�[��/(�8�dV�!2�6[b۳���T!��;�Ɵ���o���"�Ǣ�m���>���ݥ4������L{6�M���3�	������]��┎6O'Og=!J��
�D�S����� �o�h��Uc��J{O{@?ߞ��>�)HΪ�����I�_�����ʧ��V��n~�SBz���[x�G~��$ {V��^i#��ð�'�@���7�[��*��K]G���դ�)��%�d ��9OzNA�s׷yf0�'�Z�K���	�ٜT>��Z�_'��I�-F����)+��S�Fkٜ:�D	����ٲTǜ�_ à��5��zN��v�\[@R*�JD������	D��i��:;���Y!���[���]'�4� /����s�6_s����}�1��^\���5X�ց�k�I=���qu{�)���(�x8��]��D'ڙ-����ۺG}�GMS��~��`��-��D��u�	q����������N��pF�u{����i�~0\����9<�������e͍��qo����H�(�����ڊᒁpwD����emF���)	v�?4a~�����yք����ƥ�b�h=�P��&�� q��*����m|��N���������Yqlؙ�qUyȭ��s䑃����GRw�
Y3�}녝C�:�_P��8tYH�v~�u����T�Y̫=<,��-��T�A�3~\+n7��,�x�f�q���	h�b��� DZy�(Q���z�z�V���!�뿟%둀�k�r������ � eU$�wel���C�J,WR�&5a��u�:QLe��A�`��$Q֟ާa*r����C�ҽ-�9�K�+�	e-s8�L�Q���6U�"�^�� � ��G��|��?v���d��x��N��nM���~JI��i�!G��/Voz{�cN����_��]�v��q�e��ɩ���q�jܣ�>3��s�I��O\�s"�]TF�k ����?�䂒��чq<_��X[嗱w��(%��2%�Y��|����d�'�{���.;6pg�1�D��t�2�)¨�F�PL�!�O:��b� /����1�Q�W�(��|���T�������*�
j ����*��xnsF���T�BS,��`L��|vܡ��~(�p���v�/qa�'���gw�\3�]��?��3����=��]o�qex�n�a���XfDS��)nPٮ�%%҆y�UkL�S%�<D�����a��E��m���sР��o_W��x���X��@3fdx)A�k2:�g�Q��Q�����a�\═Wx�I�����j�+Y��Tj�(I�����Wz�`6R^�}����豌,����52���E��3k��qM�>-sG4��r�),/D�ߝ�<-9�5�uJ^c8�0��#�����sv?+4Y�D�-��S�$[��&����F��f����cъ� �>q"w(C��%ʕ�p����r�g>b�*j�G	�����,*��ny�	)[�ڜIr2����f��	��I�\����vz�cC��;̵@b�Q�����SU�ק�X��zh��u�{��@΃����]�/�0�#����e>��T��Sȑ���]!��u�@��E[�j�ץ�B_0dCz�)a�L�PjTjlzB�x�!�4�0]���ɹ��JqBU����m����v-��cX�4br�t8�c7�C�M�k`�?��(��><E�������?��ϕ�� L��[#0t	ȿy��캨ĺ�FТ�/2#�6�P���m�]%��>������y�A��mc��5C^��d>e��/�q����:f�Y�Cl��S�pz�(�Y\]H_���X��F#' ��X��LX����4�Ug�ހ��Mv���RJ�v� %:@Ĉ�=�f��f�+���z��]�||,|�*˲R���?�,���K����˧3���^�0����TO^g�a'+k�K/5����]��]/��3�W+���gf�=�8�E�V���zލ豫��z^[F���꒗�У��a�dg�x�!(d=BZk~�F��x�w�1+��f4op9�YϬ.� �AZ�e�PS�S��`�5y_�I�s�!���"9���j;�:�]��j��=
���^�Ζg>���qԑ��It��H�B/���<���-�*i��'D�gt��=��E�ظ;�:Ȉ(�̱Y����H�������� M��+;O'ٗ)tC���4�9Yj/j�4���X�J���`C��Q��쒟+q��!`�D�(�<��p�>��8�7�)g�O�6S�P\ңl�<4������4b�E��Q���*��\�*+�X�'yU6��A*���-v��ۅ�}�6/�A�����aB��^���cQ�Fd��������2yh���S�̯�Wv�Gl����t�m#oᕀ�1����:�6����笲u�v�N��XW��|��Nɉx�N���U�3���5���}*��-C��b�H�	�����ڍ�x�H�W���m]^n��.D�7�����So6|�;:�_�o�U���t��BHU�\/DJ�T����6��nqN�Ɯ\��>�od�5�'<�W��hc�y��M��@Q�u�S�a�ǁQx.��`#4J;��D_�U�p���&5$u�XvQj�L�t'։�o��D�U�i�1����rME�RMUN�eGS�D�fN1��60	Q����J-�$��S�t2���@�2Һ��f����14�HtY�}	y�w�KѓG���j�ӛ����P:/�����4����g�nb�M6_�(���@z�)I�gb钢�zMb�y�8Hf��=�[�φ'��9����M�~��I��EU�ꝴ�-�7�)���֬ ����k��d�Y�:��0&P
t�DV*.jT�<�<(�?�ա]m�DE�L�L�@���M\�ǥ�����}�֭$�������D���?I� x�`O�Ep�7��|��W�^�F�R��Q*^u�%UqCE�ѧ�n����;�{�Vd4LV�Ы��؞Kd�/�D�s�M��V��yiN���#�����T�ې^��蒐d�8���?'��r;8Ck����^Cw v7�����nf�??Y��Oc"����b���r:	3�����H�u�N�*��S�Cn��ѕ-��?i�����a��0l��I =��9��>���%b;8ĵ��s�1a>}����-@�Aj�X�û�
���:2jq��Jt��ܵ��<���������4��_x�˿0���iX%Y� �@^�="�;
��N\v��~ui�T�}Ȥ霴X������>���X�Y��G�SjB2 )$w�
���)�� ��5�'1l�)�6�
r<����!�jw`<�!ǥ�ZP��[C�dǛ����mⱳX�`1�
<n���횴������_=}9�6,Q�*������~M���ٱ	g�q[��bS~n3�0J�иЎ��\e�b!ZU�KE��p]��]j�������U����{�2k�E;��\�&�oՏUi���(�i��k��0�pzt8���:�C����ԗ����J�s�Z��1��[~��y������W���C9��0:e�������b��֛���q5 �g>"�rj+֘	p�r`�@�c��B��҇��R4��X�o
ߺ!H��f	�r��SU�0*��qѻ!��<��YF0��Yz!���ܸ���!Rl$o`�N3w��>W����K�΢���\� u���w��k�9eP��(�=��&6�W�)<�4wuG���C�����a!���#ߘ:L����Mǜ�Xt�X��1�-�kʸA�Q;I�/0R(�퐆�+4y�]K^���Sה��V��ߩqV<4����� q�ړ��2������:���9Ҍý����(| �+�^G�e��v��'�� �V���JK�-My�}�uW&��=�, �e�V{sư.R���:>w�&X%^ �VL|�S���')�ٙ�� ��L<�@Jn�d�?�hȧ��{�oY D��L��v���}�|z�.2q PK;v�]��Er'����8cy�R0����(���;�qc��{��#��[l�Ӥ��ScX��(��ic������%� ��T���s=���J�em<;�)%����
��5�R�����]O��enՕ�=�y�ۨ�;G<�J^	���Rdο��LԨ��(�i.ac��ړ���%�#E qk�/��ê5n�ԣ߆�|�*�7"u���B^^��T�[z��|e����j��;������<Ŋ&$���T���)"�ѝ��&'�Q©XT��7�幗��Y����|r��Ӥg�b��J�����$⯼8�\�r��KLbHھ�&����[g�#�=�_��D�F!K�
����(�P'�1�B=	G{\r��l��쬷#μ%	t�Ir\F^p�C��=�iWN��\�K��2��Q���d"HIY�@��8���K�,ϮF��4�����$;2�p=K��M�譽d�OZ �����8����L���%g^3�0�r�߳`���TT���h���}��؉� ٝ�$����
�L�w@���U�`��	h=���^���֓���_�j�%RSڶ�Ӊm#%�E;�Y���U1:��4��~9�� hTX�_�!61S5�S�oF���Y6��F���?�%8J���������?����1z;�[�s���GS�h:I�Od��P3�^�}�q{�+��9z��_�[-��������Ɛ2%�ճ2P�WfbQ��\�[F���5��K���B��v�ҩ��B�3�=p-&y]�Nh_�&@h��-�7��1:��_F�<�:D���W-	��s�dz�	4�zi��g����<v���� M ���C��MEc�%:=�YiJ�CO��Wyv����1`!����j��a!r��fL���h�c4(mk���cybò����ى���c����i;�W�}=�8X�N�v�MA��1�� �_^��J��Qx�X�*叭ƚ�����3�h�K2Y/�!��}�J�ns_`�0��RR��V#�8h�D����x�3p���G�e��>�����Y����v���ϒX�Zr�4q�|������heXu�"�xo��޶|��n�6,i�>!���骦��8a <��!{�K-GRN"+�fdB��4��{ޥ�����]�_�u���J���%����������S�N"�Dt�T-&�ԳT��8#׸�hʒ3h~���u*CI_�NvPh�7�M7�
臄ǯ>��\��!��+�R�[B����=���[��1q�5o�y�lN�q	�d_^ʵ-�Jj�=��Յ����iy���DŠUh�6g�n}s�W��Ca�i��YA�C��^U��3),�L��X�K>R'����m�����RO��v��w!���д|-��u'�P)�?SuFہ�����Bq��.�9�\�TGm�����T�X��j�˰�T���˾�
5�C���?CX_Ä�;����$t3��o&#魮X��`�D���J�-I4�kl�r9Բ�U���l�z5�/>d��%�6ID�a3qfg@��uX�����$�5�v�Ҥ�����l���ӣI�{���s� s����F�F�6�X�W�T�Trm�����T�iR�#�Dgk����,Z�3�C������an@�dԱ�A:���c�1'~Dw����ߜ �[e?�Q���K�&7��4�6 �(��Q<8E�`������)���I������R��QH�j��my��U �L��u�Ec�f��Ӗ`�Ii"�;�РL���c K#������i���W��*GI�x5S��r���Lj�n��ײV�+������$�k�MFQ.~]��,�]��!�B"����P��') �<!����1R�2�r�F���F(�~�,f��͌�>W@������[.�w ��#<��8\���E(P7�i�=��W�2��󠋹�H8��ی�������A�A���5'a����dI5�B����~9������z���r�s�\~�:[cB��kޜ=Y�Ŧ���ct!�+��M	O@V3�����\��hh��{4�+WZ@���ٻ� �v�y���
��{�AL/'~J��.cܷ򰜋�aM�m�B��,&ML3e"V�x.ЇM�H��� g�͏boU}�PZ�Q�o�g�N��n�b!4��P�O��К�
/�����S�]K����E�=>�{�2gp����c�tH�oG#7�sx4 H ���	��.�-Q�{�M�C�z2�2��s
ܕ+��,�w,�uT�l�s���i~����
���A��E��9� �����*2�f�Y4�{�Fpߕ����j�|&l,#�	���m�;�$,�(��;g�V�*���f�:v��~}�����<��j,�3_��Y���N-�O���\��l�=W��S��	q͹�eʊ#��'���8��s��Aؔ�ɼ/�\���S*�݀,���a�3qMa�䖫�x����ƚ@
j��[A��Zk����Yك�G�G!{��{1��s�w��h�nO�|�=�%�'��;��Bm$9H��Xخy��:��Q�&_[��^�Zoqѹ\68s�-�JCu u�G4{�8�������%�V�9^ǌ�R�Z |�g���_�Y�wt����H���u���O�]�)�P���lY,�fNx�W >
]XSeb��_��ʛ_����q�G��
��Ű1��%���ۖS�&�-�y�(�8�Qf�vškݟ��D,�J���(�~��P���	�%��Tgұ �"��8��̰����.��	?�; �o��xyw *��2TW+{&�[V�9֟1pFY�\�?�k���td�uVw��k_��R?n�Oe%���0�"d��fe�$�=s3�ɍ�4�dÈ�*h`,K�֩�ø��e�7�h� ��r�G��
h�U���e����!�TP���9|�jc�;j�C=7�O���);��8�TG#���� ��p/%xQB�gE9���B/�2��y��c�ɦg��ێ�,����h��M:�ӹr
�i�5;jQ�T(���HSaGt�팆�H�(_A�5�x�������,�܅��$v���Ň}Kw���A�;�iC�����lS���s������Op�\�V�`H��j��ߊ� /���2��_�R���͇W�k|J�i�s��E��PM�{��u$zuyF(R��MC�߯E��7"g-0
����0�x���}ѷ=���p,�,��'P��ҏ�;�a��Je�� c�3�ʹBK��p�����~���K^P�l�T�T[�[9Rq��BE��
h��%ƶ�4cM�ɕ��K�9��q��,ʥ���}l�l��a�:�}���7��Ox5�Jb���cmAu$��3���@/e������2g�mo���r|l�J9H��V�u�`J0I� P�)8��ZH�J�d*�d��Ho��~�{�!��]^�4���	����	-�}_���z����w�.��i'�hV&��j0`j�܊�!��f��5����mɕp<�?�KR�d�췋�Dm߁�D#�yt�2Oc��"��r]8g��]��;�L'FD�������nf��!eW�ĊL�ȮH�D�$��/�8�s���!�Yd�H��������Lsss�6�
>ˠe��G�Zb`��-p&Q~�L3���AF��I��/#�P���j� �߃����W�꽉ZD��nM���HR�Ұ�[���jB
��<l�vDp�ט<�L�v�L>��ƙ�!k`���Q������ ������1 �5q��^<�ܓK��[s�d��U&���!"^`Yh_��qw~�:/ �+X�Ѽc$�^g�n!��'�&�@R6��K�bQ��c����/���	��'v���eD?�v�6^M��^��a�C�Gt���d?��_޷�n�|ps	3Y1��$I��#���4/C;�̘r�Bt����s������qC���;���b�<[A�[R�`sfF^���%�����7�꽒��&���w/��*���7��F��Ej�T�Z}�li]G�Q|���s>�f�m:�&�Uĥ��TwK��E�2�>>Yx��Wx�U�u�}��+%���)j�"��f���)s���X�'�iix�p��8����m�/�F�;����w��"9{��8s��G���g
�ٞ��鄤��a�#%��21��İ\`<��.��F�+:t'E��E(�.��U7$��������/j`;�=���`F�����xO]��3OuE��[P���>v(�1/�O�sؐ�
)`�鋫q�^V�	4>��pE,�훴\[NOn.>��?��LOGA`y����!���ܰ[�0�/�߭�U�i��M�Z.�V-���r����?�l#��\����H���I�nE8Iy���ꈿ-ԇ�y���*�?G�o����TIĠk��<.�y�KF���e�h��w�d'~�_�ე��cE��~ bb\�M�Woe{�CZ8���x$̕�g�����)ir����@( |�d�j`�w6�(n˛y���c��8�qsd�F�]
5t�� �&ȍ�5��&��>kM�5���J?�l�n<�G���?&�%1f��]�A]�k��Y\�L����0w��5��r�ɢ�8�p�_z>�b�����8��6)����/� ;+��[z�sϾ�`��ԓ�ɹ���P���� ��+ϏV*[��& �����h7�Ԧx�= �����Z��E�7�j^��E㯖�l���\`���k���i',��T����P�H�+�@��tpw��ѾHR{g���FY��-KC�h���0�xł~e3i	�Aا}H�*ed����Q�؀�����h�~0���_�}@�C�No��O(�DBϳ�k�i��0pq�tzM��b��9z�r�?�X����
u�I?���k�:���t�l6��TS��kA�V1�Ox2�5i�5j��tN I��#0��Ej�N�q�	;WQw ��'�(1�-'SPᝅqtf�CE�A�����Gz�����r�o9�2a��^%�#3O9c����l��θ��%ܤ�3�D���@����6������a�S��d$5j�)޲/�
�F���w	���BV��xTf��s�/C�k����w�f�,����Ug;(���sOU�7�Ԡ9a���p&�߽��٨(��_��D����|s�(CKX@��z�.�\5K���T
�LB� ^Ys@���؞>��2y?�~w���]��t��F&�5K;抴�Pp�E�D�O�}���@�#�T?-��ɭ  �e�Г�?����Nv�z��s�lO�d�Íc���J��z��񎷇�NP��TE�F�&���#�M��W�=�m���w�~%�*&��/�����,��2UEo�O�T�P7���y�G}U0�:$"��ƈ�l�Q�Ѹ��"�(�Fɥ��I�#����Dt2��L������	��E^L{�I2"�[�Z��L競lp�D��p������m�*{e����ւ�w�
�s bc>x�u�zZ���?Ws�v���!��m;UT)�>��;�h�x/m��NcK�R��W�{U��_��R3�&�%z��Ƨ��α�v;����]�8�φ?O��Q��q"d��?��&7sE�>� ���2������q���&B=�߯U<!}u��W"e�0�wB.e��T �� ���dF��'�����[��<�?�Y�������3��Wj�ao�D�(ʃAJkߜi���xU�}�����$�Xvyڄ�����+�\_r�v'R�&�[�ކ��F5d|�s��lx
FA�{����Y��ælR)������f�'8����C��ܙ8 +B�0)B��O�<t��AYyo��6<qX��7#;��"@��r�7R�.�`yTmm�<rr]Xws�3�H������6\�0G!�?X�Ά���-u�m��xc�g�Q��?�b:���s�y`]�� pM��II_F����<81Y�?tHMC=��W��:�1}�ڥBe*��� �h�M+�@�H5+�gLE�>_�Ri��a@O��]a4�8<k��}r�ʛ@�0�Sq4ai[���&x��� ��8 # ��8Y���7㯹���Q�.�Y�D蟬+��L-dm���ȵ��P*ZW�<S����Ҷ�-|އ��A?��K5�I��D|�1Jw�^��c=]���6�B�!�"����#�!T�Z\S�,6<}���F��7���l��+���x聵k�[���5|���J͒Xx)�6Q$�)�]j����LZOD]G�k^a��;�i٧�tB�%����q����	;�C� %=N#G��Ȟ��3��H�Q����6v�W�"�_��� 	�z�w�T*r�Y�w��Y���JB���Z+s���$�p,�Ab�D
q���_��9�ȷ'��sA�@�F��w���!�"TM��es-1������p�m���n46�����M��`B�U~�HU�{*�6��"�������Iб�EACoi�(����\h�s�J�(��⑛8?۠m��M&�(��+#��n��K�K̐��UV�<h}p������0P��	��^�˓Ar�j*��k���� -�-��pv>�R�PM���@9�3�[E?-�"._�5ǆ��:s��՟Ge;w��!��V�&�<�.��k ��$��D)�¢C�"΁��8�z�M�yH���ﹻ�g��� Ƴ�d1>b{|��u��l�]�0�Y&�T X�Kcy���J�3��e�X�X��V�[��X��id�:%5J/�c^S;�n��~���##�zj�eVJ��	sd���*z�{����#���0S���M֪�|^ìr��+3h**8?A���(�9IZ�
���_��G/%>%[�Ɂ޾�%(B:�~O��T|I�j4b���j��P!:f��Y�^j�w�]���qY��9�	KB;b�w��ĝ��|�hj��QYl=��5%m+�m������Y^�c�ə�0�JFo$�A���%���N���qv�0��Q�į����\_9�x��sf��T���,5��c8wp@ǭܽ�k�@�B��ZqY�M�-:��Bc�3���ï;��1�K���pɛh��e+�ܑD�d[��0|gh�>��]7�7���XOk˂s�G�+	�����F���W����I�b�S	�!��G��{!X��)NMx��^��{Z{N۾�4ՑP�P�����T4m�����\�x7����,R/L�p�E�� �1V}4��Du
���2��mm?T0���D�Xﳓ���|���d��D`/M���us��[G�E����Aqc��oخÐ��5UT�}v��9ڎA"�Պ�/���ݣcߋ��3^q��#�8���YI��=�n�PG$���޻�H1nH�WpH��>�i�\m�u���$�U�0cm���p*�m�E�=nȚ�����	ZE(�ڊ?���I©�8���ʑ��,����I>3C:��f�s`8���sD��~$Dߛ]Ų�I��~WY�ǋu��~����\7���2,�&F��ҵ8�e�c�g*u��ڏ0|*���3�YZ�B+�9�7T��F��44�KR\H��҂{�V=t���{x���n%1�w��3��ѓ�
�:���ҭ��	m,�J����.�g��.|2��Jan[]=�@:|=sYk�KN�0ca_m��r\����҇}q�8�f����B!|�[W��M�p0�����B<������H��0�<L�����7����Z�L'R�9��;�!�|O�;����I�����\L�Fo+-ͽPi4�U��7�����&�q��|� ��1ӹ���j@���2�T�I���ݼ��B���7uȐB��zr\s{���P�]��e�X_��Q*�Og\b�Gl�[���x5�뿑Z� ��y��'�C^@J>f�񺚕Z2�a4��i�8ަ�b�$tMh�B�:���p�1��N�{�k�O��y�G!É:�y��w��d��T�[���p�xL���-ښؽ��Ī ���Tk>C"Ų=	F�_�Z�j����)�B��E���g=b�ʵ��舟�Ç��H�
Go�IZ3]`��5��_�m�Q��;��$��3*�LR�}<��+Y�����闐,�p��qvAf9Iȯ���N�Sfա^��$�J�mn>X��@�%|(��}�������U�ˌ�8H@��Y�-傑�h�	Gb���|P�Z�1o"ˈ�_���ص�����9#-L��� ����k�w�d�F���V}=����T�-,u���ƚ������/�q��+ka�Yd~zr,����(=g�J	���=���mEם��ٮ���,��n�H��P�~6Dn8���'H0��I�	=Q>��w7k�I�J$Z}��*ʿ�נ}ZB g� x��)���Hȳ �ɪ`R��hȤ)`��jn�ɹ[���m�fY0�S�mmvTaJC�eT����8�p���>w@i�B�y�s�v�SèS��ɲ���ģ�����h����H�6���8�' �;#u������R�>к��,NJ��
�@&9�;�(h��Sx\��(�6�M�,��ZW���Fp�7�;d���`�_E����/^Qg�a��#1ڍ���;��^�j���s��Y��c�q��ƐLF��gBф_m^u7�P���Di�/�k=�ڮM@�PW���r.XB%�+~��t�2ͷ��@�o���®H�i��������G�m���F��iH��j���V/
����{��^O"�)��Z��Ҵq%���~�X@+�)�u��?Px��8���v\��1��X������/�\Z_��"	��?i�q��dbί���Q��#ӟ�c/Z�awm^����<�y��ɾ̡����`x��҇�o�nK����I.�G�O�u�1���2�j7�,w�����g�уg�b�,L���q�H*���(���R��nix��c�����\'�R�#=�k�9�>�2v\U?�h����A�7�ŷ��f9�_o*�=�����-P�X�D��3��J���JIa�v'�5�5��<g��:}4II|ǎ����u�ܨ������Ɨ�w<xG)�kW�TǞB�Z;\�RRI�C�T�q9��>�9�����t�
Ѭ������`!�� �4�)�s���Á����_�&��.�jg(N�68��^`��i얧�f��}�8j&�k�Y�J^�Am�K�=�����7��$�\t6Ds4K��qn�0�H $�5����h�]D��S2�9�l������+4b�"y�A}���K�8�ʤ�/�+���جsֿ񚫡�b����e��q�p��Sf-<��E!o/wZ�c�xǟ=4i7'����w����4�	�Iк~�Wb�r�/יnA�z�o�莲p]�����]7&m��|��cۺV�F��|��X'�Õi��v�m��$�v��ǽ[��T��,wz�����.��Ȅ�)����
h�������7>��y]�D�S۰�5�ٞ����H�=6���+_����rP���	U��~8�v�k���0j6�PHk�"Ѓ`"����O�o�P7	���Y��G�UCxd����h�� �ޓ��3묜���w����N����ӄ�誺4ɑ̡�&�!H������D+~��)��R���=.����@9g	�e^��f�Y�n��qҵЦT翛m̂0�c��[��6�<��L[�X�/�N�z���^��\Q�&��TkxD*%�+$IZ�n�׿7�-�{�T���2+��Z)G��Y0�߶��@��#�e�d�1�XV�Dq=	n��Mf���H6�L��4�K{16�MZ���?�f��e���5���Q�4�n�Qi�_��}��<9�{d�м��[Q~�r�౧z��W��T1�޶Bt�ޕv����j�e�b���K@��+
8�#h�`����d��d��͍��b#�|ZC�ub��_=+R�2�	RP���OQ�0!"xׄ����� ���$t�L푲U��g%�SR5�?DY����Ӄ! ϩ˺���3@eFTķ)J�B��Jfɝ:Z�Ҍ_��=��:6�\�>��%�9�@O'W���-����2����J���������^�X��׭P��K<B������YѼ
�`y���DYɴ��'AӨ ��:Ӂ�c�W��u��|y�Wo�An}���
������&�����O���l��ùd-��vR�I4��c$NϤ#�4�"�N ��0t�`���A���(�2�/2V���\�4�
Y3M��(~A86<������i���%Ncj�8N���?G�(Q){O�����j�f�wI�㴃Rf���4�P�{���9��9���Ji���+r�� >���j/��v/ .1{5����9B-׶��-�k��QBH���fӉ1�s���9���(���<ˈ`�ݺ���a��α�
v�Fj"f�#q�%b�/nU;���FEհޓ���%D�0(.�la�z�H�#Y{��K%����'瞮NO9[��!�0'|v+�{|켪�|C(�:�s��gƥ^��	����^���t�iW]���¢q����X��r�����������5���d�;�1g��i$v[FG+�j9?\���oT�Ur���9&]ȾdKf@!=���v�ݪ�R�fx���ݳ�Y�:{���V����3U�U���cx��n!<c�Gc��׾���6�^����	�lb�7.o��,j:�tӽ�w,����wq8#*��*�����������3 u�:Eu���F?١�WoJ@�P�iD:�U)��K�P�I��].�mJ�ѯv��г)7Gz��[�H�({x�|��4�%��uI\L/���s�����x��H[�N������?d���-�@iac����}l�&�jr��,�T���q���r�r��\(����ɦ31cA��������$	Ojn'D�x�"��
b�!�8`g����&P��e�a`�1�qp���V!�l�׹,�=y2��)���~���p�����6�Rl7��ѫ�Y��ֿ�r*6b/W�Fl��q�w���o�>{:�WjZ�x�"�Ee�#~�?���i�	�l�O��q}�7�ˬ�섦���g����6sro#ʕ�m�M[V�{�*��\��bK�'F���<͚X�}�f7�\�"��Ԍ��+� ����������c�0r ok�m����>����6|�|Mv�MM��q��V�y�}^��eѰ���<C�t���S���}����^��L� 椣��|�'"k�.�A� o]p`�y���0���-�/��$��s����Y�QP�V�@q8�����$]Q˻3��o���Ui������-)��`��,��ڮ'�	^�_� wHr�^p*("@�mJ�9��G�̼_�5C�$�3Y��J��={���Jv����-+�Gc�F{2S�:��eH�<"@jnkC�>�,��=����we/t��j�aD�b�Y��
�_�ȱh�����P(Or!�W�}J�I[����O�5e��iO�u(�f�_6~���B;厬�^������wV�u��^�B�G9s���"�Zy��aY����/J�A��y���hb#c����H@��e
�.M$ѬA\�����LbďHFtʬ�1	z��Hбߜ�E�A���/M���ō�E�n�p�
�ms��
0К�$[;hYuZ)�Q2zei"S��:W_<}���=�(��낽<V��fW^XS���3 ,/�����y�`��,�.^b&V���_f�Ĕx��U�}64�G���6�-w?�q�R"�/�z�C�m���Jۈ����bn�֘���� �Y(�G+�_L���0���{�؋���o1;��-�M�: ��^���4��S�����L�g�~cU�b�贰M+ۍ�Lj9�k�S�k��&���S��Ws��'�C66Uhr�)�u����]s�t�`ds,��pě�����bC0�]Ԁ�S�u&ٽx'V��YcZ��18QD7��t�1�i��+�N���ݓ}]�4B��W	X.k�)-+U��2��q=��Q�� +�r&#�x�:K$Ј�vZH�+��[oD�Z����`����q�B?i�o/���6�I�8��� �k�0a���f��Y8_���l�hB���ph�����.�g�<�5}�1k���r�4�(K'8��A<
��$��'֫��e��#�5�<�z�Y���̭��\�:�ͥW�f;�+T�;�l��c	���QU����"J8��&3�sw��!ö&�ĔUi"}�/�Ѭf�C���U�z>8���dvk���b�րf0~��q_�R�������������.\7e�,�`y����c]��/U'��5~��+�nP#?���v�pm��~g�������b@&�uA���`�.`y��ϰh+�X���ym��SB�rx�Ⱥ�L��2��B���11+B�S��;�Lʾ������E����i63�޹>0�G����<��BDy��[�LbB%ͨ�x/Ȉ��RQ�:o��O������m������Z�Қ�Ə����T]" 0�Ғ]�l<��ޮW�}ݝW��RR����;UU����(�e0	~����H��oG���*-��n��*�!j�5��S�9��r�ul�S}�d�������>��b����p��뛲��GK�dF�{k`F�g����l2�֥��8���} ��k��lPY?ǰ�F,>�
�<6~����I��������k�CQ�)Q��=�|u�9�l@�Z��D)XZ3�A�L�a���pN��+Ħ'<��#G�o���I��ڒ.G�m�3a-<��[�0~�����|������>���]%~��	 B�#���)�bw �KN�_r�l������aC?X�+N��r�NU��n�9e	(Y!�ݳnͻ�A�]��/���D3)�� �lyMt��j���O��֓��J�)����o{+��m�+��b{Q��鋜�Y��I�jx�B���/��p�{l����p�k��׸Bꨓ�\�u*ʳ��H8�L^� �o���8�Q�C�"��{� ��w����� ���v~}C7:�o�@��\����F��)���ٕ��Y!�i&dBS����E���$؏l�AL^V/��	��}��:��m�#�� Z\l +�m]�U�[����AM˧D�����O�Ĺʂ�WT�������K�ЍS�%F
{�	�s�N9�x-����U6�R�#�:( ���˹�bXezȵ���$e]#��<��6Ӡ�-_�'aꨵ&��ƨ��;�6�T��Ԫ��yQ�S3���7p�$1��7�ou�Ss)w���2)�3/,����������xw!)���w%ё��rK�9͊���1��o<sG	hѫ�pՇ�tJ&��]Z	Y�\¡��_4E�^:]���m@��;$��,Y?&g������|���L��Jn8�)�����O��,󹎺�=��[�..�h�Y�S�a��o�|�]Vw���o��aŎ��q��·P Φ��[	��J.�A�b`��}�6��b%J�	k���\*���C=n�D�kGʵ'�z���m��M��a��Ć�a3�C�C������D�����y< P�X��̟<=�!�h����4w�'	@|^�#�C���A>��Q�h��ɣ[��*�wxSz5������,�>t�� 	�'H�o�� �꣺�ω6���l�.a��͊��������u0�h�'h��||͆���}9����X�l�&G���G��<�8�٘n�&���^&��d��ܱ?� RhM�aɗ�$@TB��X���YVo|� �^����Ơ���~<��>����:��!&�	&�u��E�-r�=D�G$DF���ιj[�KD����{����͜�g�ل�}S�
��˛�^�ĵi�� %�*6�ؽ.A��Ɖ�?�_VM���WNJΦ�.�m% yT	T����/eU尧�P���fN�e�������t�1F*\4���|�R.i���1* 4f�0,ɣ�%xgn��f�GaV}w` ^���\�tcӱ5R7^ ����M�B<��X�OX�.2g��-\O���~�˿���y��*(5�l^��������P��̌�ܳ��1��M@ڿ�(gr� 'Ӓ;��?��E7���(դ�":H�����2�y	�I���O?��S�|0�$4�&���D���W��ţf�80c�ue��t��S"/]�E��\�Me�f�N6S}�c޸���F��G���f��k�/��6�(|����?8��+��=\���kDZ~ӭi�ۣCs��~6��Jum��pv�F�+�Q�/�a���($�����c�Q�OAB��0H@��H4�y.���)tx0b�u���Ĕ-�a���B�t��?�Fbt#���O��/`~w��I,%b��9!��Cu�����e�@��s~�q5�ت�w�3�E��~0��8u���l#D������üG%��v����Dc��6Dy�yύ��-�hd��KӖ%�t8�z#c���5���P)6�� ˥/����M���n?D���A�cml:���,��t�Ez98�Y�S�����sA�ȳ�
2O�rKr־m��︐�hOi܊hh6N�E�G�OQs�wR��_ �m1��w�j/��*:LS�M�]�$ݟ�p*�;�S�{���T�ͼ	�GW/��a �,���.�t�����9�ښ�0X�����6^ӎ�3���R���<y��Q2 	�����߱�;|&?�9���i�+w�����R|���QN�/Ӕ�����]����IS8˃ĸc�o)����A?d��R��ZY���b+����*�V@[u��#��V�[�R��pi%��a��6Й�(��||��`f�X|˽�[���}��Ƌi)D�Қנ�A�Ȣ��m�3�Ɋ��G��k}��~�'� ���b��?�~رO8�v/Fc�Ml�^�pǪ��ՓN\�����hGR�Z� �La#{�]P��{��轺�y��L�&ކ�� geA=�HSf#`\Z��!3p�H%�
T U�Q�,g�Y=
���V4d|�0��2���TBS����nk��8�QgUK��0��J�w�.}�yG�
�8^��w䨗b��oY�n��y2���ʹ�r��p��L�"����-d�f5�y�x|�''N�]T0.�ʻD�.�|a:�g*,U%�(>J��"����'�jdw�V�_F?Pן�U7�.������t�-�l������y���p��Z	��,�>��7�b��#,)Tf�샕���4{��xAV]���Ƴ �|%\U��B�ŮS����a`�{_���~���[4�����(]>�WQM�W��¤L��%����3cP�䕈���?�����v�t��͓��hEmx}+s�S)BW��$�k@�p0t��_|�%m�'e�'�x�/i/�p�@�C]�ʻ�ē2.J�mR��Gr���^l��&:���&��W����z$C��F��(�>P��U�Z�dxqJ-с���<&�5j����������Y�Ȃ�Md����^#�Ι·�cF���i[lj�@?�����tlԗd��S�lա���]�����V[a���ب�����@%��%PX�5m%�B��[o�a����D��>�vU�Sqn�6��QNdZ�
��蛡��Gb�վ��Yn �-�,M�����2�]}tζ�����i��gg��Vg�v���m7��Ɛ���f�A��a=���HP���A d�'��E�"A4�`�{p�����6%��C�n,�W����@ ?�l%v"��fA)7���E,)������cBS6���z��?^�Ɖ �8�@ԧ�B�,w���Ëp؂�ȴ���п,��5���`�z9���c(O���ڹ	��_���o�,Z�~*W7r��
JTilD���L/6�8���dg��i��	Re|��b�[�&���ND�G�c�.��_b=�k��A�����!�l���"�ӓ:X��|���ÎۦZz#/�Aُ���^�Pث���_/�w-E 5V��i��9�ك=Ȃa�f����B<�\-�B6Q;�	�:��J�fi�כ� �+d~�.Czw��"2��IE�tVw�{�"��!N�;���)�{���,(9j7���4�?�{M��}@"P�uL��7d��>�G���i�i�����i�r�-|%u�jX���pX�[��D�/����q�<>��k�3���& �@�^�1]�T��d\���Yo
�}��v>OƼ<#7���
d�S��~G�&K�~1D�\ �J����p�~���d�X�hΈ�M�ƶ��W�W�䙬�ϧ�G^�]����5�}�d= ,��U�'v"��7�[��%�y����4t6��B�F��ژdDƋ&-g.cEb%��h{���+S��e<�"��Xu!1�W\� �'s͵��i�	�|�(5i�	!c��,_����@�g?�끝���xrN�Ct�ml�lSn��yXh��,��jJEH��ͅ�>v޸��ؓ�)���g�=2�����(�5|�h]q������Ίvr9w�Y�?r�s�!��3ye�Q�8��ҋY��HV�*Ѩv��1��D�/�&i��H�.a�M	�ϩbs%���UҫCV?>�.1�e���8�eb
X���cm)�E��঒��gcH��r$���'+��v�f���Wm����i�������M����g�+�:'�M)-�&~���N|Ys}�u�=��d�?^���d��4�~�L9$�q
0tm����{"K	`�
#�t�է�='�Xg�B2��g�Ɗ��h�P��zP~X�t��>�͙{�S$�8�S��:R.Z�1�9;����maE$�F/���>E~ܞ�9@�]�s��1�ͰB8<�����N�)��F�>�r������w��ES=:<����&�
E����+��˄}�F��"N�O�^��x��1�f�\�4Tn����!,�dV&T�G�����cm2a������>^|�����	���㴖�")y�LF!��@�#�YaA'���$5|�v;k �.��|J�<Q�H�~�b.3����� G ���gZ���Sjk���x�4-y���8�SZ5���܂��?��*�[eW87!������~ރ��V���1n�
�F���9��bҰb��B�'tW����ht���h˪��j%�I���5�vz˫*�Pk�?O�$3�'�u�G�yG##yö8~hu������=������&z����՜�6�}��/����ah�kp0Hҙ����T9>�"6�Ʀ�=/~5w��vϵ�d�3��� VT~Ҽ��?���� ���w��˪���>�*�m�6RP4�Ղ�I��ۇ&` �A�o�p ����7/GW�������$i,ro6n��W�Q��-Lgy���^��C{Qˊ��d�
�jēyz��bT�pr�݂=�L� �����G��D�d�l�r��	��sz�������4�'�ƳN�0�o��C��#]�g�-���(�q�\K�x!�ߚ�����*�S�.����tvw���.E0��{����Nt�~��M�\�*�g92�o�)=D%ڕ:M<����0��gݪ�v�ߑ�t~��o�p�%#V)��C/�R�t�>2��x��X�й���3U�'�Օ���9�K̨t��l���G6��#e�A��Ow�"��¢{������?j�!lE�%�������4jj߱C4������a�L'dK���1��}�&e�4���ʃJU��]Ecu
��}�%�Jajذ�2v����R;�P��s�+1���F�^�R��/�%'�3``*����d�N<t֗�e�2/�����p����t~�׷4�Z��[�Z1�P�le���=��<��8��z�g��^a ���:-�c0�G�Nق��g�� Ѷ�Tkl<�.&���x�E>�|=�9����b��z�s���<��B8k��=�Bb 6u")=4&0�2�;f�)$���������O4_�Bc ϖ�-���u���sn���Z�0���8E�)Z礊y����.zg��P��V��������_*dw���¬Fy_:/L�f;�7C���0J��~�_H�L�W��)��!��]�B6�$��F�U���{L6ռ~m��$pr.י���WK��I����6�c�p�� D�2��6+�~����l��"vy�f�����,�w|&��m�L�г����j�Q�}[L݂s[�	-	-�����.�1r�nhV� �#r�L#4�#@`��]P��WP~lA��k{,Wx�m2I��C~S����P��r�.�`���Y\tn;ܗ'��WO4����,Fv�B�u�����x���ې�W����KP9����9f���v���H��f��x���n��&C!��S}3����g@�G��fm`�J)�2�0'��o�������"D|�&�zMLk3hB�bt��d(���t���5ڑP��7WLY��0N\Y9]l�w��WPyb�L!�8]�F'��?m@5x�]m��'��ae���0��p���L-���5cL�zx!X�y'̶.q�HY�THh�̢�3��R�dt֕����.�ɳh��d.��ҵ���@S��~��T�:ak� ������Ngӧ�/��c]#��u��Lj�s��%N�aŬ�Pq���W�f��A*�g������e�Iuj!�
��ݾi˅�>�ϻ� f	ޗ�%�r�d̘�=\m������۬@,��h����E]>��:��h̏�mlԜ�RW���ٕ5ʧ�$I7$���h϶���=���m��t�)��P�N�N���}�/�	��FP���;��cQ��<��G��d4ޠ)���G3��d�p4w�6��/��ŵ�#5k�HW�{�x��B�c@3�Tc��~��iCy�lE����cP(�g�`�t&���q#�V��ckTs}$� ����(R��E�R�#�;��*�6�)����(_�/]��EhT:����Q�A�w��"h�IE��9���P�G�Q+���5��=Ċ�@���(.��j�3_�f��������M�e����$�?�i�������?A]�Rq�-q;X�O�u�^U�蓱���Je+(|��,GF2�m�>EEXܚ�D>�H��wƤ	���O�Ϯ+=�2�?:�a�{Nj�8��jJ
��0�{R^Z�l���j�I���:�ݼ*�J�,��#��m�^|�ڽ�S�}��l�ɣ��&�,�S�Q�������%�]�.r�X4@W�ri((h�C���ȭ1��k$�*HG8�n����V!��8�k`�i�;���>��D)��vi]�f3���^�c�g˚�~p�rt���&R��P\��B�,��}��]o
����'��k8�V�� #��T�.�l:�V�zt�P�Wq�7vʴ��O������	;������F����N��4��g�J2��Q'V��j'=	���@/��@s�b���w�5�W��""6uF�,��J��!�"p����g�z-��y?�E���-
q�`>'����$	��9y ��S����-�JJW�<��ù�P$��q�w	��Δ��H�p���-�a�Z�d����G�>���4QF���ix��>�~���uKi��+m��w��R�Jه�m��ۥ%3w�p��ǜ�+W�DB ���e GM@��b~T/�GN���z'�¬�)��᥹���	�4�g�����HTfL����t�wEL1u�|K�8;ш�r��3�A�6G�;�҄/X�-��h��h��\R��S��{�1���@Q����AC٨(�q:�C�al�M�$Pҟ�a��ph-A��o�"D����uܿ븺q[(<k���^u��.;�����o2�X�𳟔%NB;�8��L �x�4�{�tt5U�$�j�G�qC�o(�ML�s<���� x�~�j]qI�ΐ��m��m�">��=�(N��� ��e�*�����6��vt;�#�M�ጯU��0�P��@*�g�-��G�\��;�>��Q���m~��8��u���k��݃R�&��`j��E��fp�+E<�c�LfUIU՝�3��dî>����!7��y�"��12������3�]p�㨤�-�p���-�W}R�/�v+ʻ�2g��^[b.>��TX�<ǜs"�{�)������VA������\ ����K�lh��o��eag���:�R�J���Ɠ�!;v��|'e[5B4�$��s7Ʃ<�&�]�|�gك�Lu��į7�� -�qfA��i��պ�_��ُ�+�,�l�&M��AL|�Y,uK�gLo�̶Q�g�h�(9��o4]9M��B�f�Q,��fCK��م�(oHfM	��47��v7d?��0��x�����_�����\H�M/��6�-H6���P��g���Գ0��X�� �Kz�?����X\��.�O$-�vS	��-A����H��`x[hLCUp��v�����Sr��������X���S��1F�,���ʇ��Zu�����%����J�^� ��V�.��*���Z��m7�Wܳ,	��x݄gͥB����2���t4��ڭ���`6B�E-�џ��q {-&P�?ptt	=�e���2�%�3�nX��"&f�?�g��B�P��}��R�?	���8spb�~U7`N�S���NAO�M��5�4�x^^�J���s���v�=�_��b�-�^��1�o�!��**�">� ��/ |L�vqF���v B[qI�G�(&��|d��P�AĢ)D%7q!�oq���q���~�\_�����s���`�_��ob�-����Q���b2�N��هy��M�U�^�XpV�a���}�<H@�����G�<q��q��rđ��=Y "lbҳ��۶=�ѯiJ*7�}u�Ց�	�j��&�]�=�u���Xs��.�XR������;kJ?M<'X����j�S��f����«�{qW)��Oh��]L]�N|��j�W������B�k~�Zտx��H�[�3G�l�Z(#L�������RǸ��'�I��3�����+�波�R\�k��Bl�s���剕oqf���=���_�ޏ��+�|��qо3�V������B*�4e���]��I�|���T� �zF���	�8�k�O̼�肎2�;,��;�<"��fg��V,g�p]F��8v�CLmU>�FZm��ת�Qj�6���A�r�j��?b_��xEy�����\hm�7i�v�
����j�~Ֆ���n5X�o�K�� �1��:32Xq��0��X�(��,ε��-�Kf�
�:Bl��� +*а8����5��ˊ��Y��'�^<8,'I�ץ)��[��b.��ڙu��,䀖�確Ĥ�NG�BL��/3��y��Q�Np��Mn6ϓ�Tj�	���~�,U;�s��~!f�%��Bm�I��Q��E]v��c_�$i���,d���#��	�щ�;���N$Q�PJ����M�P��?�^t�0(.��� �M)V
�*-C���6%��a՚̢$C4-��
�?�����qx�Ҝ;$���hƔk����I�n��G����v9��S���W�*>�����b]1г�P���̒I�cB�\?�]qw�M��E�u޷�F�{e}K�'1��s�q�;Pp8s�['��~��2�R�]� x_#!}��p7��"ӓ�{T"����֤
q�*�P�DK���{�Oi���ҹQHp�fi�����L2j�QN)�q�e�|kL�N��:�
�p�7��+-�s��#��*������2st(�p� v��kb26&��H�)�� �=2�q*C�#��3@�p@]<U��0����UD��'�ʦ\����kH�*Y6��Zv�_���4�[�S��Ć�,���AG�O���d	��Ld��A]��DGBT�q�R#�>��!E��d�n{P��t���}�5��`���lϩe������U�F@Zy�j
�=�xC���D��8��G�[����~j��W����	�bJ6�D��ׯ`]Ჾ�'j"m�ݿw����itu@aK�賝�8��T��a2Y�/�����;�;g'`U��<�X��¼��(��[t��*��F'�Q�r���B�%P"��x?{
G��'�Q/>-��?ڏ���
�t\߽���W\3���]y���S��B��ޑ�s�I��U�$�z_� ?��8/D���}4PWW��N�q�TC�֪�$�\��<Jj�`�J�����0~�ֵ��?9����@���Av�A�[����+!����a3�[�X�|�(����n��pl^,v������5�r4~��?fA�������]�"Z��x�����|�.�C�8�H>Ȗ� 	�����W�X%q��5_�H���E'�άM��+-��F��L*��r>���x�7�9��1��_�۷�,v��Oƺ�GX�5�<q��8�����c)yу��)��c�l<u�J��pC2��7%ۍ�N?�1�ӧ���" �=��W�9*�dm��sX;
�J�zf.�ɵF�l��>�N������k�7`���E��p��Ҝ�M���O�:�����V��xe���n�z���l�������⮿���r�Q8�`��N��4���܏j��?����ܘf&'t�iP���`Oh�'�S�6�w��F�&��i$������*4"׭M�5ՙi�$�,�?u4�	��\��Pw'��*@;��"R��]�뚌;1�ɪc����G�c���)�'8�/TF�Ͱ�+ST���\	�����zD(��Vd�bd"Wj��S�r*uIl�f����\�?*�[��^F=C�g�����!�@�����91���������}9��]����Ëݶ;�,�BTз�20غ���\Qk,�()����]���eq�w3���Do��a=Q'e�c�7 �~��g���]� �,{�~Ѽs����<�ٍ�<�߫2�	Q�����B<�j�y������S���2}'̬t�u�F�����e�
�ծď�)���=�����,��4��iZ��K���s&YDE��U$�Ճ�i��
�
��qW�9�
K��S.΀�e��H��]g�L��O�[�hh��[���a�FP�.Ϋ�Xh,��h`��d�Y�	b��@��Z�W�ӽ��v��M�e;�m��e�d�>�?>a1!�1�<��bT&�_C(Iu�~t�]��I���@���,�1>���;�~�ᘹ�[1]-O9I�d��0j�H��)��(yY]�7��$��W�_!no�m[p���5z�I+Q<0~�-܀��N���rŝ�Z�f&u��uQ�H�m6�?�*^��Qmݎ���j	��!p�w�g.���P��cTj[~�;;Q]�v�99��*NwX�kr�S��^���cO�m|0�'^j�沆ln8o��L�����P���ٖS�2Ը�[��7l$q5@٤-�*��-JϮ�ś�Cs<kJ��2�8���������k����x���'`��T��K�����'4�U��(nR��
��5�^�xUN��x���ǈ�P��1��Y$�����~>�vu)�O�f��z�Z���M��1^��޳Jv�쌆	n��Fj~�����ms���V�6��/;>���X.�i�L��e5�b扁��[W�6^�Ш��:�+���*���)�'�	�X]�'���weY�U3GY�����QC��֣��I¢�6��kd�zN�>�����\�Q�w���pS���
3�~���[Dh�8�a*�l��ه1��o��/D$K�-��n{�"�Ֆ��ƘC�e!!����݆��zZА"��;�����`l��H�bL>�^�4�O�#@r��eD��]�^H�}���X�gJ2����vxĿ2]bY;��7����B ��@���H���(��ԫ�C����A��Tp��Q��u��F�i^������(|		6s��l�T�	e�
+s���;ta�Y�/)��
} �L�:��DW�UHx�R+�4���-����2x�Q�`u6DC�N���ۢ=]t��ف!�ګP4f�����{Y�p<��:�AA�g�����墋C�S�x��u�@�k��B�QkH{�@~`��S����/�(PF�R������7��b={�b�g��!����K����By���q�;�Z�Ih�#�b�T�VR~�������o�ٿ$M���	q���){���۬vF�EYq�RMlQ���1�|E�(��!�n�����l]��\n~K�	�� �ݜ��q���4�݂SD�"�]?n�Vc8\�_�<�\4Wנ����0�Ͳ��c̬�v�ĵF�
��MH��Q�-xl���J)P�U&�l�����~ޱ|z�xl50IL8����Ҹ+�Sq�J�P˔�� P41���wC�l�%8� ������G�׫լ�a�fa�
��q];$նCA5��Ѭ�4�y=|���04�N`�|V�ˣQ�0X$n'�>�ء�S���3ߘE�t=Լ��2��M,¤���@B��$��N1w�5�ԃ�mQ��=��4P_2�&�l ��n���[��in�5`A�dO�m���sM��'���l��W��Y>)�j�� �C��w��)v{���0%}��yc��+`�d� ��)��ѐ~�ZL�2��$�^��6�U�UCȚS>�������/qr�Mӝ0��|4��-{gH!��5nNu��&z�+kf��l�,@�˒���O�Uto��޺Z^Q���*�@\	b �a~��K3K�+7?�O�w�PA��]?��fj��>"0J��~�::�m�8Z�	�
l�H��4VF��w���	Ù�����nw�t(��U��2��kbã�r�7�.
��s�H���@�����ƿzF��B {�g���NE��Y|V��&�zR%�f3���^�Њ��MD����2O%��E*��"��������{�a;���^򖒪�����g�V�F%K)���S���lw4U����s�ɱE�Y�P_��ji�� �5�t�]~C�6�� �$FC�^	s��������|���0�����~:�ǭ��^�,�"�QBTT8��q�rķ(�:ȿ���g���-�#"��}<�v����N��<����DFU��?}}��0����<�O�Y��R�l��n�P���F�Ďud�oeq�;�׫�y!��ǕL���*�zC�m.`��K	�%&�w	���gdb�p|�Ij֪&�6/6�7'���5ij�=Pt(�+�������r����C�[��۔���Y��=iv#L�F�w<Т��'��%��#Y+�WF"^>�D8�ye)# ��>��@I�\/j�Y*� ���;� ��!ԟ�wo��	C�}D��YR$��(-,U�{.��mq��ƭ!9�$J�����Ah��3#��:�8���i�,wmA�Bi��wy�����3w/�wdh��o�Q�=qɍKF_�:�ڤM4P�[-�v咳��?Mv�:��UIr�M�ݰ�&��w�a����_�����^�u���y�X�Kޔ�]���N��C��5�Q��#�����p��rޱ�FM7pNԅ��r������]��I��:�� C���9�����O/C;�qD(UE���3?����i��/�/`���8�0�7a�_��s�R��:������)�Y��h �.z�7cp�NQ�s���^aBV6m�"r:��&�9����7A�2�\ep���i�D��v3��7]ނs��������ҳ��g��VJ� �X	�@c[�ϋ�)�̃������ 3��c1l\c� �(T*�.Wv��ѩ�����y
!��f��O���>|�J�����J5K����A��ξ9�2�8ij�j# �P�"∐��)�&��9%��Nq�a�i�b��JN7�·䏐��R[\��UzG���e���׊a߰�q�49$���^AU1S�.��f &� �0ڂ���A���A��R�?֞]�]�k����a��N�NB�>�{���Hk��Hp�|ʿץ�k�]FGi�T�lu�1�}�F�Qq�,RX���U
.13����~F ,��`��N��e�~wo��(A�V��˻$�k�j�\�c������T�c�EX�tu�^�B|X} m�uNx�	B{�;���R�-�E��.�kug	aZ���<i]*��(4p�Eh��%>�mi�<��6O��N8�Z�����!@7����c"̀�����!Bu�"(�&�$Op�\�BP�����n�hjeZ4�����Kq`m���L_�lq���h���h�tr�*�ή%]��NG/��b��xQ�A�V �^�Q��*���R��_H���;�*c�E�M��3漴j=�K�UfUxj��/oa�������P�Yŷ%\9��[3*B��t�5��k`n��l�M��(u�$�Ox�:t��ڪ���@�q��js�U��h�������/yr���8��M���q�_ 4,\$5?���[��m���Wc��~�F6���%��[���q��b��T�V���kue����65./|8�y��4�R�1u`�Lz��n�1R)4Y'���w<���6}[j�ñ�O�����'	^xY ��D��=���p�i�W�3�=��{�?�2�;F�����ht�K�ŏ�r�E��O@ ƚfC%\��j�8���gs��(�u��ނ��D���_}�Q/��c��ž5A[Y4�&.��:�#&S��W���8���e�Hv�c%��5|��j�F�X���4ҩ�kU9�g�p�����3�YૢHV�Z��_z�7���R���ϴg��xO�U���/���>M�]8�}M_��?��a?e�F �3�]�Ї�����>��e�* `4K�O����*����+�dHm�5!@�r6�(P��B�5���z��!O��BJl�~���ӕ���V�.e(O*�){\�f����{��a��F<Ds�"�?��QȓЏ}��C
�rd �ǅd�s,�U-��g(Ra�����[7g��MT��30��v]�wb)N�zͲB+6��W26��R��_������8!��������vٻM�����1� 	.+�-X���.h�cs=���L?���N�;� ����|��ǋ�<iΕ*K[X���l�bF*��S���A�����9#~�"%�aQ��)3c�o��O��
4Ƕ5�E/$�N���/Uᝎ��5������Z�V��!56���;˼ ��fi��Cc�,�^D;�B�u�Xs�U9X�F�rg;�� ���oZ��������o�N�0�<�����$(��|)����8���y~��-Wl�wF��q���ߥ�����[+�X�"�e3�ґ-� }��kJ��5����_�V�:�M���,A�'��I��$��%���H��#��l8�5�~C�i6ڠSm�
M��c8+��%�b'�����O�����pS
�럐�"n�kQ4F6k�ȹϤ�k[�b���Sv*[B
��v��BN[��z_��^<�<���n�U"e�{+u�=��}K8�;,ͷDW� ^E����F �T9�_��,y4ʺ�Шg�V͸gw�!����b,�9ʉN��`dj��4�h��1�>���␥��3�}V&!��c�+�dП>��E�o�y��O��o�g��/���7��k'��`2�qt��<���M�����Uq>���#'�F"��WW$�C�k�!j�cp��!|��4of�^S�wJ�'���`�s��U�gT?�]����CAM��.�+���6��ӕ�~��4Вn��x�I�GQ�x�Z���HΒ��seکz�]>լ���U#���0���T���|o��������LðVt�3(��K*���0�=V=B���U��A��o��%�G����f%�c�L����<�M���l��(�t���zI>Y:�ݝ�zة�5q��(��I��MyA�S��n)]��ɨj8NIu�6��j�D$p&ܔ��ڑ�b�:�ѕ7%}�<� ���ؗ���x��%�:����f�Y��PZ����c�^�F�d*�QJr��޺����B%��b���5ȏ�B���ڞ[���E?j9�N����!ڍx�]i� +���貫�}�kxv�_�(�E�*��g��)y�*V��O���)!�V�X:
�v	������&|wfŬ�,��sO�� owB�V�q�:�x�Ƚ����s����VA��)���?*\Drbѧœ�$�0�|���9��{�L���`��>{�>+``�6L�������Kn�Qǧ\hX�;�fDO]�ð��+��^����a6����T�R.��*�����SBpb�"(�{Vȡ�叵�oo�����h�-��Aa�����>�(J%ҷ�H�[�됥 � �|99����IQ�� �u*Œ�	����+C�d3J;g��F۪��l֑�J7��U~�A�]�5�E5g���?p�\Vj��\��2B�"���7cK �2�c��l>]������x3���T~�:%���DC�O�6�[e���X��$$%Q@"K,�G�6+\���tAm@�4��6�Y�g'|��rE�(�P�lG��q]o����tE�z�MmjЊ�� 5�]T��%$��V����A�K]��K������1�鬒�/�=��A���_Q=�_%�*��@́�8,,#�)��:N��m�/)��4���
�o��!�K�n}��k�7a�wsH���;��|[��Z�D����.�A-�Ze>�bV�c9�b���@"�~�PZq��A��٘F�
�n�~f%�e���8�*���z����M�3�;��h;�ܼ\qk^n$=���kKi�)$O�	�k2g7�)�к���x�R����D�o��	j3I�������jC_Ϲ�W��o#?�	u��tFpS;���cAX-�ҋN
�s�=�����T�YZ��=������5�C5���iŃ�FWmE���u����W�˴�x�a��q)��0F6���s0���b�S�-r:m60cd�
B��b��������G�!����H������ϑ;dB ����ȿ�W�
�P�D��S�� 8"o���iZY������d�`�['hֲ	���AGWF���}嬼�.�+x�������"����7����V�P�����p�v�y�:�+�SئJ�{B��8��j�[�0��x?��"��S��}��YB�ɒ3�p��`�3�Y���y'���]�9�T��)���g>��e�~���"X%V�/�VI�qa���SE�c<��+q</���0l��X엚����@o��(P��d8�1��b�#�Z�L�Q�u�`�`t�C�e~( خ��:�C��(V:1�&��wM�P4"���դ=�_X�����6��"�3���w�0���gdds@�>X��A�KW�jU�m�#;"�:s��r��)=_ga&�ö���պ��2����8�c��+�&ncVX�������R�V]3?��OV��Fr���4yD.K+�J96���9�:������5��+��+t�e��G��`m�=�$��g�z'�� F9����؊�f���O9^i�C�'^�5�s��*"�p��	U65�'tކ�0H��M{l�ULV��z�����L#;����1ڳ��oj��U��
��I�N�1��Ǽ^�-��f�  �E��+�*��f�C3}g�!��Ѕ4o?��aW�0z�7z�1��ԇs��<���rK_C�D���yr�?�*�C�X�p	�uVλ�	�I`�T��=��� D�f��.�)Y���lՁZ����K����vҎq����;�����duC�Y�?hn�$%�|��[�X�(�΢�/ �Aº/ݐ����V;����L�:���R�)����IAN��ƴ拀�f���ϭ�7D��
�,�������H�@���(�LA#Y��AVֹ�։�}��1��W�UMF���G�g�-�\@�İ�n���6rOvڿ��D����8!�����*�ݶ��p�A�ĳ�N"�myB�����Y�cE�?�p�e��k $�N�4���h#�9ߊ�E���0��-x4�҆�E���p|���}[~�6ʺ���fK��,�@8A��PC���;�-�s��Pݡg�``5`��`����i�SE�v=�CU?]�o�3���>$*�����`���=I�6Gު7}���T��u��Y��o3���)��|��9��+���BZ�W���(9�e���)��[����U�^t%z���s�z�Ϊ���6]�� q���O
��?�w'������g~����6����g��h/M:�qf�=gO�@�1�SƠ��"�f}�}N0�mUQ�8�±g�"��LC�['��9�
���ڧ ���[7�^��gd��ћ},L\ac��azC<���D���-q2(.�S#��/k(ugV�/��:��$�^,�z���t�M��(c\�T��/�n���#?H�)�z�x�Ϳ�d�&"ݞ����~}�ʙ$��5�Up)�O�Y�GsM�T��9f| _�����^��w,����q��,D�}ˢ���\�/p?�B��3'؉xzVRD
&�Kr�us��`�o��k�-~ $N��堣�D9Yd���u|�t?�����%S��x��*w�Q��g�j䳬2h�ݻ��y��T��R�e2����J+��R�>=���-Ѥ|���{�y�����"D���d�|�u)����� �s�,}f���b��`�-\����_� !+d����~NsԴ�|{#4�N�0_�rw
'�+y	���*-X���$����A{����;��b�����S�㴂Y�A���~sd�9�Wu��O���{�j"W�,Ȉ<�NG6ݥ<oFːS�F�;H>��/�N����G_5���E\"�,1���TJ�&�M;Y���?USmFJ}H�I&�Q�E����1HN�8�S2�ݤkt�܎_7H����������$H���%�G���7�gDw����^D�@A�%�y߸�rM7F�������j������A�׬ �Nx|_)K҉6��8�<5Un��b*��<�+H�����H���9��[���(m��E�4b��M���Y+q��AG�J�]F4���bчh�ИXKkrāL� ��	��7X��hxYU�����|�@4��B�@0ހJLmA��d+�*�.�����Q��)�r|�l�M40^�$�"���6g��7;߅��� ��pL<�v�QR�/b�����PMtY�g�߳��ل��#>�h����An!/�}vp�ؾ��x���z�z}M�`/�'���7d��B�>-̈2�8Q'��7!����։�b�uv���!Km�_���Ő��罉��dh��j��x5X(��]�B��d�fb�J05����-��R*��K�}�Iv�u��)D2k0^���%K�'����`ҤŜ�O+K0�S&�{`'��𤦮]P���(� DG�6�-��I5��x�F��m}F��`3�A(�tį��P��_b|!36ޙnb:�H�5��$��#8���=��4��_dG���q����+k���q�X���*_VPxZl����m@	�.�L�i�BKu������&��u�BAKA�eQr4�L�q�6E�0���]l�1�;�`��GO犞�����C툘�v����Q�

w��\/��H����^����Q�c����q�f��Z{Q���Zܒ�V�ý�K ��BmB!
Y6��&�8���2�_��r)��>��6RBĥ��r�).mj����@�F�2��4��cAy�,�DQV��ī��-0��:�h�
��-xn;4���0�NsQ!>����zh���RI~+�u��RҎK��x�P��6�i�/�d�lu�j�Cӓ�_��v�${�0���"�E�����p3 �0 ��b��m����>he4zz�q�?� �r����|�vެ�~g���^LK_�.�@_a�P��
�����Ȝ=ʶM�9@�M��Bb�)�Ƭ%L�XAߌ�Y=�~��������B�����G�^5=3*,�zY������k�-�{'$$r������N�zR�+a�ܙH�_28	�V#[.b��=mU����8V[���Y. SC��H�����DX9� )c�F!SRY<�	�ƨ%���!:�y� X�m&�OJ�J�;nK�1��q�It�3nG��2�c���`h�b�Yz
}2�5*�6���+B���D� ��.:=� �ȨL�mU���B=+�����*���~	���2WQ�Ti���l{-!�,��^D�ï���vwV���Ӂ)N¬���z� 	�� ���˗�k�ё=�m^H��af;7tl;��wiz�Y�Q)���܏�I<Y�eB�O�Bpy(h�����®KHMj���	�����N�T>���/�����;(0{����dO�m�nXi�n<�OV/�ۏ-�9Wn�7�ۂ�6�&��J￐�`�?��nT�*l��7�.σ�%3�U��y�5 >�N�
���?dA.��L��O��'�t�6�z�^�
�ơ�y������<��6:M�ט���`\\���W�+R6[U�}5i���m\RJȚ牆��W?u:@��DW�^���h�g�vF�������l1�՛��l(|�"��y�W�g�c��F�u���������~f�a�w7[����=pzm|�g]���~���jb�+��U�3,Yh x�8h�v���J�[��v�	�MR^p�W梷yÁ���^}oW�%��/��ʦ����}(ΦK���KH�("uig~hy��q�A�I��^(Ȫ׵��[ �9݀#�Un9��p�l8������K�t3;�Ph	R����>ΞZg�=�U�J4�i�V�b��Y���:3-����1�A	�,��_ܞ�����TL���e���Eg� ����~���J3�k�1�.����X��3k��t£�@M0˥0�JrlJ��W����q�����2A��-#\�fdRrbF��k��|��d|���[x�*�L)B����<	��c�r~��I9��Ė�0�(����g�n�L2�Vl�qU��YZ���CM�lmF�C�9�#�Fׁ�'��q�䞗m��X@�Ҫ`�d���|�*w��hC�S|m^��3���Y@�6)�ȪM���
eWbI}����~�PHV��˦���|6�(�x1pO�N`5���9X}�����?G����n{��~�_�+�0�����j��,
	�x����3�런ڨ�0���)�YD?��"�U��C�pen?���t�?x��S��&Z��[sdiˈ�JY
�ݫ�����(kgJ0��V��a�r��zp��P�\�&ykF6�Z���g$R4�Pzh������[f ���7���^큑$_~��\r�F]�e�p������}��|J])�k"j|���H.��6�n���`1�r�]'R7�3.��9K��&�2�y���H��0]8�"��+���5J�P��zI%������=��(���V�5�)�ْđ�~n�����p��ւx69Ӯ���8�J�ی����j7B',�v�׍Y�D�&�����~D��~M��Y	TJ[ =#J�	�䍽s7�3�������5
Uj�i�4��x��BR�%�H�iFþ��/�)�|�����TP���[q2�p�ę*	��g��c�r�ˊ2��+M05�5�I8#�-8��[��>e�+�\�TfgEvz�~��"�{}�=����*�����s�o7j��}|��=V��N{e���N�B�v2Л	����0�?�6J�(o;�j{���Pv��� x�|�Spx��z�'�<�D���?)�}�j��'P�3.�]�&�} I}�5�h��7��x�?�ڊ���|y� �nH/�ML���.8f�#yZ�hտ��֚�^���ׅ�o�ŉ�$��U��AJJ��v�k>8
�/��8ǌƐy_���S��-U�m`&
*b��g5C?5�!��N/�<W:�H����xd������#���kO�J4@Q4c�1I	HGGD���ǸpQ��>P�-KX��,bϿ-桚+��O�=�(�컑���i�˩d��h�Q6d�te�2�R?�rVn���/�r��d�g�i�qi+���:��Q��)�Ye��Qz��X����.,
�~H�߮����8c>��c9��䓧0K��#���Av"@���l��L�A�8�\�X��yk �\���yG�P�b�4�$	9-�S���I�J�F@|~m�Z�7��b��Z���8$��q\݌g�AG�����wr�s�q2��"�}��ح6x������=z������ʺ���,�o�����"[��`�W4�ڬ�z
Ǌ���4K�i����ϙz�z�y:���{2w�U���ȑ�}9� jL�Q��E�ط�՞�IlmW���`iX�4��ﺧ���Cj�+h�4��A�����m�ݴ������#���拄V�ۺ�7�X��SޘQـ�;��.Xꠂ$�:.ۅ� '�3
h���.�R�S��eSv�ɝ������cL-ؾ)y����R�X�λ�n�C�ާ٠=Σ��h�J�|��f	�j��2���J�f���+b{�{ʡ.� �m"n��{B�M��T�(8e�l�+�dU�x�U��	 �=�d��:�dɾX�Y$��� #�I��N�(n�w|G��@���FE��=�㠷P��z��*ӫ)㒲�����":�_��i�n�jh���>}�o%�A�a1�4�n_�x���({��=��b����Np������10������<��g�WO��G�^I���5p�"<�qj����RH��Q���4%��$;�����mH ��"�Ċ�Y�gU#���a�|L�l���� ���0���Zp�|%�ɒ3c�PjUkIO�^R�I,U1Z���i�L\�<����0������Ǣ#�~���R���o��9�DR6�Z{#�4&�4٘����Io[a�}��#
��<q
.eݹ��^k��{=�Q�'w0F��bⷞ�z�8#``<z��<���JCjv����{3�� ��P�ZL~�� ,��7��h \Rx��K�i?3�.�c}1���pBWCő�X��H 骧]>�*���5���aaFi?£i���"��iP\�@w���I�����
�rD��s]õX?�ޘ aj*�_��1�䝄�r�-�����o����=n��F�ĭ��o�U�8��8��%�aE��W��W� �}-�b�a�8��[̮'m��V��6(���	�-Ί�p>C !�X(n��mMΑ����|���խ���KY(iop���qoc��-b�W����i�����f<�&���:iUro]eY[]�� C� �߃���O��;d��H�W���.��� ˑ�Ac+�������d���@�S��;��${�j~п�v���},s:Y���beܹY���V�
���R�T�v2g�jr��37���4�� ����g�oE��Ů��CT"�����1c���K�jrջ���x��T	��b���4v[��da��h�U�'�E�fPLs+��4l}�yU�(�1q��P�<�[V�Ųg��^^��U{@��+�W��9�~�4���5����u��X\�Mx^��9���ti\��7^���I�����4#�8')�p��~��2��'֯�+͌�G?(o��o�Ɗ����Z�+*����L�&LZ2���iǗ�¨�vU4����V�% �����<;�㏆����p���v�V�:�0����]�W ������R?}���03vه�`�n���4=g�:��X��fg�<eM4�Ր��0t����9��MG�����6���ɋe=֨T]������S/��]_;G��;���,MM��?��6e,E�AEd��1{kTW[cOۨ£�`�!��s<l7Жo�?3-�=��m�``�ne����g��
�c�1��v	��k���t留^��)���ʉs�w�Dsff��&	r�^5|��L�S4-0^�o3���FC�2���#�8-��J�;��D�`�"��M�:G�n�����ٿ���4��ӯ��ߐ��Yh�/58孿���r� ����RE&r�u�. ����+ށ]Q��pͅm�&k���@!	�Rw��
b{�.���th�S<= �"m���MZ�+̴ȓ�92����q>�<b�X
2���~�G�54ß�}�t*=5�!�줞��}�z`e���ɜ����X�㤉��&�:��e_!�O�	��a��Ge-iWڒ��/�S�A�]`{l	�v
$�PϿ��v#щ�ި �x��!1�����줡��sS4CVWfDX����E�mgz#ߔ��	O���F�.9�k$݅��@����r+c�g����t�	�W��7��вx6��FIՐNIT�r$���}�qP�C�[r�<m`I'._�3#A� w�0B�n1�Q���<v�3�bY �1�ݳ_�_�y�h|�Bc��x���QoY
Z%,{K�W�/�;��O�9׮��´F�|��qh�r[�;u��G�c�X�)6�i 68^�j�g�|P��R)@z��0�4v��,cvG��*ɳ�E8����S������腁vjⴕ�I���yV�����.ј���`|�^�I�9��n�������N�
\iG�^=������݃�Ո�����7��ӃFf�4���G�@�^��">��s㫾�=��;*YcO���!3����ޱ�q�X�&%�kR/�&��h��1��}�������X�l&�X8�ڑ��q�?���(��ZJ�Mp�m���aoG����,�.~@�}m��Xb�aU��n�k���nQ��\��D?����>�?�IA\e��{OP��Wb�j��SB��qn� ڽ�p���%��"�)��x/��_$<��k��y[�Ӟ>>��S�4��1y�ŧ���^��ǧ)�b�Ln�i$X���1CrX�V2QT#��_�g��C��D�0��L�NKPu��Uj����M
a��"!�x�74�6�H=�N;�4���bc� a�p�C�,�+۰�~$��.�U4Ǿ��s};-�j�������e|*�}dO7I��p�Έ������m����Da�2 V��Di'v�..=�R���������c��)t�.��|I�U��Hu?��k�d��P1��h�Yya�ɒ��y^!��S���u9�P�-�$���
A�t�ap�Gp1]:��	7���巰~ee��C��u�F�X�x���ve�-���1�0�Ф}9mu�ǰk(0�ޫ�j���w��-�<2*��x�kJ������B�����s�1�S�&T��e)mZ���-���s��N�&s����r�{��\)�:���h���z�h�Yy�Q��lM`Qez�l�%v��a�w�o�'w�7L��E,��3�X| ����).W&� �c��H�4�[99��}�2˯�����o�]VCr��{ŭ����_��nt�52�&lV$�?Dң��<s��Z�RpB����H�HT�Ǌ��$��1�oC/>��䑳���3����'������D<���I�p#o�.~>+�["[�O�r/�W�S����	+^�%S����x�RT3T��`x DoBۑZ��%���g}��)EF[�/�2܈�\����*�m�5����̣Hv��@�Y�ˍN(����9���`��{��;�jK��+ ]�M�`�s�%S�b�#.�4�����Up�}�#K]�c�T�ʼ����m�\����Wm?�o��2i�E��k���~֟���[�`fP���D�2F:%�C�y:�[ǀ�]%���>$���|P��}���.�h��^����C����� ��ӯ�թ�Y�y
`�d��CL׶�W\ �+���#V��ٴϥ�.�[��֛t��椯�b�C	����?	ѫ�.�y��2�N!h"c�`g�����|A���mV��UC����������]��� ����h���;�i+2[�@(���}p�C��	3�錱r
W��ʃ�Z��U\�<|��K*C\Y�xPG�H^�[<��)]�>����tv��v���,?��_��@����U���ՠd�F�س���]�	�>I�I��][����H�J��1K��ռX��;+�>��
^���rE)�}�@H�ɓ't�s�~�*N!M�
[!T<^���w�Z�N�~�|,�~Zkb\C|��7�'�f���t�F�ө��O�h�.e�qQ���������*�=H"��>k�ȋg��)�{�E%�y�FcF��%��6��������W��C���8�F�[qc����*|�҂�����l��E��N\�����D/����lw
>â	��0ޔ��S�}֓�p}ΐ%h�F��ɕe�/2��ʣe�8��@CDb����<�{��3�̪��L��8�OtA ��Uw��S���1�K��ݼ��!�ED��;��O�X��9*�e�X����k��@��9�\)��Gw�Όu�u�A.<���.�8���
�؈��H���\q5{"���KwJ
j�?-&�[�?b�[�"����Y�>�Rx�531V�'�]Ni=C~Y���gQ��i�4k�u�g�.�J��FL<"�����u�t���p��5	hx��e�p�	���TG�|T�B Ӗ�`��M��y����8k6�Sb�ω`4�!��%���e,{�7j�0@F�`ΰV%�I��W7��/�C�K��+ZM�g��<��gd��� �\���Ў��	F[1�"�NƔOB�F�#>})�5�� �YFs��4�G���Z�^�!T B ��QaA�5C����˫��Q��j���25�e��y
�^�J_�<���aq���[��B@g�������*�^'`ج�A.bh�L��/R��p�MXԏ�ܘ)�E����i��?�_q���X�������� �5H�,���)�w����Ҿ��F��u���}fk�z�F���WU�I�r�z��D��eOo9�� /���?�����AKmzq�s۝��/ˡ*D��2�-�T���\�C�G]��3�F��������Idfk$#\ZBC�d��n��'L��w>p؈>����ce������Ok���<��Xē
X'���\�.��}	n�k>?��6\�X��?ȴ�#��x��/	������\9r5���Oֿ ���B�N�Ă`�������� 1�{�:�(�Yc�`�v��0�W�G),$LB�]yX��?>���ŏ�-����`Aʥo؅P��ݳ�b�����Bc��R7��O���,��S�I`X�Ds�SG����Ru��j�iưր7^Vh#A����nI�E��!kn:�}C���X۠��>��2y>N����o�H��~Hk�]V�<X��:�"f��zb��ɠ��	���*=lM���`��$"G�A�|�"�G��vC���[� ��`��5dUs����f_�x7w�_]S��B�7Yv?��]�_#L<e7r�0Hg:B�S����;-����"�� }8��&D�+M �kM��_z�f� s�����gUηi�O�1��b�7��F=�H��g��]ԫ�)j�؝h�X�C���ᖩ�q����5T}4�u������5�USU�f�d�3��N�y=s�TwL�Ԣ�������3v���u�Q����C� ��8��;�9���`*5a�Zʓ�:��vo�^��7�W��50eA6�A��y���[�Dt�o*�ϰ8�8+z�i���~�ų�3�y�}����OaϜ�c�������)�)!��j�sy�w�"�AffX9���s���?�b�rz�v"/�-�r�s�G1!����ŏ���Ŀ���K�>��t�y�R����i�E
��9�/����̘�I������v�S��\�u�77 ��=$_�8���՗i�҈�#^�Z3��P��\��1]=�FxZ-�Fr�k7��p��;a�a,S�C~=��q'��Ռ��%�����͐�w�d�BOхc��c����JGz�e1�7�"L��g'��PYP+���²�$��(aMַ,���h�-ݙ?�z�bC.���d.t�︕lq����&�­���X���,�0����*�W%�h�����0��]�x��lm���m,��6'�DOFQ1隿>V���B��� ���yf��G����=���{�'m|c��j�ys\��E@���6d�b�P���n����ё����Z�n�#B�a�T���"zE%�WT1nW<�"Qr2�D�xqi-ǽ�>�_��"F(_�A�&+�^�Û�(���(I�9�Xnv��g�tk�b�gy��UA����0�qo��ω��jڣ4��l�Q��K�q��]�V�2qS�G����e���ʣGC�b1�v����4"̙?����,d������P8ᗂ��c�I�E%�B��2a�U�[���1��Z�j�`b��Y�Ũu�!4��D�j������c/���f$Y'�+2�r*=�p�ߥ��` ��=GU$�6W�B[N�S��~���v�s9z�S�[�`e����:�>Ѓ�.�f�_�
O4j��C��"��c���>�����2oSبUr��
����o��],V�:�Ƌ���Az5~Y�i*-�U!V�I��P�����Z,#�g���cU���C�$Vz��Q(���.:�#@�.ʮ�蝧���b�T�I��y�i�)�������;�l�8ֈuk���)	Z~�y�у��G���Dv��.M�,��ʶ�F��Զ�v)MEc�p3�i�z�E8��l��Ll	�f@&�H��5r����9�H�@~.�ou��3�b����L��;=W]S�WkР�]Rץ{DT׀ڳV�Zp��l��|��&u{�u�ͮ�U/qg
XL��"��?Qr�U�&���,-��u|]qvG#y%����J�
����QR̐o�%E�`hL��pم.���>K@/<��v�#��E���k�VbTq�}��6�r9*Jy��"Ҟ�6�QЃ��yg�h���V}m�Q��e#�`����#�Wy�G�T��U����s�M�M>ۯ��W��BV�A�\4�`��Ű����+�b� ەa��͍����A�*���5/��o�{��G����]<�m�Ӓg�8��T�fڸ6��'#^�7�����U<����xQo]�R�N�Z�'�L0ǰ��>�]��:j.�5��3�c��dK"��r�u�\Ԁ��4��Hvn��2��X�:�Vu]Qo�ޜ���3#ǂM��n��(�����K�q�X�Y�����m�Qݍ�e�2�C�Y6�ޞ^�@`�\Nd��B�vPwm(�,�ܴ��u�wύp�>?/�I��̲	 Jk�lM�q��d�٥����	�(��g���Lr�&�,��"�"�/����ʑ%ج#�琨����9�v�,lE�J��Q�/ 4s5~����܏<�s ��� p9α����i���z����%r�,�&���gD���/��OF,P���V�bL�Ow&��'q�2�m�5Y7�s�\�����>l��g���/|�i>Os9=��IYx��R�b���7h���T0`Z����O¾p��)R�,ӬGP�n�����[�z#x�.Ț4B�y���	P�����FV�S�y�����ā��e|��@���2�&���|:�m�\8�/ЖeC���U6;��cQ�0+��5I_�8�-��n��J�(�7� ��(v*���"��/m�bh�öUz9v��Æ^���/d�#�ݹ�X�1����8��Lh�=bcPH|@ěx��Yxu���[�!���F������@PZ��Ǐ�&�F q�������e"r���LH��jv�R�V4樦Ԣ�k"<��HE������y]z�s�!{9�A�F�l�Z��+3�2P��囝�ލ��~�I(<����;GA]����ēj���vMN#��iV�T#\w� ��3�Z�[Z�ۓ����(�	�E5g6��<��x��ʺ%�@2��ۊ��~�N2��<�p�J���\����3�w:,�9X{h��p0z����g灩��~���A��\J��@�K K�؎V�{ޓv�����W�]�9X�:�0X�#�ÃDd2�A�'O�7"����$S���C#�oݤ"�y[�6��H+�Şef#-��G�$P�2�)�6j1�4�K�<cW��8��?�6R����0�����M# ���������Ŷs�|I���t�1���o�u6o'*@���v���eQ�]��9a�X7|D'�cԏ�~�o��i�1L+˥��T]�K�Z�AQț�>a H���L����;���XcRY�InCXc���`�Kr@�DÂ1��,Y{�$G��τ��v�U�O��zY	�k���L�ɺ�y��F���c	~���!����&�E��~8<�ժU����+"k������3�u��y�E'�w�p5ۚ���H3�V� ���'k�+�
�^**�CL#�i�zX�.'ޢ�k\s˗��Yv����ص����E'��>�:�C�l�B|���ܿ�`�4�>~��e�˵"K�@�ia����B�'�����,���w���
�wG:�p��sݐ`ܑx���X��G[�N<,�9��.�N4�t�����˼6�G�ҥ��]��&�M/R��8�s��)^9�1b����Ͱ�Z(�c�4���Xn��2�T�C9���5էkxv&c�O��"ua�l?/�X����hA)�Rd����r���]U���(�S�,�"�'SF���n��@� �}'ľҭo��)2@K�竄�Ϳ B��;���%������-�~f��Z�H���d�F�n}���y��ؖ�#�:h�ʣ�������(%�z���|D���ͷ�|p�ݢV柔"gl���SU���w崥h�*/��r�����Sȹ�Etb&��E����3���.B4�2�r].�Ů�6!1��\�ZЏ���<s���>b3e���py�s\�O'��8b$����s�*-p`��xDK|t��<w09����i�m�L&d�w�Q:�J��p��B�p5Q`h�+J��I����V����)Δ���ׄs�"�m�wbR�ȅZg�#l٢Wi���Q��Ҋ)��V��_�����Sa��OfU�A������[;�h�̗�͢���#����*�x��aOA[ه�;��]x����<_��Ә�l�lbp��\���&2��� ��gcFqg\���3\*I����ˡ��%^�;-:!��.��q����s{Q���eCX�9Hq��3�<)�^`C��q>^�	ɫy���z�p��t��;^9���#��1�p��<� ٨�#��-:�}�7~@��ቲ�6�"N��N	���n��}5�.�n0�	Z	��P��1ЭN��uh9��}2�t�΀ l]f(��c�68�w�ӗ�<Z��>��}aq.Z;Ķ�/���ʜ(���ɜ�ۥC���3ܤf	
3"M�RK����\�R���:�ˏf�A@���X��̑*�0��'x�[�g��u<��KTW�j޹*�'��I�3Q�x�4����ok�3���o1å��U�z|�kK�ae�p���Ss���"��Ub�������yE����s��	�/^��� �cjXHk'�f�����a��f�@QF�)r�\9g���N,�zxS���8�>J�5���<����˷Q�'J��}����.B%�F� =`7Pl|��6;h����B>�T��vX���<B��=ִ�Ec��9�x�:Q�mqqy���-�W�E��Ę�����1�NqK7�8���2^`��/�?a��y��V�ɽ�'y���n��ë(f?�c��6Ǘ���zGĊ�T�sP9Ibja����~�f�eI��,�[gj��[E�&��+[{�4���,9�l���NkX>��kZ���aiWMa���>�����?��hzfx�M��T30x�?��1,�)�1:N����O��XA���@{!ɾ%���Z���3����*���Q0)gsLd�dl�Y��"�x�Ť�<Q#��g 1|�PE�[�J�(Z�i�oh��O�;ux�%Y=�Q�s`$X_�h�Rڽ-�-��Lx���vA���I7,��+*I�}0�����"�
^�,��M��C-��U�����6j-ot��V+����x�A|��G�j���@*Kt�~�1](�.��at����@Yڤ`�G0��`L�~O9l��T��H�So� _�w���U����e���=4sF�E}=JC�5�p�f뒏�)�㚞����$0��} �]��	��n�	���mH̪�.\크��G�q�;.�wO�%]��dc�h	�ٳ�*G9��.ghfd��������q ��%�oK�H������p.�͇��	JO1�����tLa��e��7��b�+�P��� �r�X�g��GW+w߿�O)��n3���q0�����W܈-���� �e�&�
L>D.��e�W=	]zR���}��x��q���a��xOr6%j@n������q��ei͕&"8Á�M�� �tY��|�3�6�w�sb0;蚼��6��h����Y���}�tH0ϸ� ��/\�*��2��&�+u����se�!�µu�I��j�hf�1�	��뚵�4�F6�z�'(�h�wf%e�k�	�� �R����
0�������ȶ��Р�^����C�m#�Ύ�@���WΤ���8)�_��[@0���H�R(߬�C�WM�J��}�N�.��-�Ev�I�2I�s��'><�WZ�Ι�T��(\�A�V3W�C�A`&	�m�j� ���]���Y�׏��X�%�\c���tw[i��G�!�gā�$����9P�O/Eҏ@�ꤛ�����U"�-�u��@���t�z�ثg�h�Q�;��)��E��L:�5>��g���Z��7i0��L9m�.f~�K��g:�
��̟cU��.�S�	N��}s��F$�Y+�4f1�l>S�pt(�A����9�8��F#�,zB�c\��p�c�rw6#���x��m�L(Vk}b>4L�4Y�*�3^�c�F���.l��f��dB����VQX�T
���;�&�����@waOm��`�/Ov����cs.��m��5�Wd&�E�f�'Ɛ_W�hJ0͒@.~�=���`Rg:2*f�r��J��dp{�����hm��aJC;�T�Z���(�d%tnT�����TzP�G��_�Jl3��6���G�ЩZ"��C���9ԃ��e����Z��{�ۊ�s��8���m�.4N��jZo]|*~�?���lR�F*!�VA�^I-f����d�~�@�3�JXO���$\���-9�OH���%�(�h����!�6Uu�-�+�}w8��rt%�%o��s�U|�@ǟ�W�~!���8�+pR��؇k��P�ln<
���?#nN�n����������@%n�`}b	�Rͫ���'k�	X/;'�s���a�nQ���duf[_��ԝ=��Ֆ�ȸ���+Z��5I�W�7�;��ԣ�I�j��WH7DO�p/¿�C� ��u]��&���D�݅� R6Mݖ2�GE>� �P��6��z��q��~�,W����B�ρ���ںj������s�b�1��a�_��@%�t�2�}��Nk��ǆ��7ʸ��z�i+��g�W7��@>���дr 4�Xe�ݻ�Ơ}��y;,zk��{Nmx�~ Q՞��{�����W�=6P\Ax���Ӏ�j����������e�:	���@vlr�8��8	�
Z�������G���Q'?s��~�!��s'hQ�#'�nlq��Ph�v�tKc�/��H����� �Y�g�һ���
1���X�W�E���`e(N��54<�|3=K���YBr�V@7�
�+�����x���n#4��7x�w@�s��&/���!�*;�l�(,f�4�Ǜ�ʰھ�����
n:R{:Nͬ������59���o�3����D;�;������N����F� ��(���C�3Zʘ᪱�ơOb� ��x牡��WWT8B^ 5���XX���x��IF_���K�fį�Z��g��l���i��@�a$��3��)����+b����(��|E2�4��>��>�1�-��˕H��wlϥu
W�NW���4Ø���V0�Nj+�Ԗ�'v�*p,��͑��y��v���<�oϞ�*S�\ʚ*!��_1rŨ�g\y^�Ԁ��I~r����?\"M'aL�X-�3��OIXl��Z�xFу��3���k�}�
a�7�6�(n�{�^�WrF?�?p���g���-��SO1��;�K��8n�X\����u@X�{�ֽ�I�WL׵���`���Ʉ�C_��{�lYT��A��zU(�;��,jz�'�;��Kꢉt���/����/�j���T�qPB:z[��/T��Pb6gQ��U�ay[�� ��ޞ�Y����o��?�'���F	��<��6�	)̅;#`�ޟbj5=���d�j���#�#�f�������#�M�V��S����R�pg[���##��pCf�/鑫Ӈ]�较� A/�Z}ͭ�[�qJ%�D ڝ|#O����B�!&�Ы�a`�?��u�+��U��g ����>z������I=���ᄱ$k�)��,7�b���#͢���/<���C�d��&���n��X�ݕ
��SvO`D�S����`�g�^TbK���i�;�sF8*�}�WzE��I�)&�נ��XNeO���I��t*��;d"֠�sm�c�����������Q\CAd�1�_�6u��k���9J��.{�A�< P�2֠����d��C;Y9^Ik��� Ȗdtt��i����v<iL���V�.�V��ZJ��؁�¬ˤv���v�"�\�@��5��c����+_H��kȗ)4��_M/�<��#NJw`�Ņ ;��y��G��/�FDl���Q���z5���f�$%s��X�ഩ�-0[yo�f�K��}��F;�_�N ��e5-�h�S�I���4���nS[o����}��ȓ�?�72�́HOj�E��y��cn �@i�֡�J(�a�}��X[d��p|��\����6`�*���z�@��|"�������+�<`R�B9�?wPS�TB�*� ��㪰�nѴK����.<w~��uR!�\��>f���[[�7�#���mӻ�T��q�.8�	�uk��n~D�.���EV�)K�kA�~����F�9j��,�d���2Ǻp|��y�B�}��?UNGmH�>��4��/�\/Jֽ�l�>_b����\��ݚ�E�SHE�D�
�J�Y���Bd ��e���a���wf�Ō
�&i\���e���%���@�{��)�ןV}�
0�>@^yg��u���H.Y�D�Srj��%�3>\շ���u^<���V<�3�&�r��(����ބ��H(�D�dkϩ���ǧ`���Qu��5��G#;_af-�����suG����G΅,)Gݛ�7f%9�<�/rܳw!8�e��bE�wBi�cj'�h^�m#5#�3 %�c��Q�q{%o��w54���|͵K+<�^GR���D4dp�E7\H1$��f�$E9��uG��H[���J�/T�LOE:H�NfrȢ(��W[؍������`m�"T�	��k�]ͦY�nB��[p�C6���z���^�z�h�5gL�x$�3� b
m��:F �_�U1��<lH��.�,��D��'�Bn��W2�ꯆO�'H^Q�zl,��������5�7���8�wV�Q7G,��v 4ø�9�.��-�ƛ�-�D���Y���ɜRo|���U�}'~͛%I�I\q�s $�@s���&F4꒲�����D-��� �h(͡BP
\�X�`�)��|��1�3�Hm���n��ľ�Vڂ.����%�����Cf��������Z��-v��V]d���āj�R�[ #l$�o&ý��%�+ 5��c��p�w�;$�V�8��ya!����Q���B
P)�?�l�  B|p�ꆄ�H�RVR�;T���C	o���k�0%�����q�T��K��L\`�k��ew��&��?s��ɠω�v��j�����IA��Fz���ܓ��e�j��2w錱���-0��^Z��4p�[�6�7��M�#0)fיa~G=�����P�RYo��&�ƨ`���FP}��� ym`�7��4[nN�����K�|ex�ꬦzU)��|L�3��U�G������~�|cٕ�ۊO}�N���ї�ā����>��
�E{o�����:7 �q�e
bU-��N+=@U����tMM�i�eG�6z"��\�`�$���Z��Y ,���<����XY1��O��k.�Eyc�%��eQS����<"5f���lk����$��ƞ�`��B��W��}��L�ߕ���D5�	'�胜o	{�Y���kTq��ۏڷ2��axf"	�k_��IJ"/�����Plu&\���N�[�14^����r���v�ɡ�7g�v�&�o�ې\z"3��Xe����`����Q�:��P�y�|�y�f����ͱ�;	X\6�[7�̑���c�4w6E0����DӍ��\���f��Z:�I�~�bmE�!��3�B�(�XFdZg���~��Ү�r����6Kd��3	F��Ox�6c���]�1��^.W����x�b��WI�B�EGz�=9p�b�	U��5O�I�c2����	���7Cr�L���
��i�ީ�_)8b�ۢB�w�.ܤa&Z��{fr�_a��ت���(���Ƚ�s��Q����yo\$���rbB|g�-���$�^~�-�}��I�`��>��\d/�3�PIG�xShLCb>mE���vb�����`��*��2�3p-,&T�J�~[s��948���b;Hk��Z;�D�+��t��[9eB^�	qQ�B���p%UU��i��i+S�DgM����<T�v�tt���(x����`�T�D�����3#D�ͅU��K�c��y���~į�R�)u���<��ޱ�sH�Z$!|���?�iK���i/��cY3�������U]�g�A-*Ս-V����y�z���珋�ɾD�xDq�6Tj4�0�0a��t�P�����S�,~,�PE�H���z�ٸ�@�b�����#݃լ|6I�B���wİ�Q��$)Y(a���2w>ʹ��#Xl�����IA<�.'�>א`�V�a���N�Afr\��}�(vti9F�qIaB=��B���Z֠��y�5G�G�3��(Ss�4lh[wBG8���2��'�X��o��$�a����zZ��=,j 9M�"k�b,{���C��M���a�[D�(^5��ɜc.8ʹ�[��<�����J���c���}؏(�;m�`��W�w#�k_oٗ�'�F��yn��ݏ)w�pZ��
5�^���tY������W�)�x��s�y��tJ|�`��V�	�Lx�څ��m�
�wv:=k�BܾJ=X�QK��5�f�c]_@�d!j�Ֆ�[�h!j{>�N��\G���<U���4����R�{A]���>%�����v�%L1�~q��g�S}�ąWJ/���=�Xp�����]�*��²��]���w92%�M�g����>�
J~������7�$�M���H7�9~�b�eF1�4А/c��݊���t~�,/B�lm��K�~���Q�8�2�[�����O�=�?�Bp�X:���n*�z��3>e��rF�d|sF"M
�k<7�7a<�I�����4��*x4�unrm<�|Wn?����2�D$
=�޸�������v}~
v���h��J�)�w�G�C�r����@����J��&l���0��Z��I'*�9���/�Y ���È� 2�0��d�k�ު��yZꃃU��Z���BD��t�΂]MXwӒ��J�zv#`Lݹ����8�w\�Yj�"KY�s)���/8�
Ő���2I��o�l���5�UP�_��j-i�J~�2}��� �3օ�g�����G��:bC�`��Q��?��u7�?����t�x;����T+~���Ѵ&5%�O�A�#Vi?��V��N�ݵa�E8S�[=���aP(�|���͑��h���z��d�a��\f�u�夫���O����@L�g�s��h,<���GF7���(��%���+A���C�?F!\�+�hH���H��dnM�ܒ�ߕ���71�� ��Y�}�������$#!�e�)���N���I�K魽HH�w�S����t6�f�FJB"pz��_R]���,��w�hȁ�E�0�=����oZ��MBΜn���v%�<�_V鿋Xtڐ����s�Js�p�@C$� 6����S�lԢ>�
�\3	������Xq9_C��Г{IS�i)���^��6�I�to�שE�H����C�]&O�%�����>�V����)�^��;����R�},�Ԧ��c�-Q����T>��<7�ق�Q��RJ~�%*�%V����}�@0�hVr��pT�P9&���O��]w����99nS�^�KPeQ�b<]���R!Y���%l}=p��u�1�.�h,�s3�0�y�B�xnSe��G�-qJ"��[�픽"�SU5��mM �r9%9�(\W����p��ɘ��`�Һ=�c]Z��P���7I8�(�CqSKy4t?�ؼ������#p'�ŜF*�0h[B�"���'W���Gډ�@P�����c��B{��V���0�� Iv'�"t����"�>��s�!�'o�G.;NH�IV���l�&����[m8����u'�'Ps��#iO�A��TF�[�_���{��	ʗ�Zҥ�ܸA܋�X�����������Cr��Z\G?%9t�>fg�겙���G?F{tq�NW�z;�=����9��Ӑ�
iM�9�3�&���X_DKս��"�p�ͩ�;��э��$v��+p� ���>��ɾ��=�1�V�e�.
}q2L���k���,"6A�`昦�:G�g��?8�irٝ0x$	�d��y�k6���/
�A�2��{�t.�st-gCa���n��8���-���wd��>�iS1�o�1�ˮ����AJz�V�4I�N�ƅ��y�%=�nHw��e���/�`��F�P�UB��)R� ���KaVj����*������yi�ʾ���+}�TH���-�^��.����5���r�/�R(6ʲ�L
��W;4iȞ�*��*�\6�lg�܏�h�>ؕ�=��˭�d�[�xT�\꒸rYtJ
ZG�V���2%\�q&�ɔZ ���;�}�t�g�|��[�M��B�}̓���-���w�������O2��S���c ��}�Ɲǥ�^8N���/���q��L��`��6Cց"r&J!�"^H�R�����&B�}�%�V@!�릨��S��|�.!�g1��j���-�Oǒ��r٭ tްRDn�v�K���K!%o��h,~s�Ƚ!�Q�s����Ee��L��p�$uu�Ï��Oh���L0�&G�q:��,��%I�$��9�n�K�I}�:�)��zx�m��(eՄ_[g����m�Nf�eǈ*��	h��<S��K�1I9q��6�f�bl:ׯH v�V���0�Rn��9�C�� ���s�n�kO������{�2i)?QPt�T�E�P��"mK09Xq�-�_-VMB;���8V0='U2G�c�x������{o�bS�jMo :4�`֘.���(˼���(��&���tO��%���#�Y�;1jPߟ1��dT�<�KUt_>=P��q�����nt|�8�	�ؠ���(�F��E<225+/s���W��:E���_祄�L!8�����%�/�1m������D>�K�"�L�Ƕ�ᱶRBy��]��̲-�P�#���U�0ӂ��6Ң�K�ą�����B�~`@Փ��Ug	|՟L$|�,Q�%Ѹ��#k�:Uf� xߞ
2���p�ׯ�WZ�>h�Y���²Y0h'ҿ��E��Vd{0ۣ���O�����Kr
A�!r���<�t��K�S�H�g�[�����־���	���.� xT#��fC~�(��v�P~��������5�O��U go{d"�оK���������H��a���/;E@���
����Y����d/t��{�t&�x������ ڧ���r+���-u�d��7z`�}�ԨI@��.5K�J�I��C=ʔ��s�
���m2��k]�C˷h��t8\t�xTeu�ܓ2��<<�x5P�E#C����DY�DI�-���1�f��I;��9gB�3�m���*�5G���U�_C����v'��2^J��#_�	C�;���^X{W���"и�I�c~8�g�4얅 ��6a߅�)�f�!��2V���5�Z��a��G�%v��tqZ��p�.��(@�����O�P�f��� ��O�q.�/��ԗ����v#�C�"G)�Q��@o�Җ��p� %&!���%|;U�fH����8n�1q-�9��}b��m��[k�� �|�L_�)��<#����e���烸p��r����������p: [&�Ӕ-r�-2bBw�%!K�S��� �G+p���;\��(�l��W��	*���_#�@ɮ�Bz�/;gFX#�ƸѶ$E�'�|���|�^F�0y]b����J(�$}˜&��M��֌=$�p�	��akW�}.��Mn��DL�`D�㉳D��q?���{�p���u3m�JA��

�C�-c�)��pE���{�cx� �����QQ�:��s��pQ�M]����>�R4�q���g�^ݟ�la��,\VJ��w_�Z 2`sA��@��Q �*��U�{�1y��67�_�/��y��;�xWKX����e�1x�~RG<���]�,���k¶j����^��a	%�yk�;>�u��Ւ�u�5J8��t��t���-�V	��0�o)�b��}��q��*���o�rz@��?�mg~=0z�WԙKZ�E���7���b�����s>�p����HEE�Ȯ���d#�,ZA���ǖ�Ay��䳙1W2H�6Iy���La��v	��f��fq�O�Ec -�v��; 7S�c>}S
�y�c�ː��;�(�0g��l\�7H��=2���q.�<-�'/���V~����%��8~2���=B��_^]�t�Y��~0����B��{�+�q2&��YS��&?	l����o�}ʌ�R��%�U5�p�J�H���ٶ�/��Tt�$бl��i�EQ
ry"@����!�AA�����gK��FJB����5�D�1�K�sB\x�HJ�2'.��h%�Dp�Q�v.qA<i��i��YBY�l��q)��^#l��� ���
o��^���'����a䗥3�3k��*^�$�Gi%��U5��77u8F=�>1R�=$��E����J������<hw|lJX{�NK7m�i�u�E:�e�	�Y�Z}�n+OΏ��y����i� p�������ח��{�H����*w'�ֶ���̇w@�4�ͪ�Dh�86偙yp�8n���8���"܌���`ܫyE�3O��^�D��*�)!�y� h]ӿp''��=���<t��n������Tܗ1��g�Z�i�#YvK@�[�V���%����K�t���	���',H��X^�n�&ʮv�,�1V��K��$���ׂ�̰HC�|�),�i։�Lm����hd}G$�2z	���NN9_k��~��u����{������8a��/޶��� �G����V8xn����$���6K��DyZ�ܿ�Y�����n����֫�r>z&����w���a������	ad]�q��kT�Π,��q��d>'���^�4q&WF�2<ao���Gs���fQwiB���ܴ�B�*��ۺ�u�-Y��Z��ɩ���[���'E����YP8�
�@>>P.�Z8�km�Z!�t+����J-��r�zr���,r�#��B�jg�`
՟1$�H�9UC\44H��/��U��l�a"�.s_jd.�W�IBg���Mc!����e���R�d�X��V�1��uR��(���a�fδ�x�-��	����r��OTŉE������0?:�Nv&�='k����G�f훯8�� e^!C�� ��,FyL���x�;��s	r�@�$?�5ea&g_|��X�[u�߫m�Iċ]nfjq����]�n&ţI�Bf:DNNt��:�\������~�מF�-�6l<���z�,�.�Y  DB;^�z"��+�Mۿ�#o��5Y��5.K{ ��,�̉�hbn���4_.�4�H�M�\�F�)]G�+�߄��z��*'�IY��ۗ$G8P0�c�b	=��	�ks���u:F֠���4�2Q�G4)#�\�f���;��!l�(�E�8YQ�ȃ��i���-$��r�h+Ȭ	IA�O�����c�y��U�vr��	G�7퍦ڷ$?o���L��E��<9�
�\9Z�b;Esa��D��_\R�����2�ltJ�Oj� k1��W+�v�8�Q��<�v$y��BR�i<Lv�b��
��Pr���.3q�Ե�5E�Yh�����you��o��]��}4J�t�,y��?��������4T�$c���,�Eox0%�Qv�nU�5�!�x3��Ճ������U�l��<��l!�JS�6f�F"7� �ܘj�{���#q���#���6|�Xq<;rջ.d�,��	g�/�@��OSy�t{���A5�?��21����d���v��	�-w=�Kf�A�}<�D��M�*����g�u�_��H��)�(_���SS�Ĉָ�eЏ*��j֕�'�;�q-8!��!�o������j;f ����������[S�2�3M��k�T��p[�K��&�[��T6����4���2��� i,�ae�>̫�1�]� �iTY��a(O�_\�Pr*hյ��T�z�ҔgX"�"��P�}��8���N��:)���cnˑ~r[V�*o$��*+F�N4|P��+��Уݞ��Ɇ��ǵQ���c��9sO9�¹P���`@ZT�
��������`LKG|Y2�0P�o�ʧ���Ml阩 ܈2i$[�4�lO�o�����g�d<g�w�w��RX�Ї�q*uXo��HS#��sn��D"�h�x[����ҧ��DvBᘻ�OV��M2ҷ ��&� �'�c	�{�Q���#�BQ�D��B�����]�s�$b��do�i.��1�x�3l��}�/�	y!����0�"vg�
3#�&'^�\��aiۓ4�,B��2�x����jA�:i�^�^�.���Hq"�>�sF�-BC�N�p
��9{�Ty�1�(�������>Q/q��oS��U%�c�-��^�V��7rs��������(�Z�����I���A�16���j��$
02.���@�q%�tp_c�����`���=@�&� �,�i���`�S#2�0w���<4]QI#��'��
s� �'k��	��%��M��Yt��
^���T��I���݂%������:�)����vu���z��Z����In@�(�"���ڑ��$L�'�_^!�W��6���0����=�(��U�1PL1��+Ju�6�,�6�Nh�>�8/���1��/5�+�nZ��r�Bs�f���U1\k���'�Ffǁy'�	Pmveߏi�0�R�r�b�@3����sj��L��Jgwj*;|���j��� 6�e��ș�ծ7�hID�q[۪f���.m�� ��$�W�c���~��NXE�x�i�vf|S�N�/�� 嗟���ɻcJ����4�.9F|����-?����<�� 5;>���+ J�����|�m��gZ��"X�g֗��� �KŖ�yh��~2P7?qX�*f����"G\Й�0.p6 �z�?	���k�G�v')N�h�������݁-TT@���_���}Q���R�9���n4��ʻ���f�P��{���;�}e���f]���S���N�G�]8�X������^��9S�#���-������h���C�o<�_Q�9L�͡���/�wG�����1c�("�_�d09��p'a
��[o�y�����$��~��6�@~�c%6"����Åf���}����ƀ3e1��S��p��#��b��wwCDtց
��~���Pd�ذƊ��j���
�����h#��p(�����z�h�(Ķ�k)��_���I�F{P�8�sne3��'����s^�kޙbXv����rYi�,��rgI�x���%��#X-��D>�%v��Y�,�[;B�ꐉ��`F-~��ߞ-j g5IK�.�� �U�;aM/~��-��-�:P�g��pp����㋷�H#1|��s��.�p�زK2�:%a����^���oQ������RU��yV�p��q�~-���[7����ʷ������J$>kq)�:Q�K��р6��T�z��Zq���{�c.	�;�7�Ѐ��֟�D��8?������h~��^������7�)��4��'��9W,�7�
7R��L��L��5����)8���*��i�`�_S/�p�<$I=}cB��u [L���%�J�n;�"��������BG�������DW�.�d�0�~5K��������3v����Z�~;��Mh�q�>�ͬ�O/�G�^����{���Ms�Jr������Vkk~��Խ&�"P�{�����
�NY-�̴3��I�q��u�~�N�m�Y,JU�IDyU��yx��c`H
�di�B�9W�z�XfƭQ$��I�V֦� �Y���5�\�g[��]4�"�j����@���G��V��ϴҍ��8.v%�BK�󔁹O�U7�A���OKݩ���R�o�q�|@�d�V���0,T�����T1(�t����Z���Kf���1�Ǥx�I��(?½���c4�N��w7��P��(�Ծsz]_b_�6̫����l Dy�67m���"2C�a6a�L��.o��'���oh�Ռ#����
��*��6E�R�aP��b���j0���نq�ob�IT�a3�<��7�/�t��Q��;�bRg��b��Au�~fT=Z�J�=T�1\y`�d�:F+$����kVӺϫ�3%��}hx���t����f+ˬ�&u���ͩ��\�{��|�k��{�8f�������z����R��H�D>�J宮�哶��Y�,^��W�>�G+����4���*�Y������l������&P��t6�`@���L�4�D�5�x�U
Þ����/��P�#3�q���[>�� ���e~Ra=���@.^;�J��`E)�>���\L���;���>_U����n��oBA���W@u*{��D-��Q�˴��慘�_	�By)5��X=L��[�wF�3h-m0��9 9�[��&��'��C�kWq�#� }i}��4U� `���W-�(�7��\5�$u*'Y�7��&�q<�_�;e��.�j=OD���-r��F���I(��}u�{(��騀OВ�Ĵ�Ō��Ԇ��d's�Z�mj�`"�X̋|�:���.���(k��@�

X�U����
�1�����v[i�=�7�}����;]�Cu��,7L�*l�D��r�-�/J	����������rn�3�,�����`1XV|��`L�k�u�*F������<�}�բG;V�-��ۤ-��R��������|ќyDk����]3�w��enP���S"6��n��'��ǯٶ+�a�Hĩ���@ y9�xp� �E�E���E�j�I":7j�\�K'+�X�YB[�o�1�l��PйL���T 3�V�{p��R���tj�������+9 l Vgo���0��u��0��C�^v�0a�6��T��k{��=��)�S�> ً�&$��/G륷��tW9�K�h:����,-0B^$��(����
8O��-��M�96w���>�A$<|��B_�i�K!$8�m_�1��P2�
�J�$21��k�O�Jړ%W߸���h�רi���qF����1�M�] ���9b> N���R{¯�����	������`�92ז�4�����[��dM���@���o��oq��}�w,[F�^�j��L�#ě�L|ޖ��µ����9S�N����8˦����u�33ЇHH?5�Ԁ���̘ģ����*�!��J>�	���W�@��n�f5R�z����P��6~��
$�*ʲ�®GXI�y�mF�
xE������m�8o�.鸱��٤m��"gH��n���%�/��T݋e�%�������*�k�/��W��]�!��h��R��XU�E0�-��s��j>�?�K���"::�V�p��ђ�7�!!U�Q��S�H�+C۠ C/��P�i��� E�+>!�S�p���
�i'��p��䜾߃ZW���>��o�ph	��e����a)7��G��q�3ڂ��m�����R�΂#8��bo�e+b�Rip��X��~��Ql+�G���y�&Z�pR06�^-<#a�'Z���Z�Tq�#�Sx�Oq��r��Sq�x|�D�i(�gݳ�b�y�h�K��)�}�o�/lx�y�m`��t|ǣ2���i�F@k`��@�I�Y�+�"�5�i}�dΗ
��A͑<W��eŉEX�h��B!�
�#Z�ޯo����[p��7{����X9�R�+��>�u��E����4&r�E�%�t�e����*�8!5�%#'��^��t:��Y��C�$y�C
��hP�����{���*ZZ;�A�hS���g�Ѧ�uG.�yl/��w�E�(��2y.ׯԫ�>���tlKl~��h3���i����[d؅�		��w�����4k���NA��q�$3J�>j��r�*1�+��q`�-��f�A����*��l.��4fEl=LPg#ns/Q�Ja�.^� )��+g|xb��M���ܼ�����5K�yr��ǰ�Ej�ͺ5�Dei����_q1[�s��fnˡW,;�VK*���g��T�r=�ӘO���yL��<#��UB�-B�)D�8���K���ϴ� �)�E����⇴�v�:<QL�+�>�.�p�6B�·k�8@���7�r�M�s��X)ե'Q �#Vt*� g����q
���qڈ>�-9rN�o����A�_�\�qP�/�ͣ+��g�`n�@O~�r�31G'�9PM8�AkU�V`0#��z ����dM�`���mƫG�b�!fM�X��T"XR�=DXɦ�H(���|
/s,  ��,譡ZB�Nn����	� ��e���QF�SV�[ NŽ�\��� �.oE���_ɻ�Nؚ�v��"��|�^N�ɪ���d|��X�DWc����W�{hظ��^jI��i��\Ы��Ps�!`{�d�G�yG��:����mŇ��;	o����ÿ�c�D�'�7wO��'�+�1K��U�;���+�O	C�����㴘�����K��'��h%	�	R���GS0i��&��_�c*˗� ��I��P2���|�,�H�mk�3�W֋PO��e��\�#͌f׎[�F���R�<������+��Aވ#���l�@�HphoM�{�-SF|��0����:�H��~4���`	�AAE����)i����,M��2m��y��x���X��)�s� �{������ŝ(8�<pW�L�(Q05r �� �^��(7ތ4_�.�Wg���[1�m����G�!�u@�[��]v��LSBfTY��T�Ű���;d��/\sI�jѕ���	'}��a����1��#,�/�t�h}m=$mUskw��K��4��|�x�k�@�ڑ�%5+ƕ��6�X��\��W��V��^q�E��⾟�4�F��^v������{�2�������A����R���ճ�eu(Y���܊�c�}HW���wϣ�h�ݬ���kC�pIF��5 
��e�/�����}t�S�0)���*�)-�[�r3E�"�W<��{t"�������.�Ə�퇫W�F"�8�����_Y��-9�@��Ma-���L�׷�m�
`�g���pA��]vD�S]�HAԺ�m�Vl�~�q��MN��Y�X[B�',:�.A���2�pV��=�D�u���UQ&�@�}��=N0g�Fx.��y �Hn��ŝnol\���o�E+}�ae����� �q�gqU�U�W]��sD'q[��ZW��es�:<�h�o�ԉ�S��5wɒ!Ƒר�ʂ�ױ_.��7+=t�xk�v���AG���y5s��u�frm��XG�\���ӒD��:@�ih����Q�l/��YI�D��,˒�؝'�/�������{ 6��ق���^��Ee�!IX2.Lj!8�'Bff03��&P�S�����>Q�3�jI�jbm�e�7td}�����A��V{��߄̯_�B??㎍�30�f%���>�TO��&u�?h����Ħ��� ��A$�!���0�Z�;Y�� 6	O��nZ	1��(�Z ex�,Ć�׭�����ϩ1ݼ���^p���g�0���;�ᨕ��֏ꐨ�(ji�h�T
$q��fl7�zV^�n1�h���Z�>��2��w��p(м�+8���n��y����E݁s�g�v�@=Ӫ�`]:��`�>�Y��A5.����\f		9����'���Q
�a��Я���b9?i��/��k��#��/��ɯ#D����5������U�͝i����)z3�_��6��NKe�p:�)b�ϦG]�g��0� ��
K�b���}�A���;�܊�(FrU�r6{f�`��zu87No�e��(�=4�fOj�(~�~&#�wc�NQ���I��oPTT��?�ܟ���{�2��Tҧ�y����l�΢�dA�9�x�n����U�cdc��gޞ�|�6$EY��m�͵@.]�bU=�~T��ӝù�@�2�.Q��D��7��Y�����Q���}�U�y�#����䪝���ĵF���� L+8�Hz���/�"K��Q�)	����p��+�&D�n��s��������nU�V#�����+NW&��'1!7��"C��ܓ�H��6b�=(b��Ν&Q��q�����T��^�W�`M�w��[�S��?[�pE�A���9W�	��Kڸ,��ޝ�'�+�c\�Zjq5�x��L��3:�t���4��x�(���:�o���U�^g�T$Y`���ы����hץ]ݘ��
�`-Qb�>_,�Ri'!!�D�'�v�V���]S@���^��Bj_��N#��m���B_i��:����u��U��6�-�$f�Ͳ���S��P����}d̅&,$�����h} V������dgҡ�=���F`j�n�B���0�d�4NP�¦*����V�@V2���XJ8I�,��Pŷ���w(?�r��t}���S�~�dӦ�[�v=�y��(&��H�ʉy�Ȓ'z��Z��A�:0@��4җ#=��n����(��\H_�f��Px��rf�{7�
��.���5��?��2��,9�\����`밷LD���� �?.��diݵ�Z�eW�#2/(�G
�?���*gd���Q��uC���g�bN�U��?D�ﰯ�臢-׵���-�3ܔQN�ީ��%&u������-���	;zM�QSu�	ɥB��`)츉�z����w%�����<ǩС�H��z��e[�n��~��a�uaho_3[I$��2�b����b��Dٿ�8��<�V��e.�=p�Ҕ�]���gܴ�"�zζ	��?�K��{�-�v�N����0�NQ�ܺ��Bw�1�4�O��/�t�-b�V��HWr�:t;U���'���5�?�K ���O�Gݭ�H}Ο[{1�P�:�|_�5�O��م�׳�sW�+|�Q�s�Y��Z�1e��'܉EF0��teyA�mkȔ���8�Nާ!ߦ�eFb�~1Ղ�[7"�-]	�d��J�lbd�����%�aj��d�R�����Fi�[��O.fZ�Ra�׹)x� ��k�>]�KK�#�!
ǚ�/��x��)�Q�:�k\;㝇�4_�%��=�������Rɷ��zl��0IW�	�vR��,��TMP<��/��9{�:��0��J-���L�I<t4�7���H�v�F[��*�H�1U���Ζ7ׄ,��'��TW�����
�����vL�ѱ�����1�57'º�:��.IH����)�^X� #���g�t77�8��d����)51��.��Ϊ�,�+]���jiɷ�*eNA@����!��ÿ��jk"��~"F��8��ң�!�ϻ6��C���+�:
󲏨��sqo�����Ut����#!�C5@���s�9Jo��Hd&`���ɦ�¥	�AqA�X���1�-�d��p��bC?��w줥�k̼�\ �{(��xX� �+{���-L�L�L�T�)�W}����k��e$/�� LY����S*7i`�9�����y;�೏����z��u��8a]��k<�~8���?@��g��Aٟ`���3]v%�p�`������2��;�i�o{���e�Cq�޷�(��^&�?�D��(�s���3���]�b��"�g/����'S'��??��66H��m�_/��n'w]:�g�s��k^R����}��o}��h�U�K�c���0v�Wd�i�X�]u+<�� ���)�ݙ��B��hh�%���s��m�;XӍ��q&r[��)����x�FF�{��i-y1�X�%I����� �4����ACG־^P�]�|^�а. ��i'3�E�޽�{�F�}(��W�Gt��x isOl���`׈\�O��?���G����ߊ��tϼ�N�Q��܃�6�r��M�sH'������ٱ�� ��dQ�86X�Z槓��&,�&y��x8Z���o��ū�9kl���]��{«�hN�¾��v�Q�^��w���HƖ��-d[b2�!��=�w�w�6�i��ݞs;��M�D�3I��@x0��z�d:P��M>�ga�w}oj-�dX<(�Ow���}���(��>p��!�U��4���dB^�ly-cD(�] �"Ǚ����DBZƑ\�Uʽ��Q�n�ar���h����'$�O ����~E�\rq��1�?�
����Ţ��Sj�K��6 ���q��r:��@_�C����t�ԼBJ���q����cP[[�	�Bq����~P=H�^��oQ����4�"����/���;���b�U�j���a@O�zu�]�>>а	V=�������c��Y��US�#ܤ���W>5�|-���{�3<�]Js�y#Y�q���^���iI���c�/�a�Ӫ5�!EH4�f��ߠ����=��W��^� |��͍��߻tV13J�hi����I�{x� d�w8�>3����僓�r���xܠ�k���4�h�pS/
/J4�{���}�	%Ws�Ѫ�G�I:R΃��s����6��4|�cX��;-&�h�zA�+���'{&�y��-�; .�'v"�5W%C�_z8*Y���0�Qհ����*��ih�d�
�$�py��Ď��ʗt4���5�4}ɒ��J
C��r��&��.A����&�����,��^�\��P�����I���I���!�w�ly�d�g67��;����S�A�c�G�]̽5�|P�h����32yF�_��}(�4�*��TO�5�ٻ��f3��h����}�#w���p����tZ�*���/��<�������:����$~b�n�`�9v��,���1О�%[̷6GJ%�G҆�����/b�TZuJӈq	l����yg����Q��(���3�DkndimO�W��)��u�h),I�Yu��čp�������db��v.-CKUhA|+�tFM����]�
(r��g��=����21q*��`���hx[V\��n󹈴�� ����m���jT�^����l��Z8�6��e�%�����b?G� ����|�AiR�V%����x@�(��-��iM �Ԣ�x��1�"��X���ko����6)��[0.h�
yܵ�sLr�<7�*_�Z�~�}�������GI��	�@ F��b�2P�b�׮��ai�X(�/����pC7Fw��cq�A��[A~Vd��N�ڰ�8��	=�5�dt7PJrc|��a+z.��� ��'[mB����taI(�~w�8��4��g9�aA^�����9�x�I0��SA��*B�@z�xPۼ>�"�Âp0#!�3�� �t=QKL�К�(?O}���EW���Ϭ\X����]�f������'�
(�9��]��m[�꘼n���Fh?þ�}��+��R�^ÚvR��qg��4t��<��R�ma��&���%��65H={	y�F֬\I[�$e��A/�5lM��y'k��DH0n�j�d�Dx�I�t��NG�vA�'��6��h�?u��Ćc�3�nF���q"K�wb�Xk ���J/��m8=%�ȧ�be2�fX����j��	 ��Mv��"�c�?�\?�0��n����*��O�^Њ`�w�;+@�4^��p�_գ�&	�lCkߙn���w��L�V�c>�5���ً��w.ș?f7شb�%�%&��~�δ���*�S��5Ib�D�" �.ȥaIg��b�)*_��P������邎�Y���O��B.o�*�Mg��%5q)��3n��$<fK�b���Q���r�P�zՆ�X�����Uu��c�<k�j�l�r0���S�GHH�}�^�fm�h���Lݩ��:dll<z�$��9 v������ns�k�-��ap����XZE(~��*�X��cj��?��z�E�����1E�_�$��Ϟ�P�g)�`��^J��L��V3ۧ�p|l���>��,�l=�'-�:Ћ�N��u��5��'�@;�+��1C��A^Y��{=1Q���a���I*���p�,FA<��W،��v*:���
�4�&���EzE2�����F%� �U�I�w��G>�C�6T~Gq��K���`<!��jU�kEƠ�@R�2�=v��!��dM�^����1�����\��k҃�Ӊ��@����k4G�ƽ����ق~Lg�}���]�ɻ��|P]���%��V �����a:
�qM����s���'��$�$�]��P������*磨:��b(镱a�E?]�Q�Bq�b�Yn�~��kE�|�8���7>��ґ����~���VrH�=/�~�(�w�Ll�ݏ�ML����صҮk7=���7k\�6�2Ǵ��K>bjR����U��ÀI��SH�dPb�3�z�kc�2�x���u��ł�$�F8S�zX�����v�֧kCn�����w/2gF+�T8a(ǒg�H!���ELq�=o-�,�9�1�j:'�k��"����V�o�PMV~��K2�*���o����)�3��[O��X'\G���0?������5��%�;l�-4�
E�@�������=����U{VH�YC~�T-�|�:݁��R��we��N'��m�(�}��e�DV5]�=���u��C�C< 8�-��k�UaNm>I��T�W�%��v1n�ԃߓ
^z�ޝ�
x:��z4��܊3��c����f� Kh6�Ziز\�}�s��8aO��|n.UK���9��?�1o�' ��N�d��iԇ��YC��[�;k/8}Bb�{ E;�*Q{Aț�@*�/�u�w����\�W�_dԲ�p�Sbޤ���gO*��5*	�s�B��	?��[��\���	��:L�z��;�3����%[](�L��_��E� ��n��<�(��9n�>�!�\��8)EmK
(Ya�;3�a(��
���Q$�Rg�љ'0�y��:0���+Td�X��AQܽ�<z�Ȃ�a
VK��u���[�G4�*�
s��1�/;k.A���S������1�AI�M7 Ƣum�.�X�U��	�V:- ��yc{3v��\����5�DK�����jhΫ��Z�I��L�l5M�P�f 0FEj����qx�q�|��s*H,&�:d�
��0?�Mdl�-��@'1��U=��upt�H�� �o��qq�oE_$>g�'��7t8)��y�j�97��-�n����@_��I��`U�)���{ӽ�4A�����Y�v����/��1�j`����:�%�u���o�O\ +�\�y2N%h&��Y�R��\ޒ���n'Y��/~�POw�p���N�[�1��)���ȹ}#W|~{�ص�w��Z��;�i&��(Q3��[���'�d��D���-O,=��Y�s��0<`@ڮDDa�ruSB?w��D��X[����w9�ʠDFD�;o�� /�s	�i:27B����:�"��^�ľ�KyK��E�-���n�V�>�g����l�$9<F�譝V��"qu��E�q��Ϥ[r8�L,Ur�)���a�3���Q����Kڮ� �����o^���:��Ըǁ��S�ǽ�5?o��P��k�hD{,_���K����BT�0í��2L��}�Ǭ�t�
�����!��q���]�?\��J�Uy��|�-�f���:�O�L��e��
��ή��Q3�t�_2�6�!�9<#�� ��e��e/5�W��[����IڢM/Q�3�i�cA*͋�ѫK�����?�l���u���*2q��h�>Z�r���0f�H�����b��7Nk8�p�����;!d��������ȯ�zi�7�܋�-��E\�u��!���'�]fa��s*�[��k�b��a���V$�b(h|�8�:�P����	5�;�Q_y����AI���&����#�LT	nT�ةD�}��B�a5�s�,�U$�u3*�ṳy2�
�K��#�QXM�8�����R��"2*�(W���ć]�iN�M3��:�^���X�+s/��Q+��;��S'�u� L�i���Q�K�$C �S���w���U~�\�'B��)K �T�^w�DI�Qq�5ش�����1���!�m��I����>�{��i��'S#������w�c<�&�[�-.f�-��vE�CIvfv���!=���6�B�19ʩ�)D�Ai0a�vjM�N����n�s_|��-
5I������R�s���]r]c�O��"f��'�������T޺~��*���gY�d�u�V�����$�������+��\��Nh6Q�8��'շ0��Y�J��,��xC��[H�	�1��
��5%p$�=v�E|Sq����� 
�����Z:���<}�>����!������c+˽��'��QI�����q�ΐ���k[aႧ���1����M/dDx�V�� %z�4�]��#8F�#��m��� �6�(�������WG����t+��h��vo�����e��R�z�
?9�-+��\���[Wΐ�J
1]��u�0�Ƚ>Y�����R�Zj
����-�a�s[�-0	�EPz��������Zo�2��u�4D/�J��Z0��n��k�����;��"��1KW���W�W׮Er3t�t�^P;��Ղq4�u|��g�B
K9ա����+қ{����pߨ�qi�y�`H�1�<u�T�����{C0,��+���(��Fe5R�}���9ʌ�F�ґ��Ok/
�/h,o��D߂\U��m#c��;��27���)U� ����D�����B'?�1������s��ܑ����8o1q��<�:��Z~�ƮZ	Tv�9��S2+?�1�S��cw��[{4k�=��|N�5@Z�P��o�J?��T�b����Зa�U���.lt��^�O����/<��Tk�u�J��Q������������b)H`)��Y�~�����	'���P��jw�4	�Qm#��`��+���5��WR}��jpI}�`��$D�4i���C��jX���@���L�>��+��qtQ�[�d��я˜(��sl.Rɸ&��!�>q>��A"Z��~�-E�^��4�(ϗ�	n\�w�77З�ۥ��R��f�����_WZ"�O
��?�k���p��y�~0q�Z.�����!p/��62L*��$�o�k
��l_�|o3�٪�mU�0c��۫@��9P�;qN84��>Չ�zNξV��F�����Q�L%sU�����M(����j�(�=�L�f��k��p�_�n���1M�d#J�t�uØR^r�9����7��j~+��F�����=^/+J�a�V=�V]%� _����EI�|T���E�A5;���/`Fܖ�l�ꬋM2� �����p��z����������g���REv�8����T�
�.�'��cq]�m=.K7}L[9�H��R�0l����:��Ķ�~+��\�ܾR�4��*>�捠/�{����N�X�5 ?@�<����>/5Y a��x�]J�������p�X�6��FM�i�YWxw)3c���u&���
�Fe�%ҡB! C��˽�M�`
��^��� s���\���%��S'�nV�>��I��iū��Vo�t6��(�c2����:�P���\1�d�!�HGB��vh�D���.�s|�k����m��s�v[00^��#7i��������6<�������EFpW���HFuwB����DIWu w��m�M��@�ŕ:��CY�9nW�
��G�^Ե�+��plכ��~]T�@I���:�w]�f$�J1�%8vv S�3�Ifx_�n+�V���e8�7�%=�}@�;����Fe��4]:)�{<�L�(�%���3Yėvg��ܥ��b-�jw�xO��e��Y�����pao��8K���.`7��y���}�?x-�A���6p��T9�@;��aި�W�����<G�Q[_�JA��I��U����1��W[��YI�EQ��!O�g(XJ[��ħ.�����E�@��[�Y-��9Y�n�����e.7_>��]�@���LJϰ&�Fp��lz�ޓ��G�Y�y͋��iX\c�F�Y�hsϿO��lRؔ4G��)��#m�=�[�
xG=�@O�)����$��������ğx��?S��-b�l}�O��];>��V�ۘz[�q��3	fb]L6g���/�,L��q�P���Ȳ�ytnb'WP�Ǻ�ĔB˕�M�۳$�œ�� �s0	٬��AE�bNvF6J�H�;��7�˿���p�l��fH0�
��L��q�+0Z�$ҬCS'f���t;e��
~XS�/�i&�hn��= m�-�5��j�8�w$m�����p��s�N�Np-�f���1�4�os��ީ2.7���Fq��\���+��u�K]6��)�P"�btWS$޳V�ByrxԩHVN/(�DT-�͵����r�;�/�o�j�;-,U#܇3�c�2���N�"J@Z��,H���W�(��#knU�J�.CIW�"+�����Dw@�T~B���T=J�ֆ�d� 9�8���pq�a|0��j͓�А�$`?I^��˯���Ǚ&�����o�Q��\b	��QP�b��u��nl�)'
m]懮f��_w�oߟ���"�D3Ye��h a@�E⊎|I���5�1��#�g]�s��ᛅ-�vN$���������G���s�H���L��e�M��;���yT	?�eo���-�bU�2N����J߇$�_1�J�}���HEP$/n���w�@&��M�I���.��(����u�|��*9�u �̂@�$Y�(�6�y�ο�Szc��p��ȋ�LaS��O�D�.s��qr�ig�A[a������C]|�ֽ����͋�d���Ƕ�N$o�ͬ`DW���ݵ <�1�H�<�Du��ύ�����Y������1kheu�4��2�������i�x �����YHC}���mB��R�|>�}[��������HS>� ��hbOQ/��pN=���Z�Iڜ?>��
-����lƺ_�>]b����T�� +�A�T��(F�	-���C���WH�z�Ϣ7�48Dy
��V,n�J�\�gv����nE}A�6�[�glL_�>��˱���C/-�/d{�Û+�A7D=h��A鸾·s�{v8\(
 ���"�׼Y���(�r.�i�}�[�q�C�N2/	�y�q���m�g�����0�J_����o��y��q���Q�(CK��&H�m�U��^冮��x��V�4m��#���H݋*k��5�a�}�F�0rǨB��,PY�ڿ㧪#�8 ��$]�Vν�V�=�L�!Vn�#��w��Ur����g��N˗;v������ǌ��R0�m�M��T���m�0���bw�98�y� ��-:�N�L�;c���;1�el�cH��rA�ipwPB�͓&��_���m��	^B3g�*��m}�R�Y������a�kuیL���~4�`�e�d��ʖ�#�U@�[7�d=���Z_8�xd�[�#.���>P���ak"sM*�����Ζ��ɴ�ԡ>��-|���aM�;�|�\����g|�<EoN��
�3�@�c	ʳ�e����Q&�X�m4 �Yx7R'�|� �<c\g��d��G��r`&x;o��3gq�A�&���t����P��$�ɑ3:�grj#vA��
1W����j�뫊�d�CfV��'[���6uć��=�Y�1?פ�`��;
A���$�w�i��[ǋO���t�!����l�j�K�}�tb߆��*��H��_�S� Ro�1�X��D��)��Öp��$�J]�m������Qj�
`A*:S�M1�na�-dThE�� M�zo�oغА����_|k�&�2�-֬f8�̢��,2�h"T�,����GV]�;�ʧ���~�U��c����b��P<
ŚC��L	���p.��7PZ��Lyղ������,ֵ01$2_��Xu�8�������k��e8܁�%�D��T%1�xH�lᇢ�Šlp6F��"=I'����@�gë�[)��"ٹzvK���WX����lZ� ��XYS�0��a�I��eH�xޤ�+�U[W)W��Lu��m����L��9
t	�}C�[y��5���'��i�+�D7�z�F���c�-���>�bhA��=�g|ǧ(0t���H��
��|p�Y�	��q����w��I��?A+�?�+����c��l��}���Ȱ�\m�M���O7"��}P:��9���H|������&�r%%9���۸i��J�rJ5��H�ѝ�S�I�Qf�G�	4����tX������E�N��D���zWn��'��X�]�����j�dَ��^�Ǣ�����G7$^�h>��x[ԁl<�D��.��s�����(�*��,]9f#߾~! ��������[���^�8[䭄�X�"[��<��XC���GgR�m�i)��)���J��x.�ŭ"z��7���h�⎆.(AR���y�^�\�e^�[Q����mW����D9�K�Y{zp��{%l�.lf�FM�rJQ�pA�I�����5~��/�.�@�d'.�+�����D���q1��Zx!9��ƫYľRF6���;��h6:�B�ғ1k9�-T�CQ��5~<��o�k���X��	b��Ig�af�Z��c�{�}��Dj�->��v�hwC*e$ 1G�M�H��"ա�{���R`�D���2E�^BVae}����7�t�$�#TVo���Kw ��؟͹���NU#��Q�5ˎ%�	��F�b\'�%8�F�ѭ��5)���	����m�`JL1����F\V�x/��X���=�B��	��5��d� �rt�[�V/b�e�#��4[�Z]h���q.�J��������8[�s���Wp��LU �Vx5O�a"���7�VU6�E����"�>��<�"����X��R�'?�n���#I��D����C�^�l�G�I��<�j�oYg+Z�A�Z��*�^_�xv��yQ`�5\�u�g�J���CE+��Rxv�9��lM'ƶ=n�I`P��^SSF$i����+��L|�����ѴIݤ��z"?����Of�[�Z��!�^�o뎵��SaƖ���<�\�.{'�gK�G�=�C@%:�>�2 ���7�r
W�|���-��ަ8\-�ٰQ��A	+亙���E=Z���\�E��R]�M�&*��QxA�&K�A5��f���ph�����L*�����K�\��D��Y �GևT�G{�mO\C����u� BK4A�pl*�6�MɴcA�P]��?ǦT�C�jo�#�4ZJ�Z�3�_$�fF)�iZ�w�_䞎I?Z��cƤ��'�-[�)���"l������X�Fp�A0�J��mn��[7����7}�!�Gr?-�2��c!H�+� �ԟ.�|!���x>�v<;+�-��J�:H+�����q���K�Y�Ё�͔]O`�����3�l�����5'\?�G�H�����$t=�[�.�*�q�4n����y�<��]�h[��z�wa9��DD��ƴ������q��%=�d;a^f�5 ] x=a�|��U��C����$BlX�A����a��G���S_�;�
��sf*�1I�X��D|��i �]q_��ȮYL�~�M>F�!P�#�QN}��"(h��T�z�8�r�:'���(��WQ��nN���e����?e\Ө�pd"t��X4zxj�T�QyqN^�L���+_�����MB6�
#�'8�Aų�g߯]D8���_w�rI�O{�*��	E�ɄP`ԛ�&T�����v����<��gGF"�L��F�����h`<�f5̋;�&�9���-E�@��#*�N���(�Q>A`o4���a�2�;�xR�zx�h�z�u<F���`�����l�=a(�ɩ5��䏸b����0� h�WP�� ��g 0+�x�]U����\Sc�]_���{��NWU߁�$�\��*��v�f�e�ـtD�M��L��S�!�r|e��}P0�z�6gkA��M�c���;�6�m�®9��N �&(�`j���x �� +��\��,�=_�!�?�;:�T`YZk��ߣ��IC��VO�$�;�-Kkb����h�����ݏS�>U?��\�^y#��kʒ>�wp��E��W��fԐ��O���WYL�Y�wl�M��SX�M�뗦C� �L���q�zF�0]q�l�(�A�A��!�^�6�hr�\��/s^�?���{�}%��8�44IG�Ϊ9}�a��齃y˾�<��\�����4��O����"˸۔�.<�^�ii�#`��6��'��?Yv����^Hx7�9���Mq�lW�c�n#���o��F�n` ݉u�1yj������>���M��o�y;RjzL���c��m
�b�\�V�3�̎7�I.�� �S�4�d i��Ho5ʃ�~���=��������5]��G�6��|��ˆw��%�l��:͢���c0 4��,`�PDK��y��.�)���|�6Y.��0���g��9I�$�<�O��/��\�2�t�nߜ�B=>G���0ޥ��Ҽ(��B{��=�����==��8<�� ��|�y��)	�;���M	�V��g˥i���z����a܃�N=^���$"k5f �O5��*�ڑ���q%���i��j��}^Z-5�Pl�c�������:Z��ö;�#�Q���\l
N��Bp�i����X��g�%B1�֪J��#�v��E�{�U�x������3��6��&�� `d1����v��s���>B{��Z[�C���?)IdP`� �lZx@��b����i5=��!e 3�~Ǉ��'�L�>�{�	mi���X� �zx��	&mwγ-��4�c�ɣX䢖iz�8���)��۳�9�qA���]�i���G=�D�E�r�F�'Lc%売���M�)I�#,ڽ����o���8`�	������3	_�ې�x4B���#K�lvi%����R�7�+�w�Ly�VV��V�T\��fXs�����<\nL#丘f��N�xI�ヰ�2�D~�ʇɈ�Q:�e�LAn�Ɵb6�����r����Z*	4A#��/�}�E`�q�~J��DR�������]����_`�-Ů�b��Ҟ$��bN-���%�������M���&숃��#�:��䚑>�0��}l'G��,��+l�_3�s�N%�r9�*��F
�]~�H���Yf;jZ�x�s��M<"J1�l���m��ɾ��jV�A� $6�W>�W����=�.�)wèH��a/��T�����Ց�fᓄA-���}Јx���;��T��ȷ��
@E�q{�*p�6GW��e(ՓO2��R�߄k��w/��u��ȶ���ܮ
��Qτ����}���v���'y���2�Z�2R|��vײN]�?���&�F�T-��.����떗�-�C�'��E�s����s6]�k!�&RP������uX��8�rD�V:�D�E��oQ~�m���D�\��gE��U*��=rX�Ψ	�YZ7R���y�Zkp��2����!?��)>7�+-_踆�|Ӂ#��^×H�e�kv�����طw�)�}Z�"�P�8�U���F�$����S/����	Hdg�@Vuv�p�0�qmz�v8�`�֚���9W��	'��*�p�9PU�P@ނH�E3�c���W�;|�"8g����L>�/�6T�`���\�<Vj�!��:,��0�j�=����TOѸl�@sN�o��L��@�b7dj{'�����Z\
�#���.�Pݘ���𠉿�^��/��^�a��l��FZ�6����>����D�RdN�� �T�o��l([�O�zu��P+3��X�v�y��s�)F��Z1���G�4��<�ݔh�N��j}R�$�2��� ����m`���!���x<�S��{>���H!�C$<0��`�]��������ē�+Ջr���B�.�b9�ܺ�pi�`�x��jq�8Ikr��4n�4"q$��!M��o���!
}+<���j4)r�q
��x/k(��Z��ջ<�T!��{J��47R��.ф�a�rd���:p F	��gvC���3r�܊�x���?�W�M��\ZFU�6m?���Ʈn�x&V�'�������	VA�V�¶�}NqH�?.��玆q,���G&�[:<���;�ήl~iD��h��o�����**b�T��G)S%���27x����-�̈�)�>�;��WY���J)4�+A��#�~�3Qx�椧?�F_���^�Y�(�����P*H}m�.öC �����-uC�w.�:��
19j 2�����[�j���%������5T�aK��
KY�*{��1j��x	Y�����W�1C�ZRv�f���\p��lu���T�V���6�����܅#t�g��8\�& �b�!�Ｖ��S��V�픪emӞAJ �#�*������g��4�C�fD7��P�۶Evt52N��� IZ&��<c�I��k7To�,K�'��NL��ZK#���]�H���wO�o.}eRd�B��F��k �E�	�F�>�=���0p��_���
X+�O�<(D]�[L�EL+=>f�8�)r�+�i,��j&��\�O�ܑu�_� �.���V�'h����Z������O�(	ȎZ���l�X������i�h��^(�A��)���2&���E�-��`GS���m�$Șb�ދC�C�� �o�p��bMh�/JZ>cV�X�
ϓm���Z(~w�j0�l�]EXO�TY��N<��_zg.����C�R� �O����[��N�5Ŵo��-6�#�?��הu����.G葚[iB1a���w�:Y��\$�b���QkT֩�W��W������9<L��X��o�3
�Ll�7� �%�s$r^�m�ˎ9u��rhkqd.��5*�(z�	�ь�( 2ޢ�d�:�j �3� }���ɻd
M������Šߔ����3%������CXhd��\�q�[�W6T�����ȭd\b�ښ���Z0�J�֐��g��|$ݡ����z"�;�y4Ji�'pOzNʆ0���v���.x��rs�$?����_7����t�~=�'�pu|�޽�l�?�&�����W�!�qЌ]�b�~�n��:t9!���! .7j�)[���5OZ�ڎ:ߪ��7S�xZ!�;�~�]n!B�����W��"�;��I��1y��>2�����p=k�Q�"'���
ޮJC��a٥����.���B� D�o��j&[�<ׯ��,�#4X���bl�n�k�I�mK"t�X�{%���A�L@w�/]��ك��?�F�p12H�Oެ<]�l�jD`����� ��Ԣ�4crs��L
���҇�:�X� +��mwកB�9������u�zu#����&Y�b' 4�9?�[UA�s�9�.� VA�ְL�C%���~��H�W �;ǥ+܆����n�A;+�߃x�M��hm���}0+�c����oKņ�"d�X)��i,0$��A�rUsig���\ڜ�R#�S����Yw� ��:�r��MWbG��'H�� +H���Zo��{�e.L�d����_���v@�b�>?	���)?���5��/(��;F��pe��F�09>Pk=�f���]��t������1H�H��ʫ�	�eې܇��T\��P����z�*�Rx��A]=8�����1��[��&���S��'w-]n2Z8���Z���M�~��ғ,ʨ6bvr�W�+�"e�@_��M5{L�����n3 S��ݱ��n	}�z�'��g�I�8R=O���r��G�����K�qնP�S��&��yK���lZ`b��>���^�V�%����m�ؿ]֌?J�?;^Ʃ�E�����ja���*
dv�N�����3����i��7m9q��z�ʐ�׷��b0���]a�`ر=(�����)��^����7:�K�Z�JVS���Pj8d��@��:���qj���5����&���;��𚵆9�=��[`����%k�Yf.�m<O7��G�����!W��}��kGda�c]���ztO���c/��$P�3�Mia1�H���!	dZ_$�<��т�|�-�A7o�⸵�6\�o�A-Ҥ9̱���R��>�}U��٬n5驍�A��G�G[�5��"<U��S~�ï���2~km���MZ2v�/rg�x@M�h�M�����ǲ���4a]`�`�نc"'���|�h��S�!)������0JB{���(��'�E��9U���-'�Y+�)r�#W>�i�f9�KkTXSE�F_�����c@�x�Y�a�<��?M�֨�S�B �Ёj?WA���~����| k�B��Q,��~����O,`�3�ڨ#k	�1ؾX�����e�;��������xϻ��S~G���V&�w�mE4V�������ZO$��(�x7�
?� !�����) �%��V��F*w s�7Xs��)�n�IW����Ƅٙ��ץ�c�Qj:��;Ŕ�b��k\'�`��	��G�ig[�=�>f��{3�9�g�r�Gɨ���w#���$����L tbsXK&�r?�ާ�;S}Y��\k��qۗ2��O(ps��RT�q;%����	��f��`e��ڛ��;%{&#U1f��؞U����~��ޕ�fAy��vME<D�Ѩ��[aqF�{f��(xux9��sҀ�7HI���(G(��Xr}�H]rg�&V���x��B��T�p ��6��0��/}t����e�c���;����� ����J��;��{���,����|�E�$��uid'J���ćM}u�#�XH-!D�~	Fw���8�[���a��I��Vw��T�P���x�	^3g�Ԇ!@��{��)/8:�4�YL��or3�?T�����5�
,A�1\SHb<D
|$�D.��=ا�$�x��j���-R��F���Q����Y�&�͟ҘD���($�~��f�Ij�4�$Jy�S�-p_9gR�Q@(Af0E���I�Ƶfa|�.JV�E&�����^��CS:�D�w��C@��Za�P���p��1���Z��+&���g�x�Zpָw��v��V�o��YL�?�2��1@��͘O�H/�� "�Vn��S&/6�C��|d#w��B�a�_g۞�a�w����=�'�q��_�YKy�(�
�ao��U�њ=�9��Yu���9m)soQV_/)x��<dV��xӰ���\�H��O>\�܁C�X�l��5������{,�sX�ʊ�E0�B��_�=\�j72Ţ���5̲��L�.%fO���(w��lD4\��Uo�b$�e��0v#3�1��ݟ�i���'?�L�ګ,�#�J��,���J;FP"�nn�,�+{�3��i__��E�o�!'w�u3�]8�J�G��I{!�^K�0���+`nV��O�T��ɕ�s2��l��z4޶�o�뉔�d��P�1�A�y5�ޣ4S�v���7q������&�<��уo:r��@��,�ii����Y+#�K�w�BP��thH	��|&���!���6�[%�%�&���:�j�#Zg�\�E��G��� �>��+�͸xĒ�ok��L�u��)K;��R�I��B��ze��{���6�/�F5� yꥵ�U��e�}y!�}\:��&������="^�u�8q�U]h�Z}�:�t��N�h�:5 �+���%�r�N�a^��|��}(�t�`�z���Q��������B%�&��L~�ސW	:Q3�0�����A��*W���}��P0�#�%gY3�jz3b0ʫ9��Y�YZ�L
�G67��!-3��teE?�f� +i��	@h����v�������j���1)~�L�b�6\�!a5�����$�;����Z�rp y����|�p�mnf L 4'���6���2n�<ą�����s�
j8���@�g����6���m�O�w�J�Ϟ<��V��NR���D��ep�� M8JCCEB!���a������G�����8�߁���1����A��VA�i�0f�ċ�X�13�����L�M���,���H0y\(���^m��=��I���3�MMEH����f����A�M�}�����	�t�Za�R�E�A�M�8O������R���U�<�iɛT
�s��w�J}h+	B><��?h%5��$w���G���Qf�z������p6u�=`�H'{�D��D�dǲ*�]�[���
ϊP�7'�s���*6^��M��z-��W_8	�"���B�_�2<��SE$�E��_6�����B��@��͙<�@$��7����w��t+�TXr��gو]����Z)	}�~Rg��t <_��Ӹ���$����!������ώ��G:ĸ��Bs����� ~��s3*ihO��
6�8�:@fo��]�1�/!F(p���F��\�W՘�tags�/����@�:i�~��i���_u(��=��f�����N
o��ኪkfN���K����x07�-JIz}�� 츘���Y>ei��2��=f��\�sb'����w��)���9RA�D��S��#����$�t�����V�<f�+,�I�2m"��$����k@��a���78���	�J�N/ � ����ucp���XȘ�\�V� �+�>V�!&|q"�LFT�pH��V৊��eU�s��Rq�%}B�K5)H���ӯk��* !;d�/�9}��8����8�[D�_�J>H�SK�����d[v�d��jق	������"�J糏�l�����ڃr���}���ϗo"�ZJq�J�����h9�9o~�vdkP���WTy���1��r���u&b�rW�F�_@�(u�4���Pk��z��M�����cgq�=!�����>�A\*�Vkh����אX:�]E��(�P@<�/6�2�;M�h9�� �z�iŸ�@�X]�{*{&Ry��ǡ��Es/���ŐT�>����l���x���b��5���mfԞ9�[-LOb������W����y������h�kO� 
d�1��s2�zӓ�V-�h�3;ɚb�B�7�Ӵci�e�B�I8J���ɏ%��T|yA����W�퐮��'?�>�?Bt�u����q����g8cG��������b�L�E��C}ׂ%�=5]����π�T0���Q]La	�����X���� �
8<e���3[P���M*�1=RIDw��d�׍��Y�n���j`=߻�ZzGU�h������:�a�{7�Xwt���n�Q`6��c��6��U�h���� �`~�vt�
��N#�U[M�b('����H��UoET�^1�G�%d���!en1����.RI�ק�`��M
�u��O�ڦy]�������	Nr{C��P��Ǒm=`"I���O�8;��S����"Uvn'��χBW�Ր�F�»FQ,�l��i������ػC�t�q����H�h7���G ���/��
�����t����	J"C�q�O2|�(ki�(�%�`@zR�<T�&^0c%u�g-�駃���Tsc>tzip��8h�4*(�\A���H����Gl����Dh�`�N�3.�ҽ�:*,�/D���y+���y���-�C�MY�H�+fQlOڮ�L@`O�4���;��)ҍ,�{����yj����?��)�ZCm���ZǙW�������⑋j��|Jo�A�qM�-�.nF�j�F�U�{�c��bg�����	%t�D�M�_v��o�ҷ�7���L�������aϒ�l z�t�����k��k�>������`�?�y���0���Y��Ă���r��*��.�V�L���7zPkF�!�|�a�'�g\1�/L\�g��b�#��*M*L2�
V-Hؗ�~y�R��_>��>*8���u���S����FDp��;�����>��!t&J�.K��E?����.�>�I{�c{�W�{zy�/��(�1Dɝ��s8$���l�50З�A%S����;J�&�S�:��4�g�*�0ҵ�Y/��@L�� ~�M�$ G�DktP�-G��؎��$l�u pu5�XG��Z�9�ZG]?�(�+ê��/9������^.
"f環ig~޽���$;�d"d��^�=�䏏�B�� M5|I���8b�YIǓ-9�_��[#ό�ۧ\���H:�S��1�8©��])�V�T�����`۔�#Y lb�+x���r�X0��Z�o����`I.�׬���h�ؘlK1�9�`�t��/2*ե��+"���`�̮C�7Vj�ƀ�h����@d5�6�w5ge�Ӽ�d��$�.�Utw2�=R|~��)��?9W:S~֙EOZw�1W���$H	X�{NIi�C�}}(��6	ũӧj9�'��aoQ�0�o�#_��^������F|�X��9l��x�!�IF�(6��/�zt�|��FXjV��j �8A��`T��$@�{�AOc�v�y�p��#Tar��{������5�w e��́p�P�JG7�������$6ҥI��1J@Ӊ]�ք�]�����&�U�H����24���[�pK��5!��^�"�Y|��"C"���gRɅ�-�0wі���8(��|/�����}�W��YՑ �7v��Vd'�<y���1�<�.3��e$ `��p�]�X������~����\�t�h�Q?����n���B��K�:޸�%ذ�I'nX�+pig^�:�ҦY��-J1+;�D	� 	+�(�2G7@a�,?�"�C��䯹C[Ed��e,I_���'A�*i�L7lb�8R��<T��#�E�����X�YC�6�UIE����\g�_N�z���{��H|P�d���mA��.�)y@�1-�wt�_]������WxW�D~F���5��d>>Z�,v�'vU[je���VU��S��NO�tʒ!�8�C�3{=��� egC��~Pl��P�ø�V�����p[�OCx��ؐ�<E;�Y]��9Qt7���P�����J@�Ʉ�Q��3l����)���P�?�BN���I/���R����S��������� ���E�dk�8����8���4�qP�r�4�L �xt�9����������S5VL�{�J��8Q��#p�d@�ob�ݹ��&���8H��pA�v$+��~� -���� V��k̢Ӿb �d���3��?�^��zDJ'GY����L���'���k�v4~ �P^t���(�$�M�ݢ)���Y^0/����x������N�א4�T�a��!kG{1��|a�~L�k������7�|pSca/Ut�飋N���K��S$i5�.�d�e�E�@����~�B�Z/ҿr��٢7��6�f�O3���{l�zO��2-i�q)��˕��A<�"��tt	��6��P�op�Y�(�ԏL�Ql����=8_ߩF��>��B������+� �`��E8`�ER�y����S��m@���13�Ѷ�uJ�� e@��W��ʿ��L���2Ȫ9C0F	c���u��m�W�sV�紈��C%aQ� �w���'��b�
E��^-�V�mx�z�-�֌�Q6Q,�cr}����Ȏ,:��M4� ZW�;����ǯ",r��z^�Qet1Qee�.��*��Xp�J���}��R<�y8
4֥��5��v����)*����R�r��	���`V���<I�����s%��a�*k��+`#��v�M��DQ	����:8LSguv~��L�+���C�)�b�r�������&j+@b�Wj���T��v9��+r�mB�p]�ᆧ�N��Cԩ=��s��c�p#�,�\(�"P������� 6`���Q�.�f%sl���@�{��4�"�Js�1x엋t�p;�-j��^a@�LK:)��jZ��S��&�0	'� ��'��H�ves�6�J@��V�½�w��a5�bF���P����rڎ�h�Ы\�H�ŕ�H�<����)J�X&��S5�Ŵ�+W�k:4aT�;��˶a�S�l�X�&�3)��Ӱ�Tޫr*�v��hqH>���w��0է3��sS���0��=� ��	&�F't���w�����^]Q\�:��2�� 8�\;D;F(w�39��l�X��!v�B9�c.����O���W=���T�5H�G9��
`�g�2�_��n,u1�տ�Q}w�3<%�'�@��7��K�؃��Oۣ+�����V�L$[�ug�����Nׅ�m��U�v���'�_p[�.�{�EHoMo��n
r���i ���	7�J1��Ӗ����;k� � ���+�
pz�aZC�`d���9����XM��� ����#̯��q����dr'+}՗��Q�1�d2"	��T�!tb��߳ÈF�ɇ���r+�o3/�1Z�رd}fp�$޳����ڳ{�v�B4Q�!�S���6�u6��	�chO���g޽�LL5J�Xv<�K�z��}^�朌�������HI��낿�:���6^X����#5���C���	[-�rmBz�[���T�ҩ<���-�@o����C)�A!m؉L��}�$v�`��	zT�΃Rh��D�^�-O�-޺�~m�&(.�g�|'"��EC��,���c��]�K0аK���K e�6�M�T� ������d� .4�Gcņ1>��F*��0�~.�ոW�V�y�4���Jb&l֣C�z��j<k�(\f��b<�!�w�.�t��I�s�3"��#"��Zȭ,Y2?����jo�s���n����G�:�T�����̈�8S�Ε�O?��� ��w�͗���g@ِ�g���J�'�P�+��S�����p0��U��ť޳+f�E�y��|�>�{�&�bd�]��=&�2q�WoG{n[�,�!�\�ۂf�<�%�-jU)��CY����l��MF�D
���+�#0�w���}�+W3�"�$J�0бN s�)d��|X�4��Qm>�^�|�^��J�VC��?}�]�+;���z�D_�k�Ơ��s������B�8���@,���@��!Π��!ůb�//�y㻔�Z�O)�.̻����a8kpU�����T�����X���i{n�^m�zq�9	�[���V��0�%`<��bM��\Q��|M���2��W	ڦ����+N��_���3
Z�:�������L�oH��@���ם�]3O[��"�Ȳm>�۰}$��"G��;	��Z��ch�8��������@!!���~�e띞V����Z�uD��K��X���?�P����ʃj�S[<���V�r9�s�:��iB�t�R|4<����/� m�fV�ShR�RwJ
4_�JtO�W����V*�=g.DD��$5����*�Q�EB:z'�~�m��˱b��:��j!�'-�>4nMxo�f0���b��M��yl��}����Z]ֹ���^
OMJw�� �D�Bȑ�P�@fd{�7ב��<�	۰��g)�(����ԷߝK�݊���y��b������QK�Ќ&`�	L�T˥�v�7��`4�b*�>ܜ$�V�]�ja�!���F�t�Lq��0Cu^��uLq���1`�-:I��1{�8M{Jp�o�.H۶��UjW����Jw��B��F�V�	a�Yr���ao
0|T�)�SI��=��Id��K0���-S��Czv�c�%��G㨸\Ry�Gk�P�D��c(#mGl��g�L��Xntuܻ������C�)C�7�A~�Qt0;<s�h�Ztr����h��&��� aA��%y<��K�I|�D"�?x�xr��c.l�̋�C���Bk���m�
}!i
�� �V^{\MB�s%�.T�?���Z}(�Q�w%��iʢtD1�M�<�PKe�Q���e�A~\GkJo�4�c�{�[�MK�bMFD#
Ӗ�^�	�g�����55�g�08��#oL�����������N�nƴ��Ӏ�5��A����¤'����v]�����5U��U-�&���b����W�s�WR�N=�?���e���nCR:��b����� 
�2�8+d��f΅2���ݢ����{0�DyI�ďxe0^$[(�w>�������
�$�{Rc��P7�a;��~�S TB=G���{~���/���z;��R��f�"�h���E�J����M����Dݨ �fg�X���l�@�����plֶC��Ȝ��N:��W��=�1e��Q�R?��^�6?��W�����=ֺ��&6�iU�r�X%0YԂ3��(Z;p�gߖ�;K�J�I\�����[�~�3�	N�z��S��8dɜdD���eĪ\�}���Q���إ	ClW70=%�}�>�8G}��U�$3< Nl����VZ{�����V��>�;��� �a�ee7
�V�c���(�'MUV�ͫ�6��<�g0�>s(�����q���0p9Ԡ-�iSJ�.e�Qr�7�&�S�T�,u ��0��̘Kj�Zd͠��C��E�h2�V��D�~#�s�-��~O@���g��	���<���20f��P2|D���&t,�*[���f�&E�*M9q�ɾ��*`'�^��#ϋ��/:A����o�l�>0�����~�����}�n/����ֶ�$~�!Җn�ر:6�����Z!F�[���}�qJ���@��L��Q�Kj��m� �t�ۡ;���x F�_5�bDPE���zt��.}�Wmd@��5A8�/�?T��o'[�W�
͕+W���;���1����<!D�BL�� 2�v ������8���NV�1����o� [�*���������aJ�b'� iV����`8\����j<����k��+�z�LLዒC7jh�$wLo���$68�[�4����`e%5������H_�{����Kc��H!�.mľ��ɍ>�rI�s{�:�RȞD"��CS@ʔ�@@���օ���7��p����ڻ����j�.�Ub�9�qT��"��\̖yE�v�wڛ$�Nr�l�C���D�	�^M��@
�nF�k�#,^Bxv���e����	&��ΘǳqUo�&J�V�?��L��&:b��>���	��xq�r-;���	�������xM�i���2���=�@��x���I��}j��'+3�W�O��Hz�;��8S�V��,>�N� $4�⿕tL�.��jD���({%�S/0P�5����z_�]"��0Q�2z�}ca��e�ב��o%,��LQ8lK�A��:��0��5E|j�f�=��	l|g�I��V�����B�o_bM�I�3t.�R+U��O�K��X��kp�?<pM��6�N .�i^��,�������� �:������rf9$�	�Di�C�ьP�Y�KZ�*����W#֘��5ԓ�֘��]W�֝����y#�2A�D}�F�RǤ��.�68)��c�y[怮&'�
]Mn�lT�Ab�d���~�C�װ�!�m���=Z��J>�+PJ���r�Yv��}/�1䯜�G�WLs�߉o�^���-�����BTy���k�x�-wIv�ce��:$��FS�'R�2�U��<j�Ԗ������~���Κ��v.�%��t���{�[��:i���4|jY��j����~�bn�֞~a_n\w�c���!EGX�dT�J쿙�k	n�	��;��L�X�6�SӰ�h�Ʀ�*��$���͒��q9���0r�@��BI��c�Ł�5oh;�\޶�����=���~�%�2�����-�$�L!q�����u�a�����X�Dn�>p��߹~�E�C�դ/zsD�Mz���%�?�Rb��a��3B��k	xXܿH,�f��Ҭ����P�YUƎ(k@�{1o���hf���0��I�G)�G�`�kO'��)D?Z����v��Cik�!l��(I��^�D�ר��6�OP�oɉP�\F�~��F� �ǌVďuX[��S72�dV̘嫱K���7�Ik>?���-�y��6TSd%���*�>�t�G���WK�&ܨ���l�w���1��M0��_��*>{[O���
}�Y��{a��_��h�B����^��ӶS�r���ϣG�䈡�eX���(��WE�ת�"�滵��Q���-q_����а2�;�U��/-A�;�	�ty�m��T[�����-XOC�h�P�N!ΩO�U�6�]�Qg�ʩ&-�8~�"��);,�d��t�Mm�F�4�@u�����\��3��Eٔ��YY�Z�5c�r�EKvS9d{.w�U�,�m���|^��R<�v6��W|�u	�ɝ�oO..�V����Sd˶�hR�	3
����(��Mɖj�
CWLS�|U�Kײ�UI�q���nk	XGT�z
��mk���L
��>�����U�5�\�y;Z��B�����d�]Wz�(��P���S���z"b��m�H���k��9�l���w>^� k����Kc�k���{$��q��#H�;%���)+�Mj���E�ՖW������{���fP����sH���-�4?�&&߼r͙���)��ȿ�y�=}1����WhKa�#2V���L�
�ȴm����0:'�����Á���︄KLV�I����rӣٟ����D#�@�W�J^g3׀8ˢ�+�yˎ9����˳w���{�i֠��˄N�@�	����G��R]���z�y�3mt+ K]�42L<=�\9�ϒ���2т��ԫ,�;�}���l�Z$'Kw����z3F�ʾ�9rV9��\�����$h� ?��}ڭ�σK6�7b�(Ik��Q;�[�{���"%�a6d�P������Ir���=���3���u��!����m�� ���|~��̴j�b������]�2�В$�� �h�ImCy�Z
i��a�Ʋ>�q=�C�g�Oq�m���6ݚG*����W�F:տf,�Y'ostR�KS��@șs����9DT�Bf]6�EZ!����֧C�n��/a���\�^�	�����y��iwYI�.�a�#ZMg�#tc�V��,ϡ�)+�0*82y���o�9!U�0�C�F��F�p��%�e��y��-:���/�Z���H��VF��7H��k4���^���A�A Ș��#\�CRZ�ѕ�g!e?���Yѧ�j��G�Gؚ���)��fCu-\eM�/��Ń��v��D���hލ ռbZ���',����d8�@�[��H���V9��-�e�A5��8��^�;�p�$S�꠴-�l �x��U�� ���%f�I���`S�x�,O�v�=<�r�zwf
>�sɮ9���M�-����B%_��+:�Q�������	�����ch�&��#��o�+��:���v�X#��b����+Bn"OԎ�8
O3�B(�N��LM`.\.�5�D��utwi�6`�c�s�d܀����(ͺ0�1��v�H����q>�=��4m��6Pa'澺� ��oNx�[����zu.�D���;E���9g���̆Ȝfu��GV_Ib��x�,�&]��
7?gƯ�.,�=��֖�Ԍ����I��O���v/1�p�"�_�l�@xS�Y�{�������0f����ؠ?���0�X�ww.�u'J�B�
�VL���� �^���NIʐ���akK��ą��l�����o+����&�\��1wX��m��gA@��"䠱hh-�Բ!RM0�A�'��1$��۶��
rb��uDd��Տ�+��Y�)8!c�8D�z�X[gy�uxZ��~0�C�.W�ި��xv��Ƌ?N��&:&�B&.�?@,�h]�8����E�I		��]�<��@�������P��f����:�1��m��C��%>r�@%m����ه��<���x��A���$�����6��r���]RL񞖉.i~UKv���@ �}����#n�j0ZB/�������8�5]o̶S:hg8Z� =�����]��=?�]O)9 �'g`���IZj�54M������.�5B�Ф=�ķ)�;r�\�*cD�����8]ϸK��lA�v�I�>nxO�S����by�3�7�B��)������k6ȹ-�q�RW��[>p�S�"7o�s��ӎ͚�;]�aӈ�]Ӧ�l�����n��m��F��\:4��܂Љ��]P�~��]��&����c��Mb��|X�&4)z�z����@;�fqľ�N�d>�}���]���qbqB	�hU;��w?>���D�{�QZw��� 5KEx��Yt��S�7���;㊶y�|�`)����F����=L�Y�Q`HjG�>�Hp�f����x��/R�w�w���ʣ�).�O�<�;S҅M�t���u!��?ձ����(πr���O���!ũ
�Q�1�	,[��4�`��ȳ�B@��K���?�I�L"�z�X��0rJducc�Pԫ;@2,�S���[i;��&;ޝ�����.U��F���ܶH.@X� n��)It+�[������x58���4R'4���vZb$k���ٶ���|xZT�p⵺�E���Vw��d��}�]��� �#��y��6�&��11����Y���D����8Vj�7o�����y���Z��������O�H�']�	����G�U�1���pZM�d��Ց)�-��������}8!a�yQ{�N3�3	T��rӪ�� �b�Y!m����\�� (?���E��1r�������~P�zk������t=�R9p����}�Y�2P1Qv/�,��l���8B	�Cs��z��t���
�xxm�
1�`4��5�<�}�vq����g�\��M|	�rl��)��
v��T��̛��+ o��D�Y��5��t
��T/Q�|e�˜��c�����&�����Z�Ewy�)r�������(���)X_bk�,S8%V���@�3�Z���/��ͨ �EC���+��Q�S����2�)�V�d%7��T@���N[A�o�S([v�^Tmn�N�c�9^#G��� M�p�V\���,��A�p+D��N3o
⃱&u�X7�<���Q����:�R6�k36eh��,h���_J�������P�S����|a���Yb��/��H�b�����~[�[P���ɧf2c��?�Y����fГ�YBsέ�>YI��%���,��-�E�'�j��-����N�.��k�c.�E���n�]f��bg_����$�J��3@A�����t��TN�|��F�mq�`�g����8�˱ƍX��? YȐ�f��י��lN�|/>�o
��lhh�<��+tU�3% K�` �3�ºuYF��V�
mm���,��k�޷����>[$���0�Xh�	�~�v��u�Q
kT M��R/�_�����i�m��R�X��Fhn���Z�W��ݜ�-u�c�6�/�.�|�"#���-8�Rf�e��u�Wc�����8|2�������{�>�6ֶ�<������F�h$�\�w�b������H�B�r7�đ�b--�䍿_�UR��"!������9M��i<&�i--��U���`;����1 ��+�ڇ�}��+f���̗<k�����\��V*�P����gү���䂛ۊNt���'<�oZ�+;�Z��)�^oe����ۖ� �to߲�U���&�P��Zj�n �2e�/�ߥ�e~����	�̏���n�]$��y򇜧�5�����b�(k�,�k��Ւ��s�����&$@6��^:�ݺ�����~�g��u�d���1�� �|����	�w4iSd0-�s_�V��\4����2t.�\�Ӈ%���44o˻�M7������םQ���q�,tj��L%P��S[~�;N7����?�r������w��"�p)����p�!��Cr���)҄
����"£���2 v�9��M��Z��%�����Ȓ	&��2o�f��_6�((����w���ꔁ�� 4*9�'��T�g���%a2T���z�|8�;+�m5��V�����E�� `2�0Z\��Z�%,��FT���j��bHEPۨu��
���DS�����]	aTz��H\����8�9ԅ: �j*�ܦ�>;`���>L%:�:S����&�� �%�բ�n�Q'�U�N
8��Z)����f�dp[~/$YP���s�����(,56��fլdd6���o�*��K2>0w��(e�`l�t��w�A���
o�ň�B:�W�p�tz��3�^��N�^���G��@]N{l�Y �IC�>\C�GӇ���^[ ��z|��;�Oc�;���,;/������![��p�6bω�8H�v�q'��׌tѿ�1�����߅��{S�Z�)K�~�tC���2PW���]�(�Q��i�wG���Ac�u�\�^#���+���0{��[�G���L>�]xK��/z�cY2䩓�x�tA[�p��fx���5tk�<�}��R	�$x�F���㋌2�^Ԑ�<l#��M$|�PؘM5�v���X���$6o�)rEN.Q�5�=,�*C���~��N�߆�V�3��^nlI� ������1������X�u4��4]k�npҒs���A�A�y��\�ГU�neC�j!"����`Ò� U��Ũ��D66gz��^�ܞ�):��l�h*�:#$6z3!���xʽmZ$��Qq�F`�l�P9y�5�a�_�3�2-�)AT�P��y�5?�?<ҷA����N#�8ݬNŮ��`Q�/�}%2��?h���"/U��`�LF�7�!�%�{O��_��Np���q������F@SY�kٌ��*�}|���ܮ���3��b ���[˟,� ��]�~��1�qѾ�0��-��v߾���;*��g��7NC|> q�\�?w�_�K!8����D����3��J��R�v�f.�e�Q��[>(΁���*lH��AS�u��C�ւ�A{C!M�8��@#����q&�)�J␥��/���J�Y{%O���h�Z�Q����e#3�49�?�gE�?�%���1�0w����Z��xD�y��sKI�������a�����P���A���U��z@�����^Q�N�F�_ә?�[�uE�~��+zH�*�7���(a��X@�Sn�⺢�:E�ܭ8��1���f��}Y���M�'ǌ�:;.	�,��9S^C�z�����Q#+���"2kA�̞C*,�UN�&��*��� ���u+��g��L��;^���҈j�s8CZ��?�!�ֽ�m�v'R�6];N=�����D�d}���C(�|�)��X&&Fбlv��ڻdU,XP�S\Pڅ����ң��֑~�	Sg������:)8�]�n_G�+��_�ZC�yAp��X��K���Ҙ1}�\�=ukfvE/���)޳ �m�ͬZ����*��������T�ɻ�r����ƺ�B(�;ׂP�8<�h� �iqB��g��J�Y�`�gġ����|�e�n�$�a��0�q>�
a#փL��%���m����G>���j2�.{l~���oAk"��l�L%�6��Q`�hy�E���E#�P)y�Q�����̀�9�R2�������gl���q�7ï	�WZD�a$�͵�虝��ug�����X^w�\�A�쯉*l4�33�Sþ��+��!�u���Ü�`sn<��>��c�_t��wN��	���Tf�	�QZ}�Z��h�E���F�2�����Y�`��|���ě������k��ȑM���fw ��G��{�
[<+R���+�&ˍ�^v �m�=����)R0�#.�� 4�$�k`-yw�^D��rC'�9��L�۵�D3Ep���y@ٜX�bs�0��94t����_4�7w�7����~[l��R��P��~*�Z�:���Я�Pf��5הo�VG%Y5�,J�ǹ� 0�.WhX;s*�gX�:yW��՜�kÿY�խs�=��
2'�y(����[b�<��`��xbR-S���kI��C�oBv�V��d�� �8�&��5��->��Mzپg�R �DYGϜ@m|E�/9���P�i�r	��Ϣs쑌�~}����<��2a�%B��( ���؁7fD���,9��m�y/S�CaD�x�({s�U¤֞q�_��������̎E�/�YЏ˃�gק��4�v�ۘuT�~#�q��� ����/�8�� 9��k��{��:nYW�6\��?|賜�������l�QR�0�@�K6���ſ����h8�V��	*�x�!������];2q�gʁ�bC2�U�a���pE�%��ە�!�T�ZC��in䦧��X���)'�:+;�N
��|���-;>֚IA��ή<]_�,�����N5�ئ̈u9fD$R^���D>!ӣE.ρ%�F���z�;2�"�ױ�Q}6`L塺����#7r�������W�]�?���a��G&&�n�(0�"PFz�T���v4��z?t3����=Ȏ�Dze[�ofE�o@$\��A�j�_��!v�jՁ�F���]}\�`��X�2��b����ҕ���_�&�R�E�}����<u�9�s��8н�h]�$������ޚsx�7F���V��i$�����%��e��<B��p<A�fzf;="+9�I ������j�� *�mɥھ�I�|� ��59��C�o�5����?��F�<���������M+��*'�,��`���wB�ѷo8�3�5[�\u�q��۝��"�J�H�v8���v�G}6�dw��'�u�[�l�'��P2;W���D|��ܑ��4����n�t�������p��!�d�·͸�|h\��l�S�� ��O��dk��ԃg������Vd�%�n|�B��)�;�[�Q O��'�	j|��I������d�R�-��SG�	OA-ͳc�62+�eg�^r$
P���H�%�[�-I��)��
A�d�����Շí�P�K���:E�89ʤJT����E|�e~J�S&�B5nTy�e5��纵:�w��+(�y�s5$�^�M�� q ��w�z ��)!��^/ւxC�3%���6�z:�>-ڛ�.=��O;�ce�i;��u.�:�	��Lݗ��cR���Ts��s�n�M�0^L��߱|��YF�7��Kj����OcU�.~���U��|�AӬW�
��� ��cxmm��@�߲�Av��O^Ix�=!�� �tm��V����\�3��XnӅp��T؈��~�|ڤ7����M$�Oðז����i�ev�����D�Ȋy�hOS@m����5�%T�$s.�R��Sp�ڎ��G 5IS�@y[D�L��(��,�-͖ S����x�����~�)=rt�QQ��x�4epOVn�"H�H&����g�����&�^�5ȉ�1T�����ЫuB)��d��j��SqVlz�JL|�Mb�rM����}�L��Ou�;�i}����<�\�3���`[��|WeXUQ�#'���{�}�u=���B����9��2�j�j���I��˿�� �A�dy	�T-dO�������IR.�rjW$�J�Ҟ���;+f�R	=���5Hq\|�� ��ڜf�����Qc�qn _�LѪ�b���O�J������Ȼ�����2ˬ�tZU,�e,�ڰ!��&,ð�"��6��m��F�d�w�G��Lg��w�p
� A���n�>�<�x���G����� m�$K�z.kmu���#ḫ\�Hc��̇D�ۅ�H�y	���ו @��[�pN�D�����˪�;nO�E�q��A�����$9�ހ�#D0���b�S���o�͓�F�\�+���V/&��z�r���~�F&&�y�UYF����Y`�@9�g��I���X*�+���Yhȅ'C�̳pTVM#����k�o/'G���"�t~ؘ����;�m��`�$������=�������E��ݸ�'x���7	-�%[�Oq�F�-��
��d�L�d���z��� w@|8BنÙ}G�,���s���W$,q{	�ڲd��I�^����sS�5��c�ڎ���?V���A6����`�b5��a��,4,��F�E����	�Q,Lzx��Z֛!�x6�$�M��A��rB�ց*��_�w���R��q�����vG�=Ì�ށ�E���4ڻ���v*�|x{��Q��O#ʑ���j)�H����~k�˔��s�(��G�wve����8?���_�{�S�i��dф�8�th�_�l`���R`-�hX�#�Lat#^��]ż0�H����u$s�̔���/� /�(�_0�<�}x�c�&}�W�FJPް
�[9o�(ȣ�@�J�z�c�X\G9o ��|ў�!�<]������r����P��E!��g4��뗧u�uH��Gh���0����n�̖��(O]�2�p�����"��Et�IjGm������q5(�^�}(X�n3��3�E���NP�h�F[�U����k�V���A�H�uJ�ڎ*�_��-p�� ��A���n��_�~{��-�k�Tt�����:-޳|B}�U*
��]�w��R�?p������R��i��8K������˟'�^WS�R*�.�7�1E/�8�����}h��]��k��"ߧL�B)d��)�V[N'� x�A8��a����	Т�����7[]�n-�8֥K�n�����qi�Q)�˖0�JҤ�Vh��D������4�=+p�qz�H��X?˥�[�p!-�F�B���Wx��y2��ZyR�n�52j�;)�V�Au�Z�mDd�`��R�r���˜�-��� @oZ<�Z3��4�{�pT��(�d�,�Ѥ�_.���13W��^j�?�ゑ��`�h�I����������\v�I��NtkBN&�NE��%(�wh)�/�#m���R�G����V�W������Mj���l�d��l��m-֏��`,wA�~u��Z}�|�6�rtxd=D��D���o�m��ޝ6\
gH�%M��>���F�Ӻ�U��|����5�?�����=�Y�x�nśҊAf2��B���ܟp�⍧xh[�I��c��9126.�=���B�`qh	�#�
�����݈	����[gg�F�fJ��������k&���' X���ϕ�6����l�z�4�>g��e�!��ɾbbx+�1�vi���C[������џ��pg��w6
�P�A~��/Qo�T�2xH��{�S��򒏊�Ky���U��J
d�������m($L�omQ��KDt7��qO�^���fI��_�+u�+�9-�QRAֿM]N���������;����J�G����%(��و�+�_���}Ь�_�H4�&qq<�'@3n���Q��G�1֒�0f�n���u�D���o�}GPlE�$?�������ėqT޶<
r�����$��d`�Ҍ���a�+ @d��hςɜ��1�,�G��� 7�I�����2T�~o��������=�x-$�� 1/�^+τ��Yuʖ�G��k�!�>[M�`4�૞OS|���y��OO@3�-,M���Ŀ���N����{e} �4<�&A��x=@��R��i���GO�^�J�G�S�9��}�F�a����~k��a�J�5��ݡ]�i��K�t�M��2@eA{������p鼽tCɚ����8�'���:�6f��gh�[(��Hmt�|]��W��.�.��Yn����ߍk׿r�'���]�:*ޗF7�-����V�o�ã%����z��R�Ԣ�Ǩ�p�O��>`�����������$��	�.�!X| �'�;P���.����Ð%���ؠ�1�[9�qt�m�n�b�W9jzi)pe'f�	Lq ���h�_#���ɱZ�Uγ$i�skJ�x:�Z"wGd"�'�EJ����2{KXo���p��q��|�w���	��6�5���/͖E+�]m��#Z�!��k�$Ŀ�闼b9C��KO~:����82]\���%!C��q�t��N��t�Qd��]I�Zb�`�&3ʹ*�UH�7<1نf6o���w��7�-E���5f�8�ԭ�+W.�{��&C.��~a�[�������g2\0)��~$cq�t3 ����A	�ic��;���κ~�"0|=V�W��(�������&� �>��7I�r�,���w���^�C���ꀝ�=W�:���,�9Z�����cr뀲+o>�w[����9)2}CRu�RcLK�t��7�B���h �X�y��Zʢ$cݗn��)^���}T�͗�>Ka�AGQ���8K��v���Í�ؖ�ݒ/��h�٭�X@�"0V��M��%�b�7C�	6�mCu�>�� �%��P��!X���yYȮ\ފ�
� Ǚ݂��Y;��X߱Kd-�27>\�K�숖e������
Um����[�6;�A���
�NU�}��.gsF�����]���2���sgW	�2�֤rxK�)�+��zV���\B~u�s����[��6�n+gK
��--+�ԬI�����@��䎹��
^�QS��s��v��P�����6����D[����P���FԞ�(<�A��$E+���u�ObloLD�t����?Nw>�3� �e��Rr*A�1��%�ՀA�_/0���������7N"��u�3� o$\]ۻ�RҩD�w��k�_�p�:щ�Xym*�k�p�zI��g�(F�l�������� ��;@��%���[��@H�N@��K�����uH�+�����X�\�ub��	�ִXBϕr�Xq���1`����!.u6[�UΑ�����/�tMn�$�tq�����;��9�a,��mo�%����Ó����`<���d��Dvr��9煺h0ԓ|N!�O���gfFX��0=�L��;惙&�� �@JˉX��rg������=-:,��.{(�87��t��G�E��eeZ47��)lJ}���noa�֙�{{M�m6�U��C�/�J��a4gB�����Nh o�0������4�Q�����-�d��J�~�P>��+��{^p!�q�s˒��}ڄ�*�{��K1�t01�����,):�h�'{�@����rR������KNOic���I�
"�R/5��1H?{���+j��?��H������x,zoߴ{�{_���UY�6���t�n;Q�����缴�g՞���x�ay�
+���1�"�o��dJ�b1�[�]�aY�V��ְ��N��̉��7��r�]wQ�N�y	\U�՝l!�?�Ҟ���m��s>P���E��ϗ�9-�k������ ���'�N��VQ>tv�A�]�O���0�յ�즍�{�w�@��+�$�}�9����+#�w_Z�nyMBu�(ג��f�3�]�@���ֵV|>I�[w6�'�t�Ɓ���u7��>�W��{��)��R�T��T �[6��W�I�v��Y�2���C��g��p/M_>m��@vR?��n��.~�7�Aj�#R.��G���$Ìdog���^�M��
�����f�C�aV�t���:0�zO��ywkܓ˗���<,�4�F�����dw�TdO T��Ed5��g�j���5��gĔfG
Hf�	�U�__<! �$�����e^A��m�s�m�e�M�� ]�ɮJX���L6�p�pݛ�2*�=��8P�ا�Zj����'i���>/�[�	q�x�i��wS��C>,�;|h�{}���fAe~it2m�s)]��I�����9�(��A!�_��h�($��I��.+�^W<�ݨY-�a�#GB)� b��ԮP����O��1��";]����J��%���j��;���SK��[I����8T�]7�w\��ޡڞ��QU�K�j��7+�Wy������([�����.=���6�<Op���2w�����@�0@/a�������kŗ�q�c�)�����߷ܪ�\�f���z��}[��8�&�: ��|(Y'�{�H,o� ��P�,[!�B�kŭ����n���9+���œ;���z���Xo��U�F����&��?��W��rn�P�{F����ҋ��(��adj&RM''b{Y�k,R�S�	��9��z��e���@dN���|��m�O��0�0\���{-�g��I�S܆��J����/(>���JB;���V8�c�)|�PY�^��3�H�b��0�(#{R�1;���N���_��t��r��/�s�߮����H�Z\LX������H�����
E4!xni]����܁��[8Ux���@�Ռ��i�R��F��g�;2��Ȣ�W(<
I N�HE>Oݨ�y�$����ls����A;��v�o�#�-�"aLM���4�!ʢ��%$b�'S��q�]XE0`-s+�E�'k�b���J��k���%T��es���Ug����#=xj�p�+��&��6��u�����yf_�s4�f]G�G��> n���XK�ޓ�����6��Y��Z�H��8�]��<+�L�׋����s�g����1a�ߊֿRr�^p�f�!�J �W�����/���(�u�pO�Y/Y���S�ml5l]�V����se��43h�~Ҋ�0�E���~�n�J��ڛ$�}MTu�p˂�nw��K��U$ؔS�j̙!�%h��Ή�[��æ�H����[�Ҋ��Y����X�����sW틄���i.J bT.�k>��k�@�'Udq6�v�,?L��kW*����f?��)����Hl.O����5��
ݧX��m���i-���/p��P�*�:�&;�s����X�64��v��oρ�&ΦXrE���/�����X�%�APʱ��%�\xv#��&#���x��d�Vf^��C�`u˃pc蒷�`�?���ԧD�@��ݗڍ�e�X�~��%�c1�?����n�.���@����*y�J'��*��g��aB#�/����}=�it���D�#k��=(&�7L̓�92;�S��V���E�h�p����%�R�ð�Մ3�q:7�,��w�`Ӹ��"8t���.�Ű��4���f��p�?�÷����	�@�@�]�26M'��$���<�R��n�`����VK�S���/q�tʢ�-�'��R,�K:�U�������F�/��Tφ����������[L6u'ń���
�{�-�d�=��!�9���>��������bx�3ҕ�jbܿ�<�@]�^�0�=��O��ra��|PJi�J�X��b�1�+���!({��kQ �z��tbR����$P�����'�OB��a�mX#���`��gPֽ��24Q���uIh5B�L�?�O��A.K��\o%ű�!��l�\]@�m7�b��B�֫�++G6�� ��P}�X��j514�L͸�a7#H������C�Q�V�A`���]�L��K�&���Rq���/$$���J���1:G�2�Ha��;}g	��z��%����BO��g�^#iPlQu L�9<���iX�D��?_i����_D�P'�E5E�I���w*IE�3�'G��.�5X&��O������Ԏ/�\K V�J�x[|�K�eO9���;g�v��&Q"%��97����K�f&[��D��w�H�	���pn�	d�\��g6�45�� �8r�=�q�C�X�A�)�9�������W����hD^�K�r�\�ϟ���+�[�����oM��&�d_�W��U���-�3����q�NJ�����r)�	��~.�K ��ފ���]��}p %�U�r)= �I���B��.��憎��'+K�1�&�;.��q%�"/�܁��H6�Xx�	!���֍k�����������ٙ�ј]:����8(�{�(g�v�F�)nvl4�n���!i^�_q�A�x� �B��T׿��s(`�^58Lc���be/G-�?���s]�P���&���H)̨��C�����$<+�\�ǽ[���r�:,�#}蕤+y��%����|�@����0o'���"�������)�c.�]$���B5�)њ�è�C��*�@%KY���R`�,x�o&�pdP˻�W�H2�\۲��]�QPG�J@bX܁�~<s1+7�	�����Ee�g���ɟ�q�h_�@��
y�JPn��D�ʓ�h�%���?`t���)(�(�̳A�H�zN4v�{�
i��`w(������߉�@L�g�v�]��%pݼb��&�wnm�	n�Yׯ{1e] ���D�}z���iQ�c�["x�B���}݁c�c{5(��0��u�����;��f�r㪗O�F�j��h9(��jw���D�ZnB?�������ر���yAh_&���L��hꏉ���Ec�;�2����^���!	��rE�^X;��m�$&G�A������GqM9)�U�!c�U��~∼w��Qv0�Q���N'gLêV݇��
���ϵ9�w3�nta��S�9�^s�����P=�<��%�\n��� ԓ��a���D%�'Z�������}�%�P��@�'��J���l�vVGq����X��ʁ~]V�r��_ �<>�`��e�hU+b���;�+��M���q��:I����G!�;�K5�K��Z���a����3�N���K0F�K�r%A�yg����,�x;�$s�'y����)wd'�]o��Q�׻�d'ª��h���B��Fh��ٮ_em�q���.w���$���{G����A�5Y�(��=�ӔN>#=�{@8�Ż4������gQR�}7�z��E�� �!��e�~]m�{$�ީ͇. �0\���9?�܊S ���2���h4	%�����OQ �N �C������u����/��ԙ�^ז @t�t�j��h�$�n[E�{C�IW�>�*9�;�R���Wc8GK�-��Me�Ν����m�X.�dC���g� V�)��!4���W���?c��ʐgY�Ξ���s2r�v�b���k䜕9� C�:;t�<��l�72�f�S;6�
.ɔ�m�s�i�#Eڏ^�����]1�F��+�%���Y��eg�(D�1���R���.������Jg	�^ *��=n�xn�bWDGR�'j(�p�"������`+����7��F��'�����VVC�G(#S�J���UO�{���d$"�x��޶�BA����N���}�P�]�ӌ?l%'҃|�\�����K��=�y��q�^��`�(n��Om�Qj4�C%��	� RKx�4zz�n�g_s��k Q���St;#�Cc6Gd����'v�	u>�T��9��d�׫g��A��9�3?��E�lb�U[jn�C�X=��f�U�qgI�,(� �L��ˮ_#>��#}�<�~ (�W�����@��c����BӪ0p?��R��K��ͳW/:^v"q�"K��!�����&�?	c�v9#@��̻b|dp�;\��nS�g$zYN�b�K�bVd�)�n//���	�n;V�t�
�In"J���1�:�c����k~8C�5��`�}�&4\�V/��c�.
%>5��nZ>��.c8+q��.��9^;��`����������\�����-�����\��Z�����-��J|�l#g�eф��0I�����<�F�(r��@�i��	3\c�|�$3�'J��=���,����FZq�o�X��ZN��Rj�=?{�ɯ<�+M[�I�H.6�!�ͫ����C�KPV�>�퍩��:��7��?���Nپ����sd���p.�&z� �}F� �4O�(��m	����U�|���w���O���-�-f9 e��_U6��W���f������P��y�53zTp7��+��jH��-z�ߕ�������3��rŁ��r�ڜzN@�Ef�Z���c
r\�I�[�@=����O'n����������ċ�ka8Foy*P-��eo1C)=�K1M�&l��Q��P/�?Sx�U��9������ٕ�.���h�K��i󒑡mHSDO#2�d\�%*cbݚ�,��n���t_|���R�X�n��{��Ǥ>'�h�,�'����Ԥ��I � ��Y�E�JRu���(6i{��u����Qk��2Sqn���r�Y����>��Ć�N��`b��i�!\�"�Y~�"w{\b��k��ٲ)T����0!?`qᾚ�U]�{���R�Y[�e3�'��^�ň{D1�G� �ɩ�)�G�D?96�w��H8��|#�����`��t�>�<��h�?8i}���F�lJ/�ʌN)i��w��%X�]��o.g���r�Q�ا�f>����=X�SvI�+0���q�x�%Jz�����6���tLZ"�ރo�w�g��c�7���R�V��s|��_���El*�e1�Q�f��Wmt���=E�\��0�zgI�l�+��N���x��^a���\tc����x_�^I��nD��J�9K:�CJU=z?E_b�ܞ	+���2�im}y�����{��Q��r�zm�M_x��Z����@P	X�E�&��%��Yۿ�>m%e[���'�R�< �4�C68mӲQ�j�qfn�n��]i+��S[�3���C�a��K"n��o������W��
�'��ۑ֠���?���\���"��&����pA�ȅ�duihE�OLsú��H�acT�W���t�hw(ahL��Lн��P%Z�1�����g�a�ڋ���9����vǫ%��5yȌ�V;8Z��˱���K-�)C2j�9Hup��}�8u$����y�ϫ�r���oojhQR6F�p-�	\8�e�w�s�q�g�
�|�NTB��Ϛ�Le��/�tQ���%�(I�,��\%ѪM�Ls�QV����~��\�3�)�ݑ.\�Y��������4��C&�h�L^��f�v�.�z�ʸ,�����v@��2]c=�`d�0w���o�*�1�)xBM�1�F3R(�m����Hk7!^�w�i3��/&�0&��kϟ�^��h��©b��N����f�D�mc�do"Y�5R ��-\�S\>��l�vD�൰�y�8�i��;F�=�� �~�,_ߖ��N�6X�9q.$�����n������ �a�HťI4���8X�D/o[Uvܤ���#"ʳ�A�8� m�Uy�����K��w/,C��N2{�iF�p�E,0���:�f�O��2��*��_� �r�o|FK��'�e��bυ�aHv#���2?Ӵ��3�����3'���w��tq����	^����障-_�d��1�0�!P�`�h�M)|`)	8��}��Wq���4_�g�+�+8����h[1��!�{���༣9������gb���$C���6�h�=6��{�S�fDC�3��JH>[���b�uay�k�+���8zq�k�ج�M��|���{bX<����e��I?#2�l���
���N��*�����S('0	\�[0��*?	��U��)��4�����^T���e�du�m�Ƿ���+�́�E�%���/ֳ�"��x`�K5�$�u�rl��cGjDhÌ�rS�ګyB�=o�?cl��Jy�n��8O��k@���2W��l���S��g�(�"t�Kg�7)6R�����'�H�.�9�q�G�{˄�,��˚ސ�80��H �xA���l��ǜ��>]���LT*��}���Q� \B���977ϋ�ן�����{��#*V����[��8S����x׿�b?����@�h�q�B!�*�V���������P|�����/�>�����~��n[`���3%��pN7�,���|�Ɋ�W���$��L��;�Za����瀔�A2��;aKn�_�0$�|y�i����Ȉ�`A��Z�8!�0�?��n[_ͽuM yo��=N~��ϣƾ������G��o�^w�(ef��Y��mS���yɉ��'e�s�J]�)t��{�χ9e[��0CfJ����t�<�d�o�T�:s��4J�'��l�j�<5����W��e�@pp?�W|}�:�ϧ��!{5�73kj��I3�L���V1ӏ�r�,�y���l�o��!�n]!�(�s�B�`w��� a�9�{ok�:v���&�@�^��:`��Z=�J3���I�bt��b32i|�T$�p�oca\�zH!45i5s6�v[A�v�
��݉X�oJ��z�����R��_q�]�[����؏�/۹��r��� �p���ͷ5�)��l���ݧ|3�ߦo��7��ȘX�H���`�����j�x�{�S�=TY͵�����1}�
��t�7620�1{�I���m�r�S���}H4��.��TwJ�H�m�Ea�4b}�������a"�Jk k�6�5`��R�q)I��ՕBs�o�ф�UA���@vjT����>���U+�"���O�歉XR���a3^}&��EЙ�:����&���o�gZ�ݐ�pj����#?�����+m�
!Y~�T4���m�l�_9�w��^{�o�՞=U�u����e��dثdw����ԟ���(�Zٌo��	/T�ϵ��?7���#_���,�)�H�5�{iЭr<MU�����-Q�O��xr%��}����R�Lk�YɁ�.���N����b��d �3�jK��C�&�A?Vr��ڝ
hH�q��|U0����"L�l3�.�јdW�A�4nC0�!�2�|7\oSo� E���!�?����? G��u?m|1�����R���K�!�}:��-�4�C���[v\E-N���^�T�޼v��2��f����F����mL#YZ�I�!�1�gOx���Z�)��XilCX��)�`���LĥV�Z�ZD0�C8�!�\9.��*����"oN#f���|���6�/b���7/�F�:x�O7�.e���=�7��Φ��E2�{7���f$�t�'�[�h)� 6)��d�s;>�թ��:���|=y�5��[e1�+�#�5%xm��7f�QBu��9���>P�:15v�}p�{+%6/���!��&���(���i�(�[�b(88��k��N1�XO�F<ߧ��~ua��7R|yt�Ꮖ(�\\XG�^.�'�[�4_�թ%���tז�i��5���<nR�'�T�7<�Gs٧�}���>�AІ��b�Y�Z}�{��	'mGB
MU$��L��L �#�TJy�D�4��c���,܎�I�Qn2���i�24�_e���xp�#�%��U���Ժ_r-�&~;�hA��]G:?�2����~�B���
敋�P��F�� �Y�-��p�!���6�C��"�8��8?<���J�#%�C'�0W�F��a�j5�3rZ�+&�p�
�gѲ�� ^�Y�y2��؄���F�EJ�m�x/���Km��u]�������(�p6����Lu�H�8��M���`���BC�q��=�����;�:�ۊ^���Q�-����F��0e�dQ�и���l�7��v_��#08�s4<��@h��n�	�dc� [��B����Z�n�$QPxe�M�ߵ����?� ;�Bp��R�p���J%'�سa�}��xe��j� 	��!�qh7�[:���W�j�+>����\k��|To���#տ4e�xn���ǟ���hc��4?������) �9a�]yd���S�����xH�O��]�*��~ls@*v�64��`x�V�'=pۮ��wf+d�|[�G6���Y;S���i*�0�Vh���c_B#T�xk	gޮ
�;2�	O��G��t�7t��C��RIqH�%�-��˹Ϩ�|}e�9
`���Ʉ �����s���iX��%���bV?�=7���vPB!�^����0��T��Ý�DV�v[��v�K����r����+�(��q���8��;�BH}D��m���ka��,ov��_������H�`,[�b���`˯�����?�<�a�i!�i�~J_�S�u�$�c
�6$)�eQ��n 9�d@�gj�|�ezh_z�(�6�?]�c\R����ʟD?������c��MEQ`��ԭ�.�q����8e�t�Fk̚ɲ����|�Ɓ�B?%�L��@��lf����3>rJ�i)Ҝ��m���)�X�B� `�G�ꪞ1_|Ն~W�ą��7H�G~ဣ����$��)�0��c�"E�As}w��l&�ٻI���NzW���y��P��;�����!S�aQ��>%�:.�T�A3�W�r�l��@8���;�zI]y�Q����$�os�df��ɏ������Q�#�b�+�ؼ����:�A2�������m��� ���Q�y;������߀�J^q�(�/|�ՙu&�ҩ�a�]�@��L�@#���4q����Z��Z�������L��Z�K��B��v#��ʡ�#�b�my��*���6���D��eE�K�*`,$��Z>+��?���e�E�O��4��җS��=]���[�~�a6�X0HT)L��"gݟ%h}JX�ӵc��
;:͠�w!���,���
�Z�tDqtօ�.�i����j>���9��{� �@j�1J'��ZS*�4�+�L���ik�[�ط	��MD{P���a9��Sd{tx����?4OS�H�;�I��o�FH�؆Ћ�ˬ^��\L�Dɘ�V�J{���
w$O�>�� I]��#v8�eݖ-�������R88���T�4�RJ*�;�gY��% U����d�R�=EKs�49�B�[�Ǻ�-��q�W��J�P������.O�06�şɄK}��)m�o7였0�%�Z�$��Ս�F@�[	HJ�ey�^k��w�ͯ)j1i~0���Y�?�*���km���!!���/ �s�((�d�8�(K'�D��</f�h�h��g}Z��tN�t���B��e�����J-$;:��%�]��
(&�T�-�@{�wP��U3�ik��vNi��^Y��:���	�y���i��:1�C�/D?�5%;D��H�����8!�][<���q�Y�9:5r.1���]��	��}��XY�"Xp�0�^�iI�ţ:�/��.�*]�o��7���(��O��Q��ڕ��w}qR��ݝ��ۄyԒk~��f|$6��{�g��,X{�+�gʮ���E�0Uo����\�
��.̎�7�&0�P�a�o�:�uNT�f��p�=;˺��t�;����Ьu���Ob�¨E�N_-{�r���%���#e�?�T��kw��$�"�����nщ��}5�H���_�2˯L�O���*��c�7^�I�5�jf�jVW� GE��l�^<��g<=��m�0/=QZ��?WM�8�������#D��F�����0�(�(5�[?���\����yP�jτ��r��c��RC=RAK�e�'d�e����ӫ�`
OM�]�NZR}=i	�Dp�(��o����*x��x�3�07�����B�����&O��x�o^܁��:<ގ��=:ɽ(�llhB�4\�m�������fW{�0��S(�3�JzTI����A���薿��,:��(&5��5����PS>a��޵����g\(YL
���<�"@�"��u���ݭ)4���0X/j���13�G���`�`���f���V%�#�Ľ^\�W�ۙ�!��2�p�:�����T9kg��
���zIoO�'�����R������EGk^���id:d����7B�%(������.�l�Q�HǗ�%�$.�2W����%�l:V��nm��+k��0^���d�a�W��$T��Q��������cά�v�*3~��>�牦?�֋�Ƒ�˄^�|����<�۳��,���d�?��:�@�5=*�P�js1��
��R9��bg��C��oL)
)6����V��]\�ܯ��3@*&���!B����<x@�$_E=����;-M�Oł�Eք��`85.�f�t��Z���[.�]a/i��<�Sj��D��/)�n���	_�\���vP#��y(���@1 u�G�xa1�=�����v�Z-"�9��*�(4��^�3p��`MmadZv��f��~B�D��YǇ�]F�D�gr ����ք�оi��z�"5�r�V��k~P �8�)ҒcXh���t}0�����)�_<�݁�&�j�)�0��3�룢GS0	mg(
��|��oH�	��M���ߑd#[�ǧh���椼�����)����/HjZ�р��?e��Υ{��Vӎ�~�$ck!q-�OQ�g��?r��
�zP��ۿ_�e��Q����h���C�ˆ{��ns�<#B��o���˝��Z#�,�N�2����/+�F�Ô�||;Th�PeM9��!w�E�>���/��f���� =ؔ�]<�缡��l���������Zr#F���^��Z��_����Dx4|���P�^QF�LZ�[q���\J��?�VJ�I��m�o�%
��
)���Xע�q��7��2f�i��.;�EL>e�!Q�.@���A}P͐�����_��F A��ܫ�_> �ZmF�Nb#�4tҋ�M�^�/%�� ;�;�JK�䅍�a���4v���:��}����s:E�7�����Ő���0�ڑ/ը�b�X�i�QM�)yu�,ݑ'�9�ig�����y��m��m9����aL)���j�I�԰k�K@�$M7��L%)�׳Euwdv�pR�[�9� @͏Y�{q�F�ӈ?�q[J��E��{ζ3K����~iH.{��3�/�,[�4a36Y)#�,�`�2.����Rp�գξ̚��]����ۘ��F�"�<춍�[l[�������sw��[��Q��}���X���yMwf�FW���>:�DOv����r��Б�u�]�}��H]r�����!rٖ��H����zk�-�*m�W��qd�j7�����\>�y6@  9�Yz�t��8���arb�}�	<-yŶFn�
Kl�Č�F!/_=��[~��{^�i�I�&��*����e�5�\��B^�T��,��o�$������1�
+����Q]�!R~G���l��XT�hW�:�L�j���,Um��ΨP�Կ����A��,�eˁS����w�C�p�B hOæ#d�lG�IwS���aM�_�T$����ג{���'#���T <Tb���Ya�	��֟T��>6Xw}.8]S�FEY�������rH��'�Ӎ���LV;ރ( �������ڰ����������U�z3o���D[�����:��Y���l��vǁ����4���0�"/��G��VmA%��M\b2��3i8FHɻs�tV��;��.�~Q۫���$/�-S��~3���r�ܑ�������cT�cJL �i>UϘ����*"Ct��U�0�Ц��z��+��p��<�)8���u��	T���]���Zg�YH�~C��,_|�NP�6k�j��~�BN��;*�)��3����E����p���b��s#M`j�� .���g��fsK��xd��☛��/8r��+ߙ������W�\#��iX*T���-�l�	�nh��pcf���,H,<K��]�wh`�X�q0�T��j��}B�^��!�Ï���c!� � J�4�f����`aL������
ਣ��8;ǚ�g��\<!,q��4L��Q�vC��V	��8�������*�b��؃�m4����Zʙ�k"LEN<����7R��~�Ax��z�8���(����~��È`�o������Ҧ�:>�H85:�/&�z�=E���CL�N�Mr�,�&���5�
[dbGQ�zkT�x�WȮ���*Ƥ���W*u���r?��	UR�����)�q�ˁ�Q[O��_�kkB�.��)����˩'�2J��p�`#��#��
 ����Dal�ih�n'���������dZ���>�y��M���ʌZ�5	!Ĺ=��т��r��'����p����y��j�bI`��i?����� �v�`N����ׁ_�!�6�u�3�T.�ʾ�Oa���|)vGeI8�!�6�FI�"�4d�>)�6�\h/&�[�O+{��K�y��QN��;��~gb6Fnv�J���4q�[��t��	hh����wr�sc���{���l��Q�������_��9E�ah�B��+󦰙a+��^'!`�j�u��2�$|�2J���U'l�&Ɨ���D��˕,�g��u�y���#[�M��_��xj�[B��6 -\�8>�����ˠR�V鿫�)����wo��J|�n$���L��!8��,xq�g����/����v�J��H����g����_ɩh�^as�dzc�������#�K���e�+C<��xd�U,&PC�����7�/��F+q^v��ۊ�^��t8'^��!|-��m��A͓��W�j�(�D�i<^81����$]���g�J1$Fv,3����*�jT�,~p�,o������~f�tBu���{��тCN�㊄��X��\�u'��[n�y~#�v�.~��&Q�K'NŧrdӔ�����qC~��q�-L��V&5��-�QԶ"�C�oI�W�g�0�Dz@嚰R���y7���9�C^at��~Q=�'i5@o��\Љ��u��>�H? ,��Aˇ���*��ứ�,���HE���r�Ty�]�lh����+so��	l�\=�P�o_o�U�(hh�Q���u/N�ޓX�P��qS:�}%0��HS��a-�I��!j
�H~�+��h*�.��AV� �������|�)��ހ`�j����������Y���"a	ZN�YZ#d�q���ɫQ��[����_�|
�$�$n>ɓ��2_�������_[��&Lݖ����|��>��@;�!2�Q�6ʾ ���h�ua�1���퀩�KUW�)����B;�=��7'�yo��֎�� p�<�F��������)o9Xf6 �8�A:oP�5�2��y�e��9[�\�n�53"��Q&ք�納yA��6�Z�><{�D+"�(�}WM*�v�]�Zu ��q򀶛,3Ud��j/�̞�t�Nt��6�u��m��CV�!�\E�Tto��¼۝�a�ȑ��UX�g���$�Vk�Ȑ��޿z��*��@ η��Ēg�Ji�A�?�d�!����e4T�H$>���n�*1$yw�v*0=W��{玷Q�'�V�u��l��q��W��Lu���PP��I��_��\9S>���~�`�Aէ��!I/��wGy����ZC���&��G�IV�����2>�4�9�	)8�|d'�;��3��"����84��@�bW��[��p����>�2�,Y����ς\F�iȀ�T�%$�be�G:����~�@D�����,q�h�4t6��eY�q�8@�t��&��s �5�O�����~Pp�-�ؾXg�RHM����
�w9���
qj����%+S��B@J�!~�B{�6�0�K�)�dl}~�(�錢!2��96�|-�U�;P�8s��x���HY�|��dZ3m�S�M���4
-4�t�z�yi�E���;p�Y���Ia��ÿ��2�� ��V~�Y����⌽�K����O�b���I��S:D2��J�wٸ�����$�٥����<.�vw_�Xְ�rIiY�!2+oÄD����޽4���N$1+�5�v�#�G����X���F���Cy�>X[p_��8���T���Nw$��m��������=��U�YB��!��2�4�c<`�U;y�Z�N��V�;�#:�/�s���
�֌��$ܛ,~ķ��������<�	n��q.��U����d)�HR�����l�@o,�z�(��Ae�%�*�Yލ��k�1�\�sU(���y٧2#3��B�������nc	Gި������J�:[�Z��ġa�W��[�������M�`^�fE�Y�U��}9��u�gY���:�RZ9΢��Z���j;@�*�'$'��	ۊ{�H�q��B>��g���V���:��o1��#�c���?�u8�@�)��߄��ߍ9�}���!J��˗ \�m����������E%3Qk�]�aC���=��<��7�b/����O���)!u��Ld.8���wh�Tb��~��w.b��,�| �S��rU�#ʉ��Ƥ����0FR����V<^Ϲ�u������x��I�Oi�λȊ�r'wߏ��YR���+Y&>�zo�piVT]�� ��Y�D6�K���}���2{b ��Ǡ�AY�=�F R��Ҫ�0B(�'|��Wf��5�LM��G�5����ꢌg��2�Y������i�FNl�5	�c߂����9�5��o!u�
��Д��/����2#7S�駏��L���,��r*��ݙ��1����p�86'�tɋ�狺��X����8X���[K����S��ݶ�PG;G����Ӱ!ǘ��~��k�<�k�bȮ=�d�^,o�0�Q�I�/o8��f���h�j�uUf�s���C�	�� �-��+�(V�i�ۅ/�	��>'^m5��6���U��J| ���ڝLcn3G� Nv�X��ι��uN�厫��� ]o�O&�^fs���An��-{���Bu��suÒ+ǈUT<�E�M2T����冯����}�6���+P5�����50 Ld8�{�%
�a�A��ف���`�q�v��'���m�'��^���:�0��-���G��Ǎf�O���F]b�v�7=9��.HIT����D�j s�����=�=z�pU�c7x)�dC�\��>\�t�9f�T���g�4�<;�=X�;P/)�K��.�VkC�e} �0�0�~L������x�ς ��� D�����鑲��cў�E�C�q��M5y۪ѣh��U���?�TY}Q	߸����P+"���k�埋 �1,`�eo� ���8�gE��W��P�^�G��k���t'�ܐ�w��O+��]j�X�R�N�G���bR��n�ܜ6Y�6�C����벎�ѡ:� 
̋�&�h�Z��m_I�?��b8��q&�f�ŵ��]��M
�V�'Ik�=菳lݶ��Ճr ��H�[��A�+���qޜ������ZI���/��3bt�Zj����W��K��E~� �g;��[h_n";.Zh0�qoH7IET�-$���D�ӭ�&]�+"�_�l��������(x?y�,��nb�GL+��+8�����6�N0�*1l�x�u��-;�(�yUO�.�B�!�����2|`��M��rx����i���_�_1ay_�$�;��%F��N���]�a�P�CT0���`���	|�B��	��u^Zcb��)�k���3ysE�t�$o�T�p����'>1�R� ܬ-e�7��Xޅv�t����ĺ���+L~Z���Xu���w��,W&
����1��#F����Me�J�DGn*�B��CZ��o:��D�1R�JLF-���,��}�3R�;5H�"�&Q�Q����A�:cJ;qd̯�92���1k�S�kOU0J�YQՑ��'���z ���A�|it7W͑�_鵞�=
@�˙g��l.�g���GQ�L��+�3%��:��� ��ƫ�9N.RC�x)�������)-[L�R�8l;��3f�K����:)��n��~�)��[�e�iggA�]�}�N�
�,bB�I#l�}8C��S����a�#]u���E_e��J��F��_$�7y؈��>�0Ɏ��[*y@^���%�rEեK�n���%�'�nn�_ΛX�-g�²"
��$<B'�W-V7:1��Ł�R�h%颫?�C�o���m�¥��N�-�e2!�S�a��{�7��'�=� �rkG�e%e�|�:aHDε��I����\�{�;G�!R�hc�Cg����U���<��f���k?>�;I�K��p*�����W���O��U��Z5��O��͗Cn�isps2���^}�Fͣ˗�����c0�hsm��e��L��%LX�Q��_7�lelI�W��H����i���<l5����i�ziӈ�j�e��|ZKb��hJZ�zӹ�=���&����~����������6���S�Y��a�a9� �`j����XH|n�t�����)U>�x<r���3�|M��#7� �]�S�`�⹀���V�)O7=�S��}`pjLƩ6��9ݗ�\P��D�=��6�;�m�����{��8l�q��>�B�����c�&@ߢ,'���yp�>�M|���7�[%䷽�t%w����N���#z����KE��J�rFZ�7���^��sYO���l�)�g���v�Z��!Ħ0����'K�6讃�/v���wK8=/�ܟ�\j_(%�N�E~������bo�r��jx��L��p����3(O��>���5GU�2t���*����wc�>ɨMA]�:���o_C9��>/�Ɨķ�\���.�����������Te�f�9(1J* ��5Si�DȽK���RGB�|�hA�΢W��pY2��'�wh+�l~��)���23\0��r�e>G�ƿ����֋9�j�QK��yy���u����
�,�5Q�O�Pm��U'���T8�ar� 
D��@����{Ѳ_op>�p쁇	�J��G�y��'ۂ�L��VfJ��wn����I��zh��5ƛSi$�Cc�ֈ�G}�r�y�f~���g�,P����_ME�<����]2%��j��2�94\�5������B�f�36�уtu<�7�81�� }������A�� ���u�~Vؓa��2D��n�Q]�s�'��)�*w�%�s��s�ox�m#�Z�g����LO�\��WU�4G���ݭ��J�O��
s�,YL���x�]�<�`V�̂�X��ׅN�5yk�dia3�>G�*3YʆW#���e����];�|j����Li����FT�����D)�����E3`��eMfcC�XW����uN�l*,=�$@\g�1�f4��=��Brs08xD�����i�̍�w%&݋2�іV�\����bn���rZ��KS��2�rF�3ȫ�]����%?B~�ȴ!�	2��`�O͞�ȑ�Ǩ�{��̢⼄	������;h�h�f,����?��"�0K)?Q:	���������zm�xq#�}	1�zٍ#G�ֶmg.��,6��H�n���e�z0�>C��ܼ���X��˷+Y�ax�e�p�f�b"�]�����e��]B
�sU���P���W��E����n�рm;,¿ ̬K3���wW.i�-�q��|~��	]��rZ��+,gψNl�����/��>��I)�����ִ��.�Y^�kGz��*TG��T�7j���������'��ec��d��]`��{E� ��d��%ك���"��߅^z�yX�F*�O�w��L
hf�
e�<=�ה���=�1�	"�D)�J������7�^�Ï:��}7%tT�6���!���ّ�2�*�����;��^EO�??�R�iv<(�Z����iT�\'���d.V��o��A�@��q�@���b���(X��k���<|m���Ϥ��=�����n�Ŕ�6�Se-���LX�.���vD39�ra��p��$,)lL-WK@��x�x��yϿ$5t�� ℺��(H~���_夋��oP6��<yX09�,��I�Xi�:���8�;��∨E7�T����-�@��HsB8�}L��LZh��~�	�5}���D�wI4�<Li�E�q�5Wh�|ԡ^�za����aB�8�s�צyX���e�$Uu���*��~�}�:�[��1u��s�����D�?F&��md�M�ʭ��i�f{��ڠk]�o�?,u��anRr�uL�X};`�Y����J��o\D>"v9��0J#���E�2�*`��L6c�!�s��>�_�M�L�sΚ������w���<g��\R�~��(7CL6װ��;Ka�]>��
�P����8�{�E*87�)� ���%.唈��:�a�����ҤJ�O��^��>�(�Q<H_�����4��i�ƪ�u�炇Z�]�� 5�wW��d���n��P�ȑ��c�j��WV7�8�t������/���@ޞ������xUÞ��G�R��Z�xh�:
w���?����5D4k'%b~W�"K`Z`�qa?`�<�+�dҺJ��v��x���������뵻������"8�E ?d�Ҋ&d��}?g��dj�sO+���,'�g/澸?Ρ���>�Z�Q�Y �4��ֳ�k��n�ύ�2�L0i�E���t������BI��"iDK�����q�4t� �2 �g� �ժ�r���A'%>�}�mέ�y�WA����sfs�T�C��B���3��������`�vb��Q=V�wY43[��hY�����*�g���2�Z��������4����(ÕLkbc��D�������n��sCFN�7�g��2E�Gȟ��j�%�W�����>�8&ъErM�RV��q|2a�;B���d�hP����wg����&��w̀Fx�1���Z�r[��5k:�*1�vz�Pڐ��.ܔ1��$�K�c��!^L��d͂}�$O�֋���0/��f˥42wɌZ������,+7� ���q�=[c��X�8��cSg!�����v��8�\�x63�Xf���M��50IFK�a��d��9�x��g� ����Q�b;l�ޤ�G>I<2=����6�~�ص�,O�4�j�vȔ]	z9�y�i�j3���쪵���!e%x���y�kв	���ah� ��̯r��SAFiɅ����0�饔�zQ���9bu��K�~�9I��+@ϴ;Z�x6�]�q�R���j?��h{��[�<5S�Ƌ���ah���Gz����X��y�m�2��N���?p��{ P.SK�
�h
�.�݄�z��[�Y]���B7!QR�z8�*z5���zR���a8ף���;��0f���B � ''�� n�3w*YAZ��;�x� T#/�ε�)+Yfm�O���I�
n�j/HA��#̢�p��h]�x'滷�a���$����Vh,���>n��0ʺ��O�Vky��ɷ���y%��DC=�mꡌ�C�����&�ѱ(�r��R���V�@���9�������^�hJH�*��,9��#�W��Ȋ��2�$��0xP ֗����O�Q�7�
���T�*��{H�7o^���7K�M,Mq3\rG���9?ц��c \��!��e*H4����"a��$ �W���� "h�����5�FTE�UIZc�ճw��2a��d�4N�EbZ�����T�q	�n�F�����g$��Ĝ�;�!M�)�څ�]ʾH�U�q�U�tg,�����8v�x#Ԡ�̍]�!t���/��\o�s����W��]��O���r�E_�)����ޞ{�4���u�y���{H6����gn!BD�r �R�oj��J��z4�\�N�71��S�S�FF,"5�ݨ3���z��?��~����A�{�H���4c��: ��[�7;�,U�����ޑ�aO=�b!l�D��j49�k�hEE�����%�cS� �y�@�z��#��7D�h�k���*)6�Z}[�$�Ф`�<%�G��jU3��S�[�!k6��N]���U�Lp���|G0'�{I ~$�l+)�@�<$���/�]��?���v,�_kb�k��IY�������?1�ȝrb�����9��x �h?�t@�s%,
��A�0��^�q0ш'��Q<��8�aK��Ѳ�XfN'�Aq�F��L.�u	?h�J�.�qr*5��1J�]�� �*�g���6���S3��2��F�׊q�UHz��p?��Z�_e���*�-���ѓT��� %�W:B��IRs��=�p+͍��ȡ�ƕ*����g��*��_HqU<��e
 ^�0��$�{�E��qNUxn/�d��y<��v���rXq�{*��~ϧ"���3�d�x ��.e�{&���<
#B�����w�$o8V@/CfȲ�<�,js&B�a�����TŒف;����W���9V���s�ܕ|6a?��� A���Gv���أ����}����$|7Y�I1�I�R��v ��#X	+���c^�l3�T�-߻�#n�tt\�
e"�>����)(DX�R���,!.'(�Ӗ�"�{/��A<]��7h[0Z�{���2à ��l��7�@|G�(��$���@�mpa�% �x����07���8%&�y;���2����pƦڿY"��c��Csc�U<W��ݫ/6y����ZY-��������P�v�?�"�O&�54�JL�$�D��V$��:Q6�_����j	ȁ�Tң�ېP嶰�����`S	���<�2R���ۓ���e���0S]�sk�Ԣ�m���0B�����g����Q�s���۟@)/JmY��`Uz����5 �la�g��c���� 4]�\��/]������(����+*~�B,ݜp�R�N]�b�ӱ���j�L� ,�)��N���t��~���N�?Դ;�(fۅF4}�i��I=���K�Na�O;�Q�~�փ�m]�;�Z8�?�����t��i��Z7��-pR�82%��]j
+Xs�(�b��vJeӼ��N#j�7N)�)�0j~�F�
)�S����,�&�������[v��ҧ����nV��� W_}�G՜!s^��.�Rs��:q��B�Ż�.�RO=�L�3�DP<Ť��3�kZ�ܐ�?dT�<l��5´�FK;Y{�F�F�Ӭ�%�5t�c;����/m�����}��l�.RwZr2˻m�j#eJ���ˈ_�j@�3�;��3%��h3��\%��ո�m-
:m�[ձI�R�׌�$�J���F]��y�#MT@���Ŕ�g5+�97��r���y]� �%��x
�lC��L��4��{�ԉ]�3h��ԯ�ѵ���heS�R�G�X7�1�Ji��J@i�L�	z)>
�����b���0����ieZ&�ql\Z�:w��'�1��}�P�%,q��=���N��hI���1��~�U�0��r�N�*��ؔ$�!���/YfT%��_�x���C����Q��&�X��p�USa$�+�y2U��{�X�3?M�0\�>.��	�yJϑ�MO?5���+?��rB���g!��}[���?��?*��R1D	��|��&�����&�^#ik�4�qKԻ�n1}���Z�ءI[quB�$����=�<W�%�Ǒ�A��_l<$�1�QZ�ٔ�+r��+շR����t�����*{`�\��oʥ*�Zɐ��]?x��u���Q$�Ω�v�Z�McSl�q�22�ID?G20x�$Q��8��3�с>Tl�"ޡ#o��@�:�P�#���� 6s����*CXďI�~˷�@�X�@�i!}�xD��`,��I��K�jA�p��m�엨�s/��;x�'h|�ܢ��YY&VM���	iSBW�bۡ�t㪑U�g��'��=�S������5əQ~7�ל��r_9�:�qk:lrܱ�	��չqG _�{�" n��t���gh+�dz�w%�|#��\#�/���ʬb�FI)�Ho��-c��oi�V⛿RdpЏ3YGCp�s*W���&K�4�y�Ww'm����Y���$�z��.��Ei����},*jV�o
DBauX�m�/7���e���g	a�un!a.��Y���s�0M�Ox�vxHb��{���2y�ڙ�)j���]ćw��!ko�>�W��n�l+y�xii
.Y��|�o����ݡ� 9T���<c��������ך
�y\7^i���$�k_�Sx��VZ/F���5<��n�zp9���K��> h��֨i��������������֥�T�3-!��i�:��h�)WW�Y�憨�&Y�D,S��ρZx)_����T�U-�^lm��f�R�0l�>�7�����1]i��<�� {M)+(!�e��������U����7�� �@���YW� Q{|�{OW�}���N����t�@t��;Qn���#μ:�]�o�4hY��Օ�R}R�p��H�Y����<r9�S��=Z���ѷa]��� �Ɖ�?�Y[�^= C���lvTY�M����d����Ρ%;	\=5K�-��󧐣?�F�J �L�i��y���@��������r�-p�Q3�qH-���vR����d�]�r"R�~�q>u��.7���;��#
�<�H/���*�{dĨt(l����\�j�MTdn�sM�vį�{���d���Y���0]M���K�ث_�/.�/���[ �n�qi��"(͝D�] �?nL�M�M_9|�@��:���[�BO��0���c)��m�0�U����o�x�e�}5�i���"Ƃ��cB��A�6*�<�&:��)�6Z�:�Vl��d��ؖ\�� ;��C=�9G�j��Z�n"T7���r�E���*AT�: �"E��t�?�9��7##���0 ���ݕ�ӗ�!�,��0���|q&�*���x;��B��e�R�� ~�ox�b�g�4�&�]%��6��t���9Tۙ��
�j2w�*��
h|�,'@Ô����Z�B�A��t��Y~����\zx	o�B�Ai{6�3IZ�`�kR�����Hu҂:�FB� #e�Η�P<.٬J9�6@1�hwKp9=ZV�t �^��>�4R�r��1�F���oQ�'�|�Gt���S�of��[ڣ��ҽ@9�#ޥ��waȅ����'!��2��L]3@���:�
1$Z��>'��tO� �s�֣� �('^�!,XM��v�#O�	����_ v�n?��i8����L����2W6;��z�9&���
ǹ1RZ��C� 4Kv�0wjya��S�����iA�n��&4B���}7��n�5,�y��P&�~94Cq#�v����B�G����:�x�2���Ԥ<�.4q�ڼ�9�`�PNM�3Y�uM���HY���T3���Z�K1�Ft"�&i^�-:غ-�x��('ڡQ�E�E��ݦ'WE�F�9ϐ��g�|n@���U����>Q@QE�*�`�!�l��1�z��6h��lp�ܗ*i�1�P�QՕg���ѵf���a��I�|�
��
��fL��~3�/�)f�bI2+Ԍ�(�ϟ�FIγ#nػ���iU�I% �N?�P�ә(�~Q�JՁ0*�H�ԓ��dU�x���!B�"��,����?k:��*��s������Νs*�gJ&�a^�X�񘎝Eo�"3�����N��[�
=�M�E�����G�k'�_-�C%J���u��?���*hAoD�ɬjae��A��oXA�G�+Y�p7}���k��6��OW�@A�_��,�_���,�H��UDWp�x��b�������P<�P��rћ��E��������p�k<��]�a�bU��R�6�}ZC�F�Oư ����}��Ԭ8Yc���?�-�(�S�"�Řv��3��ӤH�����W���i��L�Sb��I1 �92�����CĿ�uK+����ɾS�~/���ڧ���$,H��w��z�"��wG)�s�y��ՙ ^L�E�c��;�*�V'��p���Y\�q��t� )�<r��ݠ�v��1���j~&�fi����v�8�R_ 1
���7R�F���:�5A���6F��H@\�t���C���[�]� ��2��uZ��ണ�_ �,����}��)O	�JcHӳg���؞�
O��5�_q�G`�<+�Xl:�u:�3N�� ��W��CĐ��yf��9��)w��1
�A��=���^�j_���Խy��`�0��$�0�w�$�+�x�:�R��^�	�!>m�C1�
� ܰ'�X�$��~�h5$4�r�գKz ��6��9�٧r^s����`a4����|���H�!Z�0�$t��刜v\˩�����+�Le&�������U�D�-[ �̦&5!/a�*EGOЌ*�*�`��"J�s0�3ǹ�m;�) ���c�`�o��oS�|N�6	V	��\7L��_%��,����3oӨxW��)�{�m)�;*� �>7�/,���?*��k���w���� �ǆ���"��a�'i~��5S�>o;#ג�Ǧ�����*t2jZ�Ύ��q�򨄜g�&S��,�6�����I�>�� ���"�S�nR���n�<�ߵ*�i8z'6����0O���2]웯�LgZ@�"3x}2��@�}д�Yl�kٌ���DRm|�-�M/]�*y,�	M!� >%�P}9�%^�8��=�~���E<P�Ʈ [� �t�,��K��v_j��Z��~�#�ރ��z���Q�`�R��S�$ħ�[֘o�(ky�'� �9�]�kVQ�6Oݜ��wEՒӌK�/y�X�~��TjF�,ѵH�z�@lw:D_{�Z���K���o��:p"&����u0W���)�(�$�ac�Ĩ{�3���S�w�����?�Չ�y�&j+^��	*K�\�����+��w��˗d:zbV,Y����2��'���1�V��3�6'w��G�{�l����q��sKqJe1�y�Kǭ ��O{�U�"H��9gD?����:n��b�GŦ�:�{B���*Y����˼"��Nz�o"j�#Xu��EՅ�i��MIG&�Ri�h�4���ޟW;
�ڟ�~|[��J}�[���04Sa�j�w�"A��6v����5��\
�h�����)�Mxv�߈?��Aǟy�g��$l�E>MJ��6mvv�C�3-���:!0櫋xh�ں�u��}�v���	R���慘�D���A:���Fw��kh3GJ��?#7��nݸ��!*���pv��P�=�P��C������,O�ywɛ�qTZˊ";�K*+��c�47DO�D"Օ�Z� �OtM�n��M���
/ܟkB�v�y0v��9�����M��Rj[�i�� �wѼ�8 8������������,5kN�i�nLd�v��IIˣ(T�[g��'�2L�7Z,��͋��;���E��x+-�����`V]�f���	����@��^9��7Z,[3^��^͊�l{H={d��{�ʖG����R9Z=dn��"��"I� ڪ�9�da�Y��{)N9-<@��H�띙\����%wc���?�lg��i��4��h��)�����he��#Є�U>�Fb`x���N�)�T)Le�
�S���.c��-!�80��Q�B7u�a�j��F�4��D&��*1���qW2u �����cz�dˑf@|�s�j1h|�V27�V�鏔	�Yݖ���O����!�	L�?.m)�p�翥NF�9����ҩHj��}���(�f	v�M�*�p{���:�b�߆���4x�������=i�3�$O@.�v;�;��lz��U6���d�u���AW�yV��L-
�����K��ǼGڥG�	&rN����w��W�Wסu��^��>q5?{�����*)ڲ�-�B����:D���1>��8DS����0GkLm\�+t�c��1}*G�a<� KN�@�-��:].��p�O{{[�~��|+�L��{y� J�	-ت��9G,�6�y=]?�؂>+�h�Ӷ^��4Ⱥ�L��'``�*�D]�G!�7If��R��yI��>k���� ا��:�Ǹ"�5�Pw3� �����+v��TK�Z3w�F�;-B0+�/k=�Rz՚[���伻.@����U�Y��$xJ=�����m���Ui^qC(���r��' �)���b:���+��_�6�Hl�<���Y�٧�j�6���gͧp�"nw��J�'.S=_�S���k��4R��+�~;����zQ{�P�!8�"��b�Ջ��;�_�X�䍤���<Y�]�E��='%l�P][R��Eyl3.���|�HY�Pxm[�=R Z�R��O�Kd>�O�����E�9�����v�(h��w�9���*ϴ���1͍#0��'������u�K� ��q���#6h|��k����X�]�;�h2ʓ���/��Kv�`Z�N��T,�ǯh�f��>`��A�Zr\��'9D�O�4Q-��	����;��^>'�> ̡��j�`�y/�b��8 �[L���oj[���z�>����!*3�����sD�P<��@c����L�rS��)णX�v׀A�~Fa�Ŭ�1v�}�s)%�I(>q�;���VdJ��9v��ٕW��9����\k.���м'*=��9�juz&��YzQ!��r��F#z$N	�χr*�U�O�&��0=}Qd���B`;�IHϳ���nmB�a�v�Q�h�Ǖ�����ɞ�����6�΁���b%�c�q���ן�����&��N��vL.%2^U�x����H�t��v��j��0�+�=�ZFҟN�.%�\]1�d�j�\�B�ay�R�0M��F��	�3k�'��\ a�r;�W	��eo���?Vv+��R!�a��4Z�]/�mؾI�7@�=0���������R�VX�O�a�`3G�tGK�5��A654w>�}�ٿ�|�J]<qw�I��Xw�a�*��t����m��B<+�
3��ީz��T},*���F��� �m�n��"7h]�lX
GT��{��2�fR��ޥ�u��7�(��Ī���}LF0u�׭�I�s��4���*�%�vh�=~�u��;���^��43L��A5Xp�~�ɺ��&N�z��2T9���oh<�)y"T'���on��ߖͨ�0ӊZ4�H�1c�d���IM�v��u ��V����2*�^a��=�~���Y���rO,�O�{#!���Kp��-Wܺ�H0�t��8������`Ks0�RW�f�b�/��w�4�>8
Y�4Ә�b8�4���Ʒ^�#/`�6����y Y��)��ac��n 6�@�'00ӳ�1�zu���]o�j��7�L�B���J���w���-HɎe?h�b]h�������(Z&�74\Q�i	��=��uY.d��t����qC��#n>/�2 HI�H�&%���)��[�b�f��IR5��N�,��#�&��*�l���E��jCZ�I�a.�U��G	�I��g�,�����H�'-�� �tBLh"�T�G�ܡ����=Z�lQ��q�*����j��̏��\ݰ�14Y����PwYj����~8sg�ƆR� LIQ��Z������dq��D5u&�Q��q�>K���2�@��(�P������-h;�	a7�hS�n^�]]��}Ղ�r�j���(���qm(��]�D������������%�x`�#�q-K_�U/�fp,\�\��OE�*�2��j�9�p1���9�;���A�f;��-�O�v��
��$B���H:�0��W�S]�}�J��W��c�����[�Fz;�k�����s��}����͗U�
E�=Le�ōS1�1�(wش��=ȏ��mڈ�, 	3y;k���w���V�>�uMZ��Pz�)R\��*V�)�Ap��n���i���_��W@�6�8Y�A�/�`חr�<ی,���G��-� �a�U���q��Yc#w�9"_7.�h�@�~`��|����|����p����������K������.q?K�����$�W��7���N�b��4������_S��Qv�	,
ig<��6���\)?Ǥ���?	�ZD���q�e�B�5�r�s���%����;"�2�����Ϯ�}WA&�m�.�n0��m0r�b1�������f��
��5�2#�s��μ�v��HM��pi�T�6�b�WH�?�~�u���3u�iA��c�c��ъiN?�GK]��Y������T�F�`5u���W����
����A.R�bz�׽kq�$#b9��9��L�U�lߞl���=3ɵ��LC��`lH���usX���N�wɜ^�3�if�R�	���� ސ��Zy�G�Ms 5��2Y�h��y���)�� ��Xǿ�5�d��������j��ȗ(	x�6_���H���B{'�m��z^;�tW��l<)cN��I�����M���c��~����8�JD��������O���F��d.]�HH��a�pT�~�������foB
1mCw&�l�K~�A)%�Z�q��P�LkئK-�࿄�}]1
�LFO_�f(���|K�"*yx[Fw�[a2M���� �����+�%��Hs�D�Л�����i�%P�CO��`w�t�e�#Y�Df@��SQc�`�p�3o�"x&:�g)R�
��<)�ST��)��t	�#l�uۛ>4%;�Y�����:N6� nWZY��E�����?���mu#�Va��*�!r͸�'b1��������޵:�K�l�'�]ufdm�0=������̶�!�BC����ӴǠ�m<�6��H c�s�~A�e"C�8�	��H���n3�J���^ؼ�k�c�� '�2^���((�t�B�n��(Vm
Y#���dxg�Tfp���N�%�H�T����� {>���� oPm������ne���a#����s��8|�"��E
�F4C2[�YWa:�a�Y���[dI��{������/f�5\�?�a@��fyx��O@��m�,��ǲ�:�G/$��3��s�>����	��e|��c,R�o<��[������Jf��C��"C��i7�(	W+o��J(*�G(�fm5f�I�~���fN��y��x�:��w�J8�j6&��vO](�OE�2p�
���y����T�<P�r���ǰ��2<�N�8I2���an&T#�~|�;�����.V��3�����0����8�3S�X��0���p�q�]�j�Z0( �'Xx\u��3���j����2��4Z�k3T�c��9�����x�~���>�"^��ʰ->�aO�/�&�3�P�&�	�����ēk%��; Z�-b��jU�'�a���i^�l�Ɇ��b|x�]��n�B����h�WGnԴ��,�9k�΂!�7���~�&[�)� �NN��j�JKY��)(�t"W����Ej���( ��Z��z(ڧ�
����� � �'��ځ6�4?"/\�Hd�|�_?�y�AR\� ����G�'ê/eg����[�^Ո���ˈ�g�8�O���u8���l����굓��+:V�ڀ�*�ք�[|&����]�Qg�����2:�dU����{�T�a�[�Ȉ��ƚh�^��y��a_�' 3���5o��بF�@��k��E�����i�0�Հ?�d�>��~�ˇg��#��Kr:d��%W���6_O'a����"	�YA/����s(ܻ<��c�~�ߝ����hNՄ�ٷM�.��+���n-e�A�q�ȣr�K��Su��Ra0���D���0���?{/q\����$)&c�i
�Ͼ�h�ɞ7w�?;�z�h�:Ay;Sp%\/#�X�d�g��?����9f\�� �����.���s.��� D��6oB_��`w��'e��!���rGM~��(�8���@	9��/��Jo�$�!����6�)�cN�H,r� �Ϭt/�7 6)?�W�N�	�t��ͺ)�(E��u�E%��Ӡ=���1�W)��W{�r٣����gQsa��)6�a�:�{03�4��B�TjJV����;5K8r !��)��#����Zπu��Q�O�3�|
��/?�G�oY��}O���)*?�T���������6@��y���;��G[Y�#��AD�(��Z��p�+Tǔp9�s�DI���!bDuX�J�!��_����ܝ���_���j��x+:*�&C>{!�����Fjꊦ��n��ϥj�1�f���f>�n��
����q�4&)�b��Sd�Y��[�Z��X�Q�.�!��D�/�%;j�T�n["H钞!���IҴ�qYD�y��L���Z61�4�UD��ƫR"z�<X�ꆚ��W-v �C���\-���հ�I�F���"���(�,� ~W(iT�Ye����3�*��A���B��d�����Y��O��tе�y��b� �[|�M{٢f-�6�e���.����q�*��Ѩ?�U�F���W_�B�L��K�8^�GE@ �C$(k�]�N�s/?~u*�Vx>���W��!���a{�L�
��G��.l��~C�\�Z�?~��'�ފ3�Q礐����y��<K��������)�;�n <���P����!Dz&�q�֯�*��<'�,���gd̻�oH��iY�K1�@�F���h��ڙ�B�T�Mi�\�u����X�h�p����Ҩ9o�-�flGi\c�&.J�L�W��>�h�l$w��M~����0f��B���>�`�݋��}ga{r���c�%�
�6#�t��:�C��G�\� �<��	e:�:���`PB��/OGe�&5���2��ġ=�j�)��P_($�В���N'T������G�fλ�~"?�[�,P�q}�P���-+��s�Hϟ��/�^0ݿ�Q�)OM1k��	ɒ����m��0��� B�1M@b����&iē�q����j%0����0��v�;�j�U�;a_��G�&���Rcj��_���7Qw�T_@�w$d�J�l'�P�^�{{S�G�q�R�3�7e1؈B�_j@y�\���D�0�R!��o�����<<r/���{c���� ��m5�U �b_������z�!2��^4+U8@B��򯂾׿��u�T�YB���������{�?;u.#�wry�;���;����L�2�c̚�^���Yx";\�4d�����v�/���� �qN�\&���$�Z��~ɓ�)�T��7e�8-e
����EP���Sg�@B��,\�q49S�7t��I���@�+X�'R�9�#	��l8e�9^]��uk`��s�FY�I[� 7��ּ˄4+���ŀ"���Ew>����@�[���ό�$�4��\�<(�P=�l턺� Uyb�U.�X��,���ڈ1��vM��O\�<����������i�+O0�5R�:�!4���Tm����9��Y�+��ū��ey��+�C!j�I�X�Q81m�e%�\_�5M^1�b@��j;&�3ⅉp�*,D����3�h˓�c7��Ab�(��H�۳.����e��'�"�b �n3��Q��ǒ>����2�z��f�7��#,���O��b䟱�� V@K�s���f}Q��T�TslmbuFe�,�+�h������#G�o/�]���wؙf�T��^P��;��e���F�W�E֫/��s�]��3��!�,yƛ���>x'�Px�3Y�%F��8��=���ަ^�{UzeIA$>T�ya۠kC��)�񿴌`���h�]���:C�w��[l_�b�I+���V�!J���%p\PAy��N��(0�|�'�}C8����D:��f:��!���Z�V ������]Ɇ9��Ja�@�\ \\֭����\<P�\'3�&Xa.��{Y���,+I��w؅�@$ʋ�����<1����CсJ&�[,P��]̞de��(/���K�q}����5�h����3:א��/뼈{�{ߋ���m�L8���g�C�Ր^]5c#��Sxd�����
ڜ�UiIU��C��F;�S�h[��'����=$CZ�� �c��Ԃ>*+��7���u��Y*:68^�|��Ӂo,�Wgm9��bt���d@j?��E��l�3��b�c]��A��.�+&UL�],k�ӏ�,������3���{=�#�-�ю�8�ɜKD���pg2V"�#-vR�B0�I\�G���R��\�u��P7Vw�5���?�Fߐ_Z.]���b�ͱ�}	~N����5�ۇc��lx� ��556�����Ğ��T/�@]���JUZRː�	2��Vz
��(A �<��� ��ϖ�W�Jrw��.ʱ������W��!��ͩ�n�^�
W��v>�����Y"�e|����%^��0qM����ӥ#�o�$����jmy�q/'�Ö1ڇ_*!��y�Y:4be�Վ��-��;a�>ĸP�w�Ԇz<����z�k~U��q�W��}-7���RT+5�}�^��2۩���* ������#(^q����Z���GB�5�p.�+>xlH~�O3��α�i��{���C�E1�/���&E��ݒv�J
�x�!��7J8Jw��N�_�[_��].6D�6��-�↓+nG��JA|�f2^��=��.[8H���7�щ��1�J�>A��U;I�?̧%Cŷ��~VB��v{,mfP44���p[ĺ�"�Ӻ�\����,��\zҴֵ���LI�jFKh�X0s�5ˎn�]hn�B��R�7	"v��x&燪fT�B��3��[�Q�9�HI��l�(ݟ �����\E������G����c�"�6Dbf�.H�K'�~��T)*�>~�~�b�E\���lˎPRt��.�`��l:��*��}�xD�����J\<-Lcr3�ﱽ-\ڝX�A��"�,
����f��Hf>Nي<!:/Ǆ8� ,D[�٪��.��袼UvY�Np���U?Q�	�]&�/i������ط�S�3@�^%0;�N�C'Y z��Qo�u�'�d��{�s(��s��?��:�αKQL?��9R���g�X#Ȓ��^&v����J�~��d������A�y,��@X=N�E���:r�zJ=�S ~������rwe*��45�3X�m%lR�+(n��Z`�6[�E�p�<}΋��������R�����b��^)��%'Uغ��*W����]�G��)ς��(�@I�c�?�Y	S�v�R�E���k!�xU�@�]��\R�&@y!�+��=*QTj�?r&�O��H �_C�n�`G,��8\��w%]��3\c|k@z��^x��CކD`K�[ߚr�a��5��9�`�+/KU��-y{ H�;�'�,�W�LEE\�Y.����Is�r]���+�9���m��"����s��1'�~z�g��J15m�G�z#⺜���x}���wV��|)K�9l\lC8�!
�"��������D�~��r�F�׌ ��R0�~8��L�sD�v��ڴ�53U�%�s��
s(�K�y���?����]��8�n(i-M�`��r$$�/�S]KRĖ���-⨙v/ER�l��V��4o���j�jj��A3�h�)���l�G���fJR�2]Gkf�'�i��r��PϊN�`�>4��4�ս� ��ttcߍM��o�^"��d���
,��RHmE.t=/�vo��H�3$�q�M|�u�-Ö�i������Yn"(����f�x޲2����1E��� �t�v�S)c;�%/�"jm�
&'CVr@�4���a�4�s!���Up���Pӛ��F�׊PKƹ��!څ�]4	�F��v�g�揷�����LM�;(��^���zO�
�M�;9%����\v0 nEa�etpo�	ob���7<�����������_u
��ŭ�qL%�PxƘq�#�� �.,���Q�]ϡ4eTQv9��i�KK�]�4�u��1.������%�yY��I��5疝�Ɍ��X�!pY��M�u���Hm!����uy� 0��*��:���8��)0Bw�\l�"j�C8���S�+�����n�_ާ���9�<�QZ�-�u�;g�O|[3��Px�o�5������@4I�l���%����B~��:�~\ Z��څP�ø��ѐ��F�3�����kƦ>�-�Pø˿9�ލ3�O��WP{Xq{�Rá�%`"�~���@Ħ�il��`B0�8Y�T��Q�&���y[�KhY�+��ؼxǯھ鴾���=�M��~�n������]ai�oM�?�}��Ͷ?lr�X3�Q�b˯iJ98���$	��M�C�� ��_���1������8����΄��Ճ��xsTGh>��Ӣ�Lgx���}�)@<��~qZn��((�2�����U��#��x�1�	�ċń�*p��R}���Yٱ����\MH~�.paN����m�ٝWx� 
�B��q0�o��7!�%���В=$�<⒇˲�a�A˨M������a^��fS#��&�Ggkt
V�q���e۵��e4�����
��c'#p����jG`����k��.w�	�æ�$q���x�ڨ�	o�M�G�;�2��2�1oeC9D
��	��5��[A&ǑVJz�y����W@��7��i��'��`��<��ϙ�CL ��,��C�����S���9�� ���x��i({��q	�A����Up��7�$;S�7�b���ra%Vu���3�d8��R���%� ���r�Ou��|�}O�d�g�#���_a8b��ty�^���r�0v��;7nFK��r�%2��u}��4U8�j��y#d�P�x�k�z�D�)X�g�Πѣbg���&*�ż;(,��&	)�,
̃�v�6�Y���n����U����l�e�nQѦ�n�L(͑�X�`�6��Ȳ�P�4GZ�+;X�NHe/`��>DaM�<��"��7U5l��V�_�P�HxPH"i<9˕����O���@݀�2MIG­ԣhZo����B��5j�����>ϊ�u=#D�1J�I[]�Y�?��ͺ)�2i�zdmO�}<�]T�!��DݚNV�Pݭ�umJ'2��ɐ������D�IzU�M{���xE`�W�(fd�1�3^2S��[�#���yl��z�d}�a��`S�^Kuv�$}ҁٽq���B�&�cl?�t�D�(ּP.����J@��L��.ʳ'���ߍ��nN������&Q�&�<L��f4��S9��mD�>c�|����}h\��9�ӻ�I�h��j��!�hy=E�$��[ߙ0*·b2���L-���7�F�z��Dk�4b�{�3w[��U��Ȗ�-��	�0�#��L��M��ar�fv��Ձ2�\Yww���l�Q������ �+�Ǎ�Sy����Q��-���~,��#!�`�����yZ�[���ߑR㌴������5�W����ӳ�����(3u����}��M�絮E%G��W�w6ۦB�s��C�=��N55mF?��G��������l*�,0>���#Ǵì2�:�ϝ��v��5��e���J�bX����F8%�2�9��C�s�����y�R�0�1���|�k��y�/x��R\��_�fISK-_{FtY|df�&0�)��i�F��8ڀHJߟ���ö1�6w崫�,��6�Y���~��I�Z[v$E���b~�D˔��,<�$�F��"%?�9�`J�8S&�i���3a{�:y궡�(?�U�7��)V��H�:�x6~^GD�C��d�������>vpl�O�[��L�����zF�.
S���N�bޅGp� 6�=�
jO�x�8�r*�Oo��E�_��fXF����9vH���kX��O���[f� W-�z?Xv��[cS(w�u�-A!��� �����@��ÿ�>���.���QE�J�eytE�$]��)	�2<)�I�`m��e��Z���D��^`soY��V�'����L9���h;󿰭�ܡV �_�=q�ƨ"O��E��pʋ
�&�O?^��!7��K�]��ܞ>���W�4=rA�5h5��Q� �c�&x�Yt��nٕӣʆ4QL���@�W������iI���lk����o�Y�:���j!
V�΂s��L�a�8�*Ԯ�0M������S�_�n������Ro�a�Z�<�@��(ܼ�̬��Q/Kx��79�l�&T���ó.FV����W�XS˲S�#l���8~�*�du�i�T���A`��$}��(?�Zى����Gh���D�>��&�j�uʝ�T���,tRt��
�r*f@-���۵<���麫�O����X��������0Br��tr��ߝ�u��~/���ІrIE�,�5&��)�╎�ƀ��f�:Oj��C�7=�r�,�!lX���E6�v+�e��C^~�N�{.���lv8~��PhD�8T�J�S��x���qF�.
��ZQϚG���Ϣ��X[�ʮ���&��Te�i�ذ�~�
�
3
�*��kRd�s�_�Lǉ*K�b���d��K�w5�L��'L�~�?A��G2}�����I&Ě���scR�6r���I|�?8I�]#�2�6��u�\ ͂����/���8V���0|��. �M��3�)�����.�n��>J�Q}`�'&�-k�W���]zS�]S�K(������7�tjf7�Je���>�tB�N]Dɮ�ݬ��&���j�fO�ruQ�%�i��9jv��'S���¡�!��]��30�4����ݷ/Ui�~�B|�"$p6 L�����`�>�3?涿�E&���:�6�G
�.Q�� ����ϓm�6�j����]e鐴J���U��'Uj��� ���wa���2=�;_Ab�8�h�;d��qW�	@�؅���Xm(�G���/�ȵ��!��,*ܨBЀR�Œ\��:��l�����jv�G��$jޜ:Ry;��H��]�e�jCU�?���@	M�N��is�
e(�N��̙�ZS�+Q�:$
���׮���E˦��dc�5����K������>	dέo�b$��o�W�ErH����2�e���b�(�u6��#��]{Zq�p+d�r�eV�?a�?8m[��9��Bh��S8�j�f�4wR�:�"@Q��(�7�&��rY���y����о�/�����$b$8�u�r5�sE�y�#�D"&��Q��}�̣�WG��%�^�m�y_���|�Z&V8���PI������I$t�a�RU��7��En��4��2���jZ��cAG�3B����� ���\�p��������ltv��^���9�E���F -�R�a&�
��������#��AF)��SlH�د�c��Sʭ"i��*��8?�����Ү���W�a����;����_
'1n�F%�t�/s*}�F��c���jg.��ak,dW���Xr�P0��&�M�*�D�?�_�70w��8E�P��T����ې 9��Ǥ�,�nG�^=D�M�dJ��I�f��lC�l���Q���/��5R��v��-��FM���Sj����򤌌i?����
}�>G�\�\�;�EmOϛ/z�?�N]<i�\�u0Km�~D�Pʖ�U��dP�o���)�󬵯w(���eo�>�ww����SJ�|�%p�ս�ͳ�IL|]$��������������!i^�U��M+(��n����$�\��k���+����dR9���mi���DpV��_�g~�QoZ@,¹��aU\��
��';�ѕ�����)G��"������7��3dt\�S�����N6*�+���(
V���S�'� t^��Y���۔���=+�m�s�Գ�N7~�k	~Z�{p�lw�Wj
�sP6[�FǏ&���@R��F?��렱�;٣Y�&�������SO��6�C����_B��kD�ݖ�U��ٺ������ ��.� 5�g�-O�=ů��H@����33v�w255�*l�*�r̢�+`Bճ��H�䳐�.҆$�U�L�R��$�}�Ω�D��,�����d�ž<<���/2/�,��7���h���� }�O�Xb"|�6�U�c�;���H4yH�[K ��d��l�p�є�T�T��MMv�\ �rb��>o�op�����-[2i��. I{<g�v�ryγ�����HA|��<��0G4|�
�3��X.iW'0:�$V��!"�����3Ѵ�k�~.�B����7�u�𳦖� ��~!�@,6?��y	#�[g�y��)r�G}9{y:�d�����h.�fL��CdEH����IN2�g�V������%�� ���u�	�ƳS�ʚ����pn*��9@�����dTs8�L=ź4�p�s�scD����� �彳��q�!$�r�}�y�zj����ks��PClV�D}3����D���@@5��z�V�q:>x�cS֝c_��-c�\��u�/Jo%�1�#�^�c^ʄH�����̎�����1�/����l�a�C���#��$�\�#�}g��]�l+��<4;�^��D;]~#��ѥ-k
�?��l�h�i]�*�]"k�����]��4�0a��p9���Z�tB(�Ւ�$'�ۤ:�w�i�sHIT�bT�<���S*�k���{�N�����v@z��Db�Aw�o����i��L"����/�%���ʬT��s�D�l��B�|�f"�#�|��~�[F��ƹA2̐z��IF�����u5��sb�dܝ�~QZ�
gI�L��`���6����Gu׺ʝ��u�X����p��&�Q�6U���p����=�����9��=���u�K!B+��I_�t�������qv%5ڦT�>������V���H�9�t9�w���z4؉%�@�-��6��+�w����Ϗ�����Ua�/]ز��r�W:N#r�]Ed��U�;;��	�:[>�>fj'������c�:a.��-}����j��Z��3=H���uεN�(ع@�Sj�B`�Mhvu��#�6���/�y!FaP�ي~���\`�:���ҏ�@��	�'�`֪�}���䘣O�
,5Jd	۠�<��,;�"�fd@�f-� �4Db��м��Ԯ��d3͟~��L�4��˸E���K7���۱`%/�+�����\[�A�1�q-:��^��k�z��K�@uV#��q������X��s��ᠡ�"/�n���a�z�[�:�b�������j-��K���	�&�4­DZ��Ƿ�Otc"�I��P��pi��e�-@O�	ή^J��:R�����8}�Cё�g�U(�'��8�GIмl�(������D�R�?Dw�������mCg~��+ؙ�1m����q��jzE�S]���wwF�\?��e^�߶� R�!f��	��0��	������z���lV�Gi�pj�+����#3~W�t	�`l/��24B �u�p�]�f��x��<��0;�^A�C�l����Up×�,�(i�<��_^�;��^.�E�'&
�y���P�FZǌE@���rȬ�v�-0I�ʜ��cnM��+0Ʃ-@S�s�K�K+�{��ሗ�=Q?���i�� Z�q�$�%�̢�RƗBH���|o�-�A.~�a�x�C���E5��/�ǆưE��;�6Az?WEj��1���fe�2P�����p���o�`��q��Նޒ+銝9��"����bIg�\��F�e��^a���[�Q�[�@��Y� h�b�<9 ~V���=�O��IF��'b�R��')F�D&"�%a B�K��t:����氆^�u���e�]���(���,���Fl���4�}$��'���2��Q��o�9)�]5��(�!�*T&� �U6�"�1�﷙c�!�Vy�%r� �x�a�{T�W������/�%<O����	(�9&�B�Ug�f����T�j���/Xgs������'��v� T��u�5�^F�_kw~�����'�����	�2?��/���,B��(YU!6�[E�+6@B*S��� �2�U����+��0G ��f�FN��`ugM�i���/��l�R�K��/��|�s�~`ײKN�7��S�
9*�4���r�p��� (��>����/������t<&��ݭd���JH��f��d3G�f��Y��T�U~:{U㰀�
'����ژ��<�<�6��[o>�$��|�硰�ل���+��S����h�I5�3<7�.�}��|�x�M-��e�ʕH��e.��~FL)Q6��!�����jZ��P�E��\�{QȜ���J��)���� �@��4�_�ܓ��d%u����|+�y�[����74��E�h�\�1uD`��ü?��h�m�NL���fsq�͏��%[�����~�x ���W����u���m�4�����!P�n�%v����q��,0���"�f��t��3=#�P	Vg� 'ڲ��J�B��Ma�8{B*߮M3�:*Vi/_T�üR�^����q3��O�jwY��_iU?�j	���i"G3�b��o�bqT��� 
���-���H��l�o��"焏�����,*V4%�&.���O�=ݸ�c<c����e�.��9!̉R�C���d���.^�<(��`�H�$��^�&8��H�A_�Yg�dZ����K� /��:¸l�NhȅK@���#9�y�PƤ�޷�>Z͍v���\5�O0�T�5��Nv����.4�c�cPI�(�S����@+𷟉��"��)J� .�t�=�B���#v�����N��콅w�GC�R��[2'7f-���S����2��N"G���$$�����.p��y��y����g���,c���\)"UԦ+&��ʪ����:���D ���������\��NY��;��&r��s�~�n:.Lk0R�5�Z gv̦J�FO�1gT�%��@CZΟ;�����bT%|�ɒP�򮥵��o��ۉ��L�����Dg����F�K���NLҾ�D�1�6����I.;�?w����,�>j�k�/��/����۶p����D��#LRw��CR!�>Q�I!<�ٺ)���"	pð_K*�,y号5̇1,NA��|���HG<��J��7�����6Q!�Y]�����y��KØ�*I�l������SA3=dJ.�m��q�g�Ǣ��&�vL���`�i�)@}�(c�]�2OgäYŵ���L�a�
KN�3�|5G�o`J�dE�s�O���?N�-�1�,�����t��h�s��γ}�"��nC�I/��)S�>��.`�y513e�^��U4���(�I7�_|U��x�
E�^���2P��F�+��#�R������B�N�P��!����-̍��=
��V���/�;�tj.���.M��5MT_c�/ޥ��a:��(\hIBP�N-jrw5�4����c'Tv$C<�ͼײ	�����d�'�\�-�r�EPq�҈7��?o�=q����a���ժ��mm���^,
��C����Hp  �vc�-=~��B���jZ���f����-0��5S��@�MN\�*:�\ڭ!�j���n�q�[L*��AZW������g��<_q*\�ջޖg�\�ˣ��Mm��c�RL��qK8����x����A�d�v��ר|/9���H�����N�.�|�>\����GB��Y�o����b )&Lr�T%�u�Rg��?�m��_x�:�3��e�o�]��h�P�{2����Ɋ�T7���]����C����i�$��Y�3.�T��m�>M�����RxSP��ͽ�s�����~�#����ŪvFn3K�d��=���)�}�I�����0I�03X��X���x��!����FP1��#O�B)"`
q,q��o�k$ �Z��h	FRB`�g��@����f�hS���џb�l���g�$!��,?Cy��a#[h�I�˦���c`����ÿ����@x����Y�*�o��)��_#bޔ���9ܮ����x���ѓ�b��9��4M��פ�-��X�<#Xj���q��p���,T3@��"���%�0��ux����Ա(� �
7x�s]��l�ܢ����Iɝ���I%BH_f%\~��Iok���Z���q�)<栟��1Xo���cԧ�*�-
�%��U@�!0�Ѷ�t�ұ&u�I��Y3f�r��:2v3;?|L�x���=����8�9K�����V��Hԃ�� �{n1�� a��Y�f[+w�;�ea,4��|���!��Ó%��=J#g#�w47��=��J�֌�oh�E��s����pX0K�����A�2�ym��I�5�i1�.'�'+��4Ò0�`uo�0s�.A���A��%�x����XP�8�N;�O�R���f��C�<��0���]w�&��I�&P�.�C?��p�:���q9���MWӜ
��t���+�i͙�c!�1�^/S�:>g�dű����A
9�^ �Ch婄���o�5�N�?��G��gݚ޴glހN�K�'�qK��K��Yy��J)�d�����#��7+��]R��ʆ�~���F1�9l�.�ϫ��f ���1]2\z�49i'6��?�����6q\EAW#�ޜ+����
9�	p�l���߃Aܷ�>�>�$��?��K�^%�ǖd�h˜��4A�1���f�j�n,ٽXNYP>H�=l+${�n���X�d�)�2�+�j��+�Yҹ�Ձ4���ğc��a�I��ĉ�2�M��'g"!������?~��G��3T*�5�5*eި=�K"��=�]��8u��S�?.����2��w�1)wў�D.�Cy�d�{��F�6 ���:^��ʙ��'��� N��p��9'���!�����E2��# ��{l�E���se�V�R����_����>�DAA��a��$���P["_D_��,����!�]������zc�X5�<����u��L�ң�?8�I�%�/$�����D*�h�f0�n��	 1�h���Y��HIX*�ZbV�+�|vgHa����'���goX�?iv���o,>���H�t$���ձ	�Ʀ� �ꖡ�G;�n|�O��a8E�9�q�*��ł�O�3�$T2�K9�N�%�N�R��hA�/�M�P�0�Y�pX��z�Ӓ�PC�B��p��Y�I2lw� �h@�. �t>2��5s����c�Qߢt���M�|��ؽ���*��F2s1��{�p�	S* Ȁ����h�d95>�/���X�z�"��!/0|��̲�s�hI�:u�D�S��E�v��ȧ8�V������7����II�@8ge��I��h���8>L�Q̓?�*oe�컩㿝�=�:��JE��*� �Y�pʥUK��XgN�O�C�@��.������G|��'[������l7�i]�9��m��O	p��[^$�2=��q1�Hm"%�)k����CV�������+J�ó�7 Ȃ(�ET3�2�L��Y��dȆ��7~.�����"���C
���
#:j�)z_�Q�r>���A���f��g�eJD[4y�x#q	�$�l0�Ώ��K��S�Ӏ4��V~�36�	Ń��L�P��`�#��0��v@O �s{S�l��d��F�_���b���^�Q��t�n~�#Έ�&cno����0GYD�`��e(\�6�q�Rɽ`Ur�}���f��f�6.��i�يa �d��%���ڕ�N�Eά{@��[��v_F����{"��KO0��X��@$U�dS�,�\���+R9�p�@�OS6�B������0 �r��n$���l疘��	E�۝x|V��R)ʡxvsov�tE�x4�"s����>�T	��TΆq�DƟF-��D����I��SQ#3f���%��Һ�$���di�p̼ b�W��������m�K+y�u2�3S�H/	�B[�ru���7�ag�[1�|�B��Oj+�!Ϟ�),P�BN��T�����W�(���)�G�'�6�ዌu��<�}-ⳛ�A�����}��0mp���t�F�%r�C��3(�~��E[UT�@��7e�Ξ?ȍEp�.��'��c_|cG���'د�A��5>�5A�ە��z�}�gR/�% ���ͳ`��JCW�� �ݎo�~�FӯHt���3[��ҖO�^7u5��!Bh�anH>����,؄`	�n��Js<{+��60uq��.H0���C���=[��)=�=�LjBUL۝����u (jHhn�=g���Ɓ��x�$x`q���VK`p����T7��̧��yi��Y������!��z�΂'�DY�������x[lI+K�&��⡿�=!������Q��3�i��O�'��Gnf!Ӝ3�tb��q�@8��%�D�������z�_t��bD�/F!z��P�����z�͚R߳���țo����a2z�(mY`�Ҵ=�-�։v �c~�\V�W}V����6M�<�xk����������q
e/2/�n��tR���Amd�v��[Lm*-f�ʑIg�W;|FKM�˸lpmf�!Q0�j���(QW�=Q� �P�jc��(��c��7���Y�����VVZ-f\�ڤ]�f�����f��)���2�,LX��6ؾ��{�۱���`�% c���P}�>)��oT"e��,"�="�G��ň�z�����SȟIe���ʋ싓djmv�>xE�-�����HXc����7�I��h[ܑ�΄��#�o�Gc��¢'ɕ��𒷵(Ti���ʌ�t)�.�8�ʒ��\���Dm��j�Quisk��C���Żi��^���6f469�#�8=,���ϵ���Qx��b5���ȕGV��IV��u�aq���g30��Ϳd"$x>��B��u;�!Sf�݊k
�&4��!���mÎ'�������Xo0��7G��c%p����MBP���W}`�I�)�f���+DZ���C�=t��o� �5 2O"�rou�ה����%���A���u�n�J&��`���@X�2׫N��i��J\�'�2�7��I��T�/�e(ئ��W>�kF�**��t$A<Ϋ����)��'����Ȁ�����j[j1��7-~
k:���F���K�I>ijp��(3���G��߇*?�F�-[c��h���4�+��M���G��ǲ���t�H%���ܘ��A�:~~g�A���������zs#ɴ?����3��ii�0�}�:�����`7}��p�G�(�����7囆�Q� >�z�W	�
���1̀���S��Yv�iE�
���|��n�K2��8#��c����6�2�6��)��J������O��Z����8���~^��IXDV_��8Cuާ�[�f&�:�M)XF([h���Ҹ��qM_��A�)B?TU0j�9�c��K:'�͋����b'�r쎙�T{~ٚ�ؐ�7C���v�i}t�ze��I��]5L�H(48�C3m���d���,�x��6�S�	���?���C�"�nw$��,��&�v��U$T�!��n�N��.�C�U��&�����DAlN���}�<�2`��.>�N���~ w���^�p��_���6h'̌f�Ɩ��@[�8�9A�I]�riB~�����ɼ>qS @#֤��@sm�k�y�+ο�B ���.��W$K�H����xY��T⽡�ͤ0D|T�t��O����,�� 4�Y­�[V���R���]�_�ʹ�޸I�ح������_�Z��6�Q1�+���}��Z[[(\��8wꘄ�Js������a� �m�g����>����I�I+'��%�E�K�:'}�1�4��s1�
���������>x
�ݢ�en�ՠ`���*����8߉�����e<F�}u_��mz3��5k�u[��x�=�,A��5j��@���$�'�K�@L�����'*�5Y�J&.�a֏9�6p	N~t�<��6@8�23�q�EI�;
9ݥ�ῸT�M�'���1o�mU�/���B�oe}��>��D��e�/*��ЙD= �/�P���Ff�ٗ�����!��ìv;͎�̙�k�j�Q>s���N)=[䏑}�n<�'�S�t�@\���W����WW�Oct~��F�z#��x�c5�a����y?��F��H,~��2����"�@4�ؿ���&����Ǔ�Ni!�BA_�`��liR���Iv���a3wJ��+m�?��E�?�'� �MR���4NN���#p�<X��@�}7�9��lO'�ZQ
j��%�<ƶ���)������2n�|>sao��UJ@�=/�Z��.:kВ���e�7�n�l�?��"��yRiZ�sY�vqu��: a ����p�^1�g$Yƀ�wmp/�36>~Va%ۤ�ȧR��<����1�}�s!����&��8p�vw�lD�9����s���\��2�ف1��'�Z�s��v�W&I߂
B�>���!��؛�_b�b�b�[�O�s6ߚ+��fT��0Z����xA�w!��q�rV�f(�&�zZ2��e�^]�NE؆�l�\m�QHʟ��o:�=��Wɘ��f04v+c����*WWX�����mqۣ�BN}��dtҝ!Uab�®�N�#&�6�����zND��:�W5o.�;6%���NDv�ǟ�*|>�t�䈐=z?�O(� <M��C�/��N��Ģ��=�r3�*_�p&�qVp�(7�Tr����Oiv��fOөnU�\�2S��WprD��$p"Jp��$�}ǝ ��$S[��q+3��.�E���+�~�_>[fC�d�֭`,���jַ� �n�	�d���ym��Sh��|��� V�M�6\�zbes"�;|�a���_gߦ��3G�^29��,�7��$���\��s�e������Y&�.Um��~^?D v_T��:*�a#ʹax�>�eUʒ+�ȅM^���l��I�h*��m�-�4S=����QŖ���L���aNE&�]��iF�p\ ��qA|�Mk���C?j��5O�q곛宂o�ߤ����� �e�xOZI�A���Z�fĬ/H)E7d�/}����gŕ���D���>!A��~�ZAa��s��`f(&l�y��V�6@�4���-���#S�\��j�F~��	G߃r��!,�W���&˱Y�I���v�/�X��Ym��nS��>���W�D���i�/��iwj��B��mysz�:nrبy-��dN;1�8@�-�׬-'��.�p8�l\r�|#&���^��?���V�5�7�L�T臏zy����E�Ό�yV���ෆJ=����w��}D:���L7K�D+�v0�oDe��5������� �&�^\߬��\i���S����)���F_B�Z��.���X����>=�v}e�}����Js��z�;4��H�A�P.&�h
��<�'���yHhx�=��PA6�Sޮ�{yĚ��T�I�~?��$���-*���1\�_t��"�3����
+�����]-��ݻ�Y����Iѐk�:c,�=�9(
��$�3�GV����4Jk�����&��9E|02��a��µJ0�-�V&>'������a�(���	�7	=�F�I|{X\A�q��$�0�AQ(.�.ɀ9883��;Qp���e�g�ݶ%"w��2�8 W�J�yX'��8�Q\I+.GkqI��vۼ�H�V�:>Ku�@X��|�7JU�Z��	V'�r9}m1�_1��<��2�Ić� �O�Y���ע�8����[��:�J�6��&72L፽y��6�&��]�ihE`�G�Q��#����<��`�r[|��:*u�/�*�� ��[�B2�nF�f�<�:���{����ݲ���nxu�ql�=&��w^m�Cݒ���U��A�"]�P&�qR�fa�[u¾��#qY��n2HT�����9й���<͋su��	_�xZ�-�!�t���&�5��2l9�q$1�(l7���Ak߲'��n��ur��^��e��<
 �!3����Jf°��}a�o��]w���];H�� �{͖lI��r���b��^�wرÉ5A�M��u�%���(��鶮O�[p&�_��C�a���X��F��e߮C���&�{�&S�_�i?I��q��N�{�B@�Ii���F�������Y�0%�"�ykf���I1���[K<Ġ���VW�e����$u���J�[�#*�/>�3��đ*��b7�!k���ِ,��j+M�s-q?N��b�Z�1�4�Ӝ�1�4�` M��rb<r��{N�^�nn8�-��Ax�w��]�R�7�,�Y��:����@�	?H�O��W;Cԧ�oaJ2��U�0�����`��^:�\yJĠd�� �S���i��i@�O�m��%�&���Ģ�ʲ�L�"����O� �n@��.n�CU�L�cv��K������q�	Y}�a �~⨧T��L5��_A�.���-|���|P�a�󇢛+���L2������ՒP=G��>HJkqK��1���Y�n�S�E9�����TK�b�_���KzUG�7t�`���֔�n�ChPIAW��~6�g���.�Jgz�Ow��(M��!�W-���;LU�`�D|E�<iQ���7�.�/4JZ��t� �mY�P�CDV��Ӳ#(/Eެz-ٹJ���	�P�;P��i�6��mq��x�!��һ�C��?h0c�(c�0�Ѣm��^�Xt��?Q��I������P\�Ӧ���R��(>1v��ƒ�$�������u�$��vO��wB���2&�
 ���� �U�b�4	��~�ڻB(��U��M�'��֮���?�^�Gu��� ���JjHT�X��7����Y.�	"J�2�mc��)���;���=��c�̈���%2����r̦/��{�kUOQ���K:w{D�jL���4��g����y�d/�aAD�ͺu�첁�N��dG��H�>Q{gB�q�uV�e�'Xʯ�g]=�� �?D琣J�@�&�ҝ(YV������cW�a�	0��Q�k}%p�%z楞��C�9��A7�!@��_�[s�uP4�9��\*-F�)��Y�6�U��i�9���g�i��qu�g�c!����&��K� 'kӔR)t�TT���Df�2E�wM�T#<���;X���6.`^<�,<�;�uq�'D�phV5mW2��02�����F�����z�,�O�S��	L�.Y�|�/��@�,�!i��Hh�%
��\٨�!�,�rOh��,o�(�pt�S�'���d�_H4��d5�&�>?�@�mf�'.6�a���o�;G5�u:g=�[Epo�������a^�R�^wzMt���\�Ԛ�0@Y;�[;���*!]w2Wu�FQ�S���ſ����t�D�+�͂<�:��p��������k��s8^�?��"�q{��n�KF�,�ib����s �I�3�f�W==^���.e�\	2+�����ᢺ|V/�~�=��څ�t)-�8	���'x�n��HP�Vd*)��'�a����	��$�� ϙ`�w��� ����T�����Ar�[$U���e��{�G6�7�q�9��0�"��SEn��޺����7��B�m��`~ 4��*����7|?ʙ���:]~�����gT�eeSv�n�G��nz���~���s$�@��S��0��%\���g�xrq�����^|G�Zg��j���S6���(
�����rJ�Y��K�.������%ó��D��%䑗V�����*%A�$>;�%�'����N��A���IiV,Њ�j/)�����s?���|*�`�8�q�˴�L=�Ϯ�U�R�G�U�]�%W��p��v`՛���O
n���o�.�~�6���ô�ݷ/�;��]�)x�^��}��U��
��m6ZO� ��֟c(>ع���6F�d�%�3L��>��,�^0,:��Q���=v��^�J����W�1�ѣܨ��H����Ϯ�~�n@�����[y���"$�Qz~��6|��U6
�1�r��P��&�ܙd��-�WَSBf�����C6�$��z��i��SO�w\�7��!\�{�zaңV��娔t��`�{n5���M�u]&q�O����Q��q�x�i+�Ζ�4ۨ��Ӣ2Z�����]�a6XAf����,���D��Φ4B㈇R����k1�Ѽ���<Q���i�i�	!s�b�bW�7"B������?=���v�y-en���K)��w�m�3����cO8��j��aI{v�Ltr��>x�EU�E5S�AB�̈M-̌'xN����)�|E�D�xR�����~��X0���:!�/��[��J�-� ��G�+��cW�X��7�^�cz�˱�Q�A'�ɩ�\;؂&�.�:>�?6��4iz�N���~�L�\����c����|涥̭;��,Gwt�@uJl_�x�O�l�2��`�����s-�؝Fx���˽4��&6D\@f�(���T�x�/@��թX<�*�U�6�\?{�@|��Q�K@烦�#�^�Fv�
���p��4v_(n�&˞&�������~馲?Y��%�7u����DF��4f�]N'�]� �/Ӣ�����L�@�R��b+��
ٗ���;ړ��z�TݏZӀX41QΝ ���[�s7V�D-�f�c`Gm3���!���{iB��m��n�abK3�4�PM��g��P���z����`ΰ���9O�Z�#����,�q#��A�M����T�~/���]B�/)���*KK���v�u�v~:��'�x�l���ֹ��[�˼�7��⊝]R��b�@0�	�' rH�L����#�n��(��� �<�)�E�&&2�zQ�f��p9ސ:�d*J4��K	�u��"�V�1��&�����c]�p�""�ճ��T�QL{���M����=�j<l��aN���T���~nU#x]Q�6�ߝ����-\�LS�]�A��.���R�~��<�/�� �,�A6���v�JF��c%iLo��7����Yؠ��S��.h�*c�(v�����<f��e�e������E>3���v���(�|Z��F� �������^XY}!?5M�8�l��IY��䇞rQYPR8kc9����C�ա+V)���S�����0ѓ˝�.�����p6��80ϤO�SU1�%����M�Mz�L�l�@������"<�ϙ�Ň�3�nا��������cC��: J$�N��)���d~N �Yм����1��1h��!�Ҏ�ɷXLu�&��K��wf0mNV�U� �����Ʈ�E��e@�#^��lR{�$�J!Oz<�9���֖��iOC)ܰ�$t�5@@�Pq���zYC�Sg,c�J���v�%h�8" X�|_S���?�fi�Z���P�E>��S�Ωg�8��s���n��s�!v�j�.�`$�'U�:���@��#�޻Lnɼ¨�;����oj�����};�Im}�� >���ẟ����NI!:��dH���In|���]K,=�o��p\��ne��̢��Ii�Mllc|������If�~+=<(�R��$)IW[��<F��� � O5@�B�����{+y�����&����-��"t�٨v�k]���9۶�,�sm�E�k�?7G^�䛅����o���$,��%Q�T�K�v\��>��z�wk	*�=�L�z:J/�6�z���U�mV�����|	�3xuƈ�
M�a������IjI��+1+
,jB}c�;�1�����v�S9��#E�8�$��s �ԛ��ir�`�K���FY_��!��7.�4^y\f�j�#��{�	��g~\����s���M�.n��Xwm2��&0�x�IK�lL��gV���G�82����mؐ��"��A�`�w�-;\��d}A3��h;����Eou*��3��h����q,���[�Wi�"�B���9&��]�؁-���0]���4&*FdT%3/�vIYqr�%�9N�<�:(���:���5�%-waP�v6o����pm�'B�����nA٤abj}HΌ����.�9��Mh��>�.����j4Gjdn��w�\N���+���o+@	w�%p�Q��W8
%�4 FoBXü!^O6&:���{��4�ԕ:���h��A����x�x:�����������%C�JU,d.�������Y�:�z����f e�5�r�l�˧@y_�g�w�?����|��/��ZC�t�q�B�F8�Y[���状8C��;E"4��{C7����Y��U��b����ゞ%����Π�~�����	O��R�"x���E1CP��H�p�Y^K�+��{O���ˢi/�Hc�M����t��t���,�p���$�ގA�k����U�)�A؜ �d�$�z������u�?�g��t�0 �1�Op
�~\э�J�$�s#��uo�H>�=�43�����Rσ\��H���[ߛb	���8��"<N��� z��r6LH!����b��)%������M��>׍5B(����S��C_��o'o��6������AR(�tc�T�1����`�oɈh�NJE����P�ߐ*�V��3��ŭ{�VB�_��=�8�b��yk^q�c����O�ĽQ�jA	kH�#9�����B1��>�Q�v$)��0�TO��ǫ/��^�W��6I���@o]v{��ⅻ�')��� d4��R�S��tYrpx�G���hH&j�	�t��-c�+�n���P���Ƹ9�8_�/���JĜ|����M�{�ݐ�&\S;�Z$�̧a�f<g V3(�P��0��k<nP�ڝ�t�Z��K9a�W�K��"�68���Ih�uyk��3��B�-���o�w��w���3v��v��ִt^!�Ö�2*N]��߭�Q-��=����Ϸ`%�J'�O�����6Q=`�Ѯa@�C���`�6A� �����G��>Ѷ[r.��s��9҃����7ȍ��>cٵ]�m��A�iS�@���'��Vh^1�_��d&q���F��Y�������}~��p������Ek���5~�W�'ZG��t����#�댭MBk�׸o ;��9~��M�<.�A�azӮk��ԁ��K����CQ��XJn�Z��F-8��R�`%�C�E^q3k���ܟ�Jf9�����0i���jm>��e�/�[��x+�ж��%������v�`M�O�)�u{���[�'�'M�G�f]q���X;���W�u0�W�_��΂$���6N����$�d�k(+�]&T	�;���(��$���)��Mó("�i,��5��]'�t'��
�R���G�{��ޮ"[��@%s��x�0�Ï���\1�Re�)*��q�T/���IE6i�[�_X0 WB%Á��C� �WP$�|�_�
��17=H:-Ry5�0����F�]��Fm��G$����G�����A�.(��ڗ0i�.����/�ּ�u��������ߣ����J�6%C��O<,�AI�k��Y5E��g�sT���Ęg�9Qp^m�mGL��ۢ�I�-J��3�]�/���V(����~��({�Qp�Tk����j���'�gл���S�U�=� ���2@q��*%S[��Xy�T[��{['r͟��li�jU�I3�vhk���O��<S�	�jBҳd�|�/��g���	����r�V���W�a�δu*%u5�ת����gړ���
bI�*����K|��Ell�M\�9��Y1��@�W+Lp�;KXm�W���}�*(�=tTҫ�����1�����!)5H)D7Q��g�A?!T�C��}�����0-�	5Z�w,�?; �_����2�s�"�6k�a�.�h�_�>�4L`Ȼ��I�P%jxtT`Ϧv�l�֨����ϲ{����b)��'���*u��{S�'�|mL*�Ȯ���0��b������9G�c�S�\�`=p���q|����j�354�Q䍪�^�j�kn�'g�o���?�M��t��x4�u���6VB������f�G��WDzK���r<f��j��Ÿ�[O���2T��#�F�U������2�x�{�%s��9C�[j�Z�ۨ��)�l%Л�qւ #�H��5�����m	��s��"v���((����ȏ�7E�2z>�(�пt���.�]�>�$��,�v�i���"������W�ON�)$�kG��6��܏w���(N� ��;~��r�l���/����\�P[L�d{l��!��A����<�Q�A����R���1������
�����c��9q���r���t ��i@���5�%����XX�m���ǜ�F��}��Ơ=�w7V4_soGhf��؀�� j�� �Y���td��a׍�8��\g����!b_4ͷع������{IC*�ԡ\��W��B���Gh��7��y�ԝ�`� ϞЕs�/*l'b˷[D�Uc�:=
��@70�-���ϝ]f�l�9=�	�)�e�8W�![?��%��iw��SC��	H�(s�{�^A��_(��V�Vu��h+0l+\���Kv�����>������ϩ�6qal:��F��\�9��2��ۺe����Y�N��N߀*�$��o�n���i�`���h�i}�]�57���$����{O�K��?���i\�n�j1/l��i[K���c�0W����<sGT	� 얦��MZ�+9�÷fCY���D~\9�UX��RK�=���v��>�^K�ȓ'�H�y��p3�nON�Lw$�\@P�?Lk��H���ϻY+TuU������Һ���rr���:S���DB��n�AV�S��񛣠rÚds/jj���v�g�$Hi���f'�8+>Eڊ���nҡ��u�����O"��di�������"e�.�g��m�'%NOzBjp�H$?�~��}БRyX��P�%j�Ta"²V����`��68Rp6�ُ&�c����R�R�!ʉ�7L��eA&�����IC��A@ݵZ�����I%�!�SȠH]�&�v�4�8yG�Y��9��������o�w�����#���ˆ�U��Y���Hů9 -��&y�ހ�@�;�0L�R-H��ʻdY�0��.�(�b��� `���[B�M,M~�'V�op������3��
K1����$9 t�������F�]�<T�\3}}^#f�>�E%�r��͎�6���S�7�]I�Q��u�R���Q����"��d����®䑶<6+�#m�.��`#yc��E9ї±�JU�Q5�E������8-��C�VO��>:VTN+y%
�ex�����uCm8+ot���	��*(���l7��=����T��aO����^����(D���@;g�#v�|j\��P �$.���/A��`ʡzb��A,Ɯ�U���eub?e��uT�wR�%��?ln՚��/X��Q� ��.�|�qU6&�bZ��l��=����;��pG��|>�o�w8���=d�bKc�JEٟ��Q��1�k1c�áq���umҷ���ep����%�kn�"U��p#���R�Q��v�vH�fhF5�;�������9��b�@چ�4�����/ԝ� ������vp�����ㅡ�S�&��X���N�}�gg���!�Ֆ��}������~ɱ�9�#��D���:�-�H��W^(�e'~O$'��j�����ʋkD�"��z.��U��O�8�1)�V�
;E��DtX"��Z@(�]hǹȶ�OWx�+I���n��ik�b����ҕ�G���i�U����ނ" ���5���u�K䦗�$���!�
6:����_Y�9OD��"ƋM�*���{C1.�)�4#��}.Q�Up@8!��(�!�2g���.���?�R�ֲl\#�K�Yz�}���YZ���~-B�=`��	K�����N�vV�G�t|��/%�v��mC;m�3;��?*��5��]�P��tߣ&�z����M����U�D'��FE�0�<q��|4�G��iӸݓ MURJ����Z�. ��4#n���������"pE���v�3��t����ScSqr���~���ao���kýCv�O�A5�c��F`x�������D�Y�%)��.�<�`�L��@�����aSKg^7ѷ�ed�������K�x͡y����yT�����P�ߞ��	r7���T=�fNw��Ά�.���Ԣ_�����%���x-ݎGq �m qf��h{��O�'aڤI.
PU��yS�L���{S��o[�PZ�*o�/�m��}�h�4�<{Hz!u���܁ҬxrE�p=��}�?��Ꮱ��^f��H�n��I���W�>)f���L�-
&��̘%�F� ��/��v鉡��w����kR�ϊɆBE�-j�;��s���,���|f ~��_	x�1 ��g�O�X�[����A
P]�+��pT�S�%�_���e�9���PR�?�?����0��.$܍�*6� �\�@!�Q�6�v�K�_�ŉ �6����ⵍ#�js`U���ň^����Fa���x!��H�T�:�Ƙﾒ(���6-f>k`�:#���Q6?�V����ĩ!f�/�[��5xң���^\��Q��s�>0��Tw`kZ��Ls֒ؗ��W�H�B�h�)J\Oaߪb�<�xk������tm~H��Q;�Vt�"%*$c���L;�:�5=z��%�u�LuI��R�T63�Ђ#4Z?&b��*�I$ե�ꏽ�b�T�mx�g*��:ԧ>�D�r��j�[�ҕ��!"�D���VB�O�֦x�:� �}$c�w����Y����� ���#��r�O���P�'s凘[�Ԝ����;-a�1kؿ]�q
4��IP_0�]�+���|���558���%^>��Ҫ�t�6Sg^!�L��C3(�ќ��ٲ��^f�U4sh�#}$&+���L�X��O�֥��^�q���Rx|<��M�<7@r�ǂ_�li�j�۴*kH�L8CS�� ���q5���d�0�ô�h˵D�3�ts��q�SP�W������M>�@Ѫӝ���� ��p`�'�Lގ�3��f�������`ư�u~
��rv��Tf�<2��v! ZK�!R$¦1|n��%�o���7���.tD4Mo?����/� �Y�v�e�[�.�<2���lF�p�`ͻR`S�A^dr=��-V�{�5����Tl�Z�,C��?9��QY�_)���;�&��-�L��A���3Tg]D�sF؆zA�	��8��7��t����r�g��H�Q�J�����F���|��3`c�T������U�O�BQͅ���Y�)m ]�m��-J_�No��ݣ���{*Z�	NS�)�}4ۄ�s��ǈ�P���^K=����jP-�NB+��K�{~ ,���v�UM<���(�#����}�bD �����mB-wM�w���J����K6���;Q�+&����^y��a"a��@^;�q#���.b���R��A�-J���j��	�E.�>�傻$�,[k?��X_�c�V��򁢔�����h5�u�߻2H� {������UBXU����[yF� Ss���`�L�k����!�Z_�T9 y��^ۤ|����V䤏mU��ٸh!�� ^����l�-�"��H�����-�>ko]�Ø���,�Vć��P9?;�,{;�E��F�<Le`U@�2�YΩ�;������D��壻Kr_��`�6�*�B!�*�+�>Q'��Tkg2ˎ�≓#�(�s5���%��׍�s�1KI��Q��=[�789�.Ql2t��c���5����Iלn���j�S�'=z���W`�.[�lE��?[�Ȣ:���1S�8Y}��ƫo��M�(N>c(/۠���o/P�}��)��$ۜ�Y[���! ~m�*%�g���&�}�}����Hn��M0��^"���,}b.�Px=���}���!�&�V�_��i�U|�ddy��?
�T��^���t�1t8���CB0_�x$ѮY�,
[t��M�Sk�P�Tf%	�K�e4]}�S%��ؘ<����_^�:-���B���˅��)^>���~���������>��<�q�>����YU � �2[G	�q:��%Q��U�9 x�ձR��ex�^K�&��9�l����-|� Á��ߕ�m$m$���=��, VOL�޽Xb�lr�M^.�/�[�W���I���Upr��:V�{"1:�|�˃�8j�����~%\i�����\��	j�Z�UF^a��0'��"ח�@��ǧ���zmK�a�9�4�ڋ �$�
YwbK������$}W�5X�u�)���ic����v�H�Sj��Ѵ�=���,	74GU	;I[I6����B ����~�!��H�YyQ�I_�����iB%�����}T��7��w�bMs���:$���S��崫 	�dLy�Oƣ~�OUM��D�$��3��;�&Y�8�5��`�6z�.�eM��εЫM=��V���w��;��M/A������b�zBKc����
�0�g1I4]q�V�8�޻�I�n3��2��B�N�B�˼�@fВ��?��c�k���8?���1���\v׎�Q�]!���:�HG��홮xX���~�u�ˤL;��o�ⶮ���g���T�F�_�m �6-$:i���
T�$�B[F�b�8�*����Q�qvU)�)���c7��<H�'�&���{]��{(����7a>���W�H)���9��/
,�˴`�fY�4�d�4ɖ�VR&C�G15r��v��B�3Q���!��>��$p�Q~��^���G��1${��-T�$0��~P�Or���0�.��)L[6Ze�i9�,���<Q�"�q�Sq`\˻D��sU�Nj�o��np��b���4��"���6x��=ݒ�~C2��o�%�S=#b��B�x��vj�"����p_#)��Mhm���b#_�C���t�s\V��]��P�v�8�ye'[����C2#Rw&��
~��4�w-��y
�7-:/��d�R>��K��XgIf���s9>)|,v����$c�2�X��Z9�AY�5�͘8�@-Z��P�y��8N��Q��.���
�d���W�p$Xh�� m	#��C-����p���j#7&�Ak���=�wj�-^���H?5F]�<#�||>k�#E�P�/te��I��m>Q7��}�T�n_��!�e�p^6��.3L����1�63_U(B��;�4u",��/�*��c;��aI/��DA�}ZmɧDY�*�XXR�qrW��Kf�~y8�QS�9�ozd"���i�t篰^@��Jn7M���dy��rb-Gd~Lb��@��M]��sI9-q�.��;Щ�i,��9���uaiק�ގ��Q����g��;<���0ikPR��v�������9���櫽*�T�����8���[��E�v��7ާ�9=�I���*��g�u�+��&�ښ���G���Jo؛88�ɒ��g�q���T�����NR �e��;�̂=���m�.���Ml?~N����F4aZDh�m'D���`�f�O���)�i��۬���q7Z��'�T���	��B�;�8���sý8'��	@�fhH�>|�����Ϋ5ktyÇ>ao����3�zƘ<��/(�Ev�
O��O9Y3h�O(��xq#B���c���'E�Fc�O�xQ>�^l$�̊�JE�L1{��鞽5d������ozݐ<g1�*{f��|c�*EXgF�7>���j$�g�����>����$�*�����4Qk۝4)Iش������(3��!���?�8vp�v�sp��6e0���K�nn�_��_A߮2���KoǟPu�E)�B�tt	d��������B�(*�����g�`�Zz6հ���`�Wi��M�M|\�����ήZˌ��X��_|��iȕ~H��]�ܒ��U/�/)V��Z�-����D��@�����>UB4��ћ%a7������˴G1�r>R�ʤ��t=Q3g��m���X%����z�)���p]��gs�b�f��|�~FQ��R�,o�*�!���6Q��wl�G�#���o��k\�������m��d�I�Kb�a�j�n7
�`I��́$Z�����P,��Fe$<Y�*��43IQ?�{|�sJ@^�be�#~��w���x�T��{���)h)���;��c�4м�(����4=���E㽀y��b:���S^��
��S���R�j�Wo�i���1q{,g5�3dk�j�p�+�>@�-t�ju��&[ֹ�Zۍ�j��=8SB�P��i�W��v�L�a5'�K4�?�C+&^ר9�'�:�.c�.���	��%�]T���
۳�@��Vǡ�g����CUC���F�=r��[a4bM�+	%<�g�r��_|���G(�W���<���G���LCs	�Ј��FS�7y��o�I}r��a�߭�6������S܂3�`y+�w��Įn�/
�����8*�O���{����ϜK���6�)Y�����|x���퀲�;4A[D�ƪ
�s�/��?Љ l�4��^�����kۑ ��S��sW �ƪ?b�˦�Ip�j����=?�O�ʰ
����SC�iȐ� */ѫ�Ұߞ����#,*�W+^Bf�!zz��K"�V����}b�\;K�8V��e$n���(��=$a�
Ʈ�a�}p6���9�6s��j��vTH��C�(���juN�&p^�2�C3�CK��0�󅢤6��N?i�#/�1K$h�]�C��w��GE���Be;��׋#(˷#�J��S(^���)R�zUt�0/��9,�m��,�˧�����67*~���x�=�:Vh�տ���J:��4��t�/`LF�^ְ�:[�F8;��fn5�s2�s�g�J�����9`�݂	HƗߵ�z
}�1V��lQ�6j.����dr� �o���f����6٨*��B��zcFh�����I�#}��*�E�n�f�Cc��;%v{nT�Gps;�G�	!Վ����ߒ��1[��x������-#j�;����R+����y��t��D[�1⸏?�l������@����;�c�����kɦ�[��1��3���ʗ�B}�̷���Jܵ�Z-��x�<��P'��#Y0�T���,0�dp
�Њ�[�����lVX*��<G�6�Pd�A��+:XN�V6��� ���HK�a���4������z�fm��0U�35%|
��g���Dȵ%]=� e�Ȏ<G��|ܠ��@������f�zV���H��c�isQv'����NTd�f�CR%����P�m�4�_i�k�<qd*Ù�\-wQ�4M�d��wf�Rx%>J��t�Nb�������\欖�Θ�h��[�P�^L�~�J�j!�1_io]��o���B!�jpS@�a4�V�ƍDo�!g)h��+F*#�S�?I���C�`ں��e?Vז�-���.����0�X�>��$�:�
��������U�z����I0G��XZ`"t:3{O��-��¹Sڷ������P��i���� }W��"��VB�8��֜I�g�g��O�d��"6�[�%A~:&`�c#S�=N�/<��X��>�⛔6�K�-Ų���K6eA{^���.§c����P4���͕#}��1�Md��1�̱a4���W+��kn�=|G��P4��˧^kmJ�؃���w��n=`:q&�t�<5�nIE,�.I�i��^�/�o�QY�[Y���k�����aV���W�-Ś�_@���?^}��WPXV�`�g������m��n1�6�%D# l2z���fZx��
$�\�[)�1α��&�ΎPD
i��lt/T�Pϡ�Ӊ������3��*�l�\J(�8R�����l�՝���xKۤ�B!g�Hj����;��e���ѡ'uC�n�3Q���X^
��^Y]Y��WUôM�����%�h�gOpD5�8C��X�T"\{�ۇV�Z&o�����ēB]�(�偶+H�7r~3�'FO�V� ���yBu��6�B�nJj��@���G���]^�6�K����I�zZ�D!}�����!��ĸ�td>�dZ���FI1�������z�G��S ����ׇ��'}��Ul���w_�J�-0y��̅Se���H��YӘ����C\���:w+X�L�Q���ۇ�02C[����	K���7ÈR;vtY�]��~��*P}��S�k��T�\�lC"郠�����hشt�ž�����Y�B*ʴz@9�v�te�"���p�}�F�>�t��I�)�$�z�"C.`,? +��ͮ�eQ�2�刘�Q�J�`���8��E�J����D���Eޒ�� ��.�Ťr�*�$j��]ª�s7�������Mx/��^@��s?��L�[b=�s���?o�ߓC�q|y��ԇ|�.�m�Z�������d�Х4<��'ϪE7�P O0�lu]��$�e-�ƫo2����x�R-�?2�Rv3RS����ۈJ����$�I�Y���|껚�+�،��T���WX��aP�^�m��=߼�K2�ƶ"�Y�lr��G"`�ƕ+o����6'<��x(�]��uL|�� �X��W�M�R�y������}����<s�ыH{8�Wq�����v��~N�����]TJM4��hwD�����)����'7.'A� ��3wd�(��1O���\�'k'M��&<�e�?�
��'ZL5���o��[���N��jJ���og����dː���_6%&����7Rwc�2��"��z0��:^�@�����@�n6�U �:3*2���ᇏ\t�k/ʹ1���?auY[����pÊ_L�+[���WVp�%|�������[ �B�.�wqf��LBE��:����[�ιD�����Ҏ�B�{.��n.洐�����~�3K��/�#�=�֮:�$#���]�Y�����$�&�&�1G͆��7�K%��!i7HF"V�-Xg��7�ٴ�ҙe��� q�~Q�[�TzV}cG��6#Ε���ങ;0�>�M��J���: !^\7-�
?�*I��&)ʵ��z[����b�("�3v9�C��g,z0��?��[�C�ζ�x���+`D/�NJ�����P�l
j�h>8�̌�,�B��LD����DX�2��O^��i�؍D�Z`�4�֑���`7��ŵ������Yq(\Y�V��GB�����h��E�yƝ�k�|"<��1�1�#x���L��4KU�f��Š~Q����~�W�1�z ��X; ^p�(R����F��Ґu��c��p���	�aֿб_Q[���d��J`e�?�zhft���o�]�5�q�1@d�Ն�c*B;&�	E{T���렓{\�N<^�f�X����/�4lbO��#M�]�Q�����4ɾb�������wۋ6�-��4����Ci��H{�� ��h�-��6�˽1�q�ɖ���&<�-U��u���	��Iv� �@����>N�ۻ��Y�����zk|Ȯp��U��X#@��|y�.���&7�]Ǟ�����Թv�b���2�]\��j�$�1��)�§�}�����?�*$�>��ŀ����=�K��n���Ӵy�E'񼵙��F.ؐ6�8���W�Ӈ�3&�?�uW1�P�o\E,�d�̤��1��|�2hm��4Q���J�x��O�'ʵ�h��;9ɔdc�O=�z0%͹G7	�v����&�8���IP�_��Sa׿1Yy��"��pz����	��l����0�7���!GT������D�P����cz��?e��)�>�E SXjڲn6J�k�O}�	���tGr��������m����_��|V|{�d�3����γ��:4�gt֜���e�g��1��+1���F�	~x���Ei�[�R�Z���f����!�Gv�V�`�,8��^��q�6�p@��1w�3�b�0��u���ac�$�J)J�=�[�]uT��{���a{����[�K|./n`v�#���s͂���Ua�1��<�h��<��	c�p��͟\�(��".�T�m�T�4$/u-��(�N�n7y�Z/���?E5��Ѐ��^�݀���|��Y�ϓ�S.M{�
Y�2�~��e�Z�����S�s�~���٪Tv��z�.��hR*��S�<�|��g.X��m�0"7ѿ(�+�f5��:�Z��4C��'���d��O<� ��W�Us�T�t��ۓ3uh!D��S�����,�Ft�w�QW�<�Jș�Ӓ������Z �0�����w�z�#����X�9��i�kZ1sS>�o/����	�ro�v����92K���4ћ�ghQ��x]���XTc%x��/� 'KRF���k�ė&Jkd��P~��w���˥er�_��q���'���gV�vm+�uԶ���3���N�>A��so�{:߆
}/�H��Ưn:v��>���"�+�Zc�����=��&7*`��"�^�	N��ʭ�Ȯ��K�I���$�xkY���e�5n-83�BlJ�#x��m<	�ٓM&�^4�]l�9T��3�[Bg�i��{ˀ����@�ĵo+(�C���n�W%+O�y����B "��.�H���?�(������]#��;�m��@��7^{.��Y��|�zc?�M�� �:���'��h#��nķJ~�hc�����Y*(Kndd���g�����oCtX�㉨��|�`�E����-l�V&~(�-`���e �	�{�}�X����7����!~BELK��-ӟ�T��p1P,�����-�T#Џ���Y�t=���dȩ�,��vJ�R�ꙣ�R����4�4)T�pV3�91�D�
 @+�T=
��o5[�V�s�KcR� �&���kf:c���u"0Y,4�4��AO:C�1z��F�0Af.eu����� �����$2qI$��RVUg�kU�7��f�i�_=�8W��l�P;�~��3�?��m��ɏ���Miĕ�T@[B'��h��s! �,��s�q�;@pd�ƖM6������f��;����ń��2��u��l�>�R�7�%��v�}$>)Z�36RP:�D�����y��|'M��>	}����~��X�\rAG�I�0��/U^�t�ۀ��7V3�,�'�7p,����4b0�"~�黰�]<�J�����wZA�w��D����#�Nkg�l|�%�tD�<�A^�}��& �e�1]�l7vom���M���S�R	G���<�]OT'���m\��PMx�u���!��W}B��E|6��<ZhdE�	�L��Ք��NF�JN�ݒ]�g��A�"@Ñ��LC�����I�� '��ao��a��t/�}C�J���߬�����/B+��M^n-������()���$< b�vY=g��
����A#A>�X(#�Kq�}l�#6�JMW�L�<>󁵄��AЫ��'�Q	�����ʥ���n#c4$X+h�]pTf ��{-0�W^�٦�1ɥ�M��|v��"�j�����z�<�ӿZ
r�=�Zz:����S�����M���3�h����9�i	��a�Ց8�����P�¹��c��tB�zŁ��pT�%#\�3��H���YBog'a=�Z�SG��532�k��F�CH��U�l-CE ��E�.a�Ǩ��,�X�����A�lSQ�ȃeǽ�(�/��/��hn�������|�T<����]:�뿕G�� +��Kx4է.
9��������Ig5I�WŦq�ӵ*в�9���^��i��lII�:�r�]�q��L��������"�Z�x�Ӧ�z�ĭƞ�(��J�^��������%�JlV@U����&C�o�FPa�~���y�����)@���ҧ��'_Nm�&8����k!����}�3�f�Yz�m[���b���J���u|�I�N��r�p���/�H^|Q�����H&o��$S��EU��}}�-o@X��Op�$��\�,��#��pA�����a��&�JSI�NT
�O%>���g�F��@UT��`�L� �<�95&�D(�_2�c9@M�H�g��[fB?5e̥3�+םW��i��N6�U�����#��G8��3�~�^�ej�¹���?�9���0��{�3������C�f�K��H ���lN:�w�ŶQ�~�����@Ė�:�!:�ͭg���ŵ��ϛ��<��W8Q)2E��G�w��B����P��x�AT�t�æ����޳�RV	�R1`��TG�8
Z ���.2�cВ\����)uCr�-�'(���N^^�9 �G��$�d����jW*�I||�nE��C=��Iƫ�g~"<	���}5&��dP`q�'!__������)kci�TZ3��l\�x��2�fb~����������e}�Z/F�\���z���/�+�p�� <7�,@OI�d�l��p��zgL`�vn}u����X�#M��=B���#�����@zH��L��T9b��&P���_��R�tk����H+ܪu'��)`.g$�h��vܨ���z5-���}��� �b��u�ׁ��̊;6#�ٌ&,κ@�V�k�'l��;�u\y��ߦh5<b��e���Յ+L�.�a�S?=��9�����[�v�L�h;U8�%e��S�Nڧ�=�����.	�L�\�ˋ}�G��.F��w���P��?71�Im�$A�z�A�X�Ys7�A���`O/�-t��4�l��%Q%0��d1.�3��g�L�ϲ*�FD4���,��Y����]�1�-��/WS�����b��Nz������2z	Wۉ�r�Ɩ0oq�ye����~M���F�TPG�]m	C�Q/@���]ξ��#�ZQ��_����A�!Ӕ�b�:�,�?��?�>#�`��uE_ܒ����G�leHUm�{��lv�DX�w���y�6�S�M�vR�m<�t�Qb�q��L��@�%��Y�dP�˒�f����6�b�&�� �g��:�>^�xQ�FЋ�ev+A��9-��o)�-^j_NpX#|�;յ����p	���e��=���2��LS8nSȻs �^=M�ko�Q}E�$�r��o=�-Ec� �W	�����VS��U�͔)I��t�f,0����n�Ks� ���I�me����6�3���t��������l�'J��k6���Y'�#���5����uY��$3z�tp���s:���j�]�+|9���B8*:J�Σx7�\�"W��m��s��������茳P�,��4��0����(L��o%B��4R�+���'eFc��������w4D�.���5v��P��@�R�im�V(s����y"B"]���9��Ꙑ�r~Qz��O5|/�2��~�3=d5�8�+�xf8E8��^Jզ����/]�ҋ�yn�"�\���=\�`�,�-�L�)+}�NҊ�ܬ�ـM��}/�6Oo���wn��H�q���m�Oܮ��� ���C�+zE�%��*���G�h�,fɑ* N �@����-�~ܺ���Z�t����J�2N�໒~W�l(q-��f4i��s\N��PF�D3	���"��<��#�O�MM�q^�too=�A�hX�Z>�FExs��{��MA���y��J�԰i�;�pMir�Zٖ�X���w.�ﺅ�^Q�DB��Ȉ�ZlU��||�6������'������2P3���<,��)Ee|�2�I�:%�D�UOo%.�7���+��r|'��PR[]&�$]���ȡ���&6��QD�@=՛^ۗy�!�p�6�PЧ�	��r=H���`�\k<*8gnc*�qDW�d�k���������-q�gݻ�V1�;@8�{���L#鯁EC� ��#OB�T�^�K�����ԟ8�W:��R�7'����Y�u��.��̳�����n[N�b����Fj�:Z����:��pUmD Ll*�ذ1�{�;�M �q������}:��I���ԅ��3ã�'���&��� ��j��v�sA2����LֲeC��A9���7��v�x̏νQ��Q�F�ͫ� ����/���#(?A5֋s�s��k���� [�ߵ�Y,��1���t�[�	<4�l�%���q�>�U��{����]ķ�X����1Eȝ<0k�G�"}k�{V��̥�ĮC�#�j�Ƿ^��d��1Vx�`�F�����.TG�"�PZ$2�8���Ӱ��t� [̹�gr�N>��r��(�0F�������%zAAVi۶�y�Ҩ�3����˼ds/?soe�[���+{�]\�'�S�00Y[�6�?)��ܪ[�Or�b��v��h�gn�z#�)�HG�a��A�4�̅&+�r����K�ݻ9Q�К9>v$hKO*�}@1K��s��g,�ǵ)�Ӆĭ��~[�P߲u,�7i��0�^����z�w����׆	I.3���n|�q�%���:)(��������aP%G&�%$��� ۍ�I��5X���a������VJݙ'�_Pio�����R���'L�˸��B5X�R55Ě��B
$�cE�aDON_�?�O����s��D�I�n�˄F]����WnȦ�Z�Ґ���Z7m:�f�xӨ�@�|�i�:�����<29!�Rlt3��H�cOv����E¤bI����rQg[��iw
��UF̕�8�h!�����5с̥BA,T�� ��%��(������?�T�a���٣7N�����p@�)��<��� �<Ål���$8�F�! (����{_|���J {��w*k.�A ~�IԖ6��8Y���=�y��DB{�VyE�R�#;��H7<�U5�v�;��_�noāS|XV��œ�5���F�;Śd�5�>��|���k��.n�
GƄ����R��d�`�Lg��,-'>��s��zA��� y���7�m=��#���Mo�A�&M��dz��� ��ቢ�o@���8���#��R�b��b����������ن"�`����@e˩f|�T�ڒ7n��iL��	��D��㥧�}��#�u����ۓ�Y��-Q-��^��	b?�U�ˈ�M�G;S��F�ѱ;��=Gg_�� ��7�M0\��K����Y�ȈD^���SH�ka��̀���b�%g�d@y����z�u��t�a��Dǳ��
�SM��M�g�h���G�ƩX�麻�+�h����5�%����7V*B�V��<0�3�S�-[�	���ϣ��䤭�ܪ~+����ėJ�-�?��v8b]�~��Q�h�+��^��!��r����P�W��:HAp��'��\&L���\P�E=j�����=���?��\
���)�u��uW"{�z�r%t�U�=k���*��+�c�wc�CJ�?���@/	)�������6*�!첏{3�a�,���,��.^�
8< ��"�I�n�'I=�_����W�7����l�C{!�/b�g��+[�Uj^ l�^Ԃq�Mj�(#��3;�F��>esV\J,�1���Ӈ8���}M�p��\�$��b2f`@%��!o���[QW�.@��N��q�A䑂�#�/��+�c
��*�W��|����m�3�&#U����Px�m%�8��R�i���YX��߸-��i)�u��$�?9pe�F��KF�؟!&A�Pl������0h?�A��u�u)��әFN��u���?�A�	�s�)�oD�.�M�F�4(:�v�R�ׄXn�/�l�?��/M�nK��P>p�O�B�ɓ��&3A�`��߹`]���7}�-�5��	�A��Eb�o�V����Hx;�k}����	 U5�������Ap��z6�U��~�&Z�?al�U�#��	��*�,JD^B?���@i"�*��:-C� �ךj�T7kj�M7��"X��Yp$�dT���:���o<�6�B���'�Ͳ[�����yݝ7)	Ɍ�}��X�슖���̍��a����[�A!`�I�'5g+�?c��/SRR�J���FW���p0��F�J^[
���`�v��cܩ�r��]+�(�E7VZ���!
Sm�S�� �I:��5���C:-�q����Ok��M]z�!8x��,I�0S����[����A�����")		ys,��T<���g�T�\�g����uf�^�Pqx�G���wd����ǝEq���;�+0KT'Ł�*���@���lWK�آUA�Q�)�^�Z�A�>����Zg_�B ���Tmn�^�]@_�|v�a��p�v�ӎ�&���n��z�������F�`n����Ӑx�R�˞����qJ��Rj_
�<�M�s� (������Ɣ�T�K���'�z����%�U��h!y��&0Nq�<���wY��<v�:�nVϕ��k��҉fA���1��$k���ҷYȢ]5wn��A��f?�U����v+ဈM���ҥ��ȼ���r�h��P7D_��6���ˣo9�FzB��0����I�u���>��n:ɷ=�g�� Q�Y�pO���wq��/�)_q	��MY�l���X�8)�^xf͘.�o���ҁ;���[�A�
lk1LU��J���JK�߿�UŖP��SD��v�nV��p�0F]D�i"���$�.]��Hџ��2�]U��E�yAؐ>���%�NV[k��|�?�8�K��yv��p�ȯF���@��ҡ���4�?��݀�VP� g�F>����bg�gc���ĕ�ߔ�F5DT�&le{�
΂y�Sn�&��诔h��e
�� �;s5e�JI����@K�T�xU�vqգ;֫j��x#8�0*Ȯ�	�:P>s�s�6�a�N棞g�--e��A��-d�DH�	q��M�ʦ~bi]YG�4<s�0�&$A�<�s%��4��	���YP��6Y{i"8���¯��
�'ɕi¬f���/�hw�br/��w_syi�СTx�#�g0$Hܹs�d�lXV��w~�cr��޸/F����c�tGW��Þw_е���2���z|�;��$�6� ����ȸ"����اd��w�-8�&��2/캶�g�V�Wv*���R�x��5 ��{-���~$Ӓ�M!,�'�J��ſ�4y}"�
����l����Z���یT�܃@��Q�o�@����rQ��$oj<��,	�t�;��W�83�W�Z�K3�$(S7fk��0"=�t���4(��q-�䲕��)���2���G��]>�"A+(�ޥ�(4�6G�!��h������Q���-�C��7PU��-�GY�`j��h6e�i�H�F�l�ǚ���t&f2vd�l<.�O��M~n��P��K���e���B�$}����wY{�h���J$;��U�zt�1\��qm91M�k�h����#�C7��A+>������|0�=r��U\�X3�KCd0��������s�;�J�p�+�3aҪ9�ю!��H�
�cr�������̒�fk��8���8W�t���,��0�E�����l�@�4@*;x>բ}R�i� 	}o2q���_�#�X�Z��AoaV\H|���lI��%Bem��#�Y��X��(��m]Ὀ��plIC����R�mB���b �q�6�zB�^����WD��=�ޘe�U&x���5_��S�Q���\)Y��lX]�<h˵\ww-${R�[�B<0���ǖf&>Ù�tj��s�4� ���H��5��P�;?�}���e�o�if߶�t' ��" �m���$�$�8<C'��6*�G��!�(^��F�����qG7�������*v%�����y���[e�?����.���ՙ��T�����.CĜ�7�ĕ�EA��y�PĢ�ݰ��Ϯ"���9l4���g���IkL�%#�h���dҫ'���÷*��`�Q/+�-�͂jĉ��WI� mB�f92?�c�g?�>�q��]�m"B{���'f�+���-�����,y��%A��{t��1��>��
�zs���M��n�8���E��Ֆ���F����[��jL	�(��^������
N� L�D��B�2*��/�h��pvc���7�) K��#�k>�.nP㙿�usX����)��w"߭ػ�ۨ*rA����}��2�9���EE��n9- ��c�9/�7H�S���ts�%�j�7j%}C���H	�c7�j8���~���-SgéwKp[b��![)*�x�5����Ԏ)��VM�8��J1q�~�����v�
Lr4�pt�s|#�-�X��e�,�8q{�<~��4�}e����~���s�r�%B�9��9N��7qm��r��F�r|_�+}"e��r;63U�v�I-��
�T����PɆ�f[{����B�����3�Qz�o��h�Z��+�,��)BT��P�P	��7Z��Y}ic��}<��B�8m
G��iZ/A���z|z��}.
P�Q�j����x7��f��ۚ�.P�Ze��2s��M�t��F�Vɭ9k..z��1Ed�B�l������C�g@�6�������)�%z{�Q-Ɵ�Y�*y�H~Ȓ�Z�����5����h~"��>p'Jث���JWGm��h3�����;�$fq}S�|��	�����*�﹩Ho߳0�'��=���г�3���r����k3t�kW��)S�7˅!�:޸�F�4�!��BY �@Ow���y���כNi
S�-�ǩ,Ĕ���ु��	�/4�3�2�CK��p�e��Ү�a]���g��s�̄�w3��I3kxxx����	�v�1c�ӼoL�~0N���!G�R��º�V63RU-�c7��v�޺�x�0j��I��	�Lz��l¡�$��7�&�a[�T$�c�64�|ZM�l�̔in�0�&IQ��'���4��.�2Qf�����U�i��#�1G�l�BD���������듮`��?0�?����3�n�Hec������O#���l�t��y�U�p�ߍ&��y�f�@�N�a7l��D���6�#D5h�K���p�A� =�qɂL���~�����(3F�Oz[��SN30�� Z�y���D�	����?�PF��x����๏�a�n9�fq�<������� ?��}�z��:w��8��k��E1�Tw��ʙR"�?N�2,�=�aKφKZz ��(��=Mo�1k����h�#%/�!�5Hj =����fv��5���`��s���[w:���|�v+ �f�AЁVoҊϮ�O �*���-܆/��i¿[m��o��f�ڜ�E�U������r|d�-츓�'U����CеAI���AZ2��z�����`j*�8Ŕ@���n ��q�k	�>T!�����������qy�Vo<M�yCU[Fև�Tk����L����+Z��'~>>��/�g]`�����l�4gڮf�<1e��J���>�yQ 3ǅ��f�7��{1�-��1-L��9��*,?MQ���&�z�N9QjM"���/mk�l�#�M�\����+�!��W<m����`��aǨ��E�q��"�n�MaU�n�������ې��j]ѡ���?>��n�<�.Q�;Y7��؉q;���>��+k�*������Ns�6�i�L�
��E̹�֘�O�ht��"��E`T�������I/�'nG"Im#q!���ι�Y7�@�h��r�&X�r-W}x�;�K�tDsf�H�i4�9xu1꽮��E|��?~��݄��M���@~d�u��9� �٧�yE~��%D)yj��D�'פ���N���HA�5���p�G���r�dl����o_�Vpפ��_O+�We�u$�n�sW���7�,�m����pkQ�Ԫ6�qU���Ԝ�y+`����n�v}���4PuF����`�����R3�� �ԣ��Z�`�ꢙ@c��p=M�G!?��ŘuT7����t/Q\M,6=��b�����L�2؝>6�G����@�_���$!�g��#�j�9a�5{�8�q�qCC%���*U3�6�z�]�xy�})�zO\�e� ��?��=4�W��xEe��De[n�s�J��]�����:�?s�
?���H��=�f5�#̳��{i���J�������5i��Q-�̽A[�fYA{��I�e��;᦯�ʭ歈ܵn�6H�{D��Tr��DO��� `�Nw�T%NC�^F)���Ʉvz����g�ZR
7�7;\xw��=�c³ε=�B��pa��)syF�	f�%V�s������L�\��Zc���K�+�&��		�	_��;�v�H?��<=�o�R��*FdX��������K��8,r��'�k��״}KL�?�EV'�������(q݊�$1�5+�kT�QI�=YI�W�����)S�v��Ǭ�H!��.KJ��p���x��"1��}
M��غ��670���@|� <�a5#G��#�_���,ki[I�vR��W^B���b���2��R�朳��螬A~�S�LM�%���mN�K8��BS�&A�I�@��u���
��t]v����b5dxD4U\t����Ft�\��)��}��eL{���T��64G��,�^�7sHd��wm�ЃW"��O����{��琾�]� =��ll�
�VC*���%�q�k�N܆ࣴ(O~sCx왯Z�y���h_~{{d[݆r<�i��c�S�KX�(Hy,H�֪阸����}p+jA�UN��u�����j�����H����-�KJ���f�G�Qv7|�� �p�"��o�_��ܾ��+�9ӝ��e���x��L['�O}�L҃��v�h�r�ư3�.n�7�2$m-d��G��&׹�X�D+`om��1�|�bB��K����CGӼ�]iPI�'b�¼_淀7�`�>-G,��}l�^!]^c{B
ϋ�ȶ�ugR�r����e��@ .y�����m�f�_�	�P`9`��V��ӣ����Y�7�����;V���,�����D�N��ttMZ�ƕң����
$�2垪��?ʧ����]���:|J]�~�V#�W:կf l��0A�I����<o�@��vH@�e��Z����r��j|W���<�8��K4�d�ǔL��Rq`��}㮇���>�`���o���ԁ��v�η��n�;c��"�²�(�o(�S�����E�2[�@�r��v�i31y���P����ܥ�w���@��w]�䍃�|��=�MȪ���r�VT���L8�8�f�47����4ΞJ��@�ڔ���t_/C��lx�Y0$�����<f���-7>�[	��$�>��P�.�1,�!�
[���5\�:ʔ璉�/4��ҟ�I��`g�S����v�z�U(���4���a����s��0� ���Bu�Юd�g�@��d��A�aŜ�9�|ڽ��N�&�f!<+[�A�r�X$�k� Qwl
����X$䔏ó�ʮhrH����T2C�$[�
�A�&�N^0�+kd�qg@���F|!p�Y"�����P�XW���p�n<�ﶅ�_7��{X��Ci>X3���GH�̹�W[ f�=��0P{���E�����q(עV'+���c�ɿB6kkII����%;W<{^�F��1RZ�0�q���mH�Q;�.M\ln���^�"H�j\4�._�%ގ˃�r7�.�	oZ��*�#�l�
���,� |Q��Z2vׂ�B��t�{_�M�\�^s>t�``���;��S�ƁZ�Z��ʰ��'r����>\�{4.F��(B�@�ݸ�G��D8	�Hɒ��4��ٓE	Gt�9�����Q	ͯ@���V{ˀ
"BB��D}����'�T���9mW���m2h�/녤E�w򸙦�oX����@��ٌ�) ��W?��~ҶoXV򬭣<���Pt�چ!jWe���Ru�?�nk��*!�Ӌ�ݽ*gz	���8G�����E%b�O�{6��-K����oR\	�Y`�-��\9jB�(���in��(�����>*�[J�Q.l���n+.����6��K�lYn��L��L�21�_��.Ю
����v������!M�&�1���#a	0׺G2<bf��Ff�Q�]Đ'�^
�\s�nT��Uԝ�Y�n��)�	P����/�ىBׂ��f��ˌ\-8���n����@��=�-��W��/�(�F�ٓ���li�Ҙ!' ��g~�\ri�U�,XKm#��X�����Ǜ����S�ݍ~H,d^�E/|�A0��gU�_@��T��E(��ͅM��-.=���\m����Ӟ��+N�sdIe�3qj�k�2��4K�j�_��υp�/��2qf<Đ�
6ê���P� v�tZR��U�S��a)nБ�W ;�U��"��C���~����#���↟�ݞCPh��ӷ�xƕ��#2����j�
�-�w��K_��vE��x'�+8���lc ��Z&&}���Bm����R��f$��IB���|eB�g��l�r��J�_%�p�h�b���],O�������5K�|���q8���놵�A([�ۇ>A�~od���wy�.|v?K[<�оGS�|�q�$���\|-��oٖ��F=2a�_��%�к�Y�&'xʞ��wj��&�;[M�ݢ��불�|{���e{Qe-����u���Ǻ�4�Q��y6�f�ќN)z�Y��h~��9!y�@ڸI*��.6��Tү�S�yb�崌��k�K�/��;��%{�U�A���$�{����KbF�[g$\��`��Ȑ]�q�z�m-�^Uƛ�����gtΙ���#�7h���.�H� �4HC��b�������%��M��ĵ��K��gEp�i�Be��������n��4Q 5��x��ބ��w6��/s�Z�&Mb̨v���k�k�8m��0�g>lR��&<j]k���P��ˎiu���'��>;.��K6R�;��cO
2��]� �]��t�h��!�Ӵ��AzNkc�`��ׄ���#�("�x��P-��GfƤ�4�n(�8eݝ,����b�Og�o%x?�}	jg&��cr�˜S lieD������5um�ؐ^�s+\��62`b�:c��f�a���֤�Ŧ5�@H�Qt@E��#�_�jF�� �; E�;���lr\��������v02�r�F��AP�Ks����b'��a�9h�+��a�-�/�!C��L^�q���u�����NK '����-�ݯ�v�ґ�j'U�'o+��R9y��)N ��ZY5Yc�r�wĆ�\8�X�\_}3���`�v�F�J�'K�~h�>;�#�@���s�OY�R�����~~�UDN��Fڏ ����D�lHMf5������M��=�C���O��v˗�yn&�ҭJ��6����ڹn�C�4��v$�A�HB"�ƚ��ֻzNVutJ�B�D�aw�KW����G.�V��Ka��E�M;v����]�{-��'(u����{^�׭t�7���P��^Z��NZ,E�gY8GX��nzl�ӏMK7�1�)`� �8\�:td�O�o����` ��o�p�|�5S�hH4<����B��q֡+�"`e���F \��Ŏ�	H��Q��ĥ���?�2�(%E"��Y��vtj�Z�X�^�e���~����Ԯ|�w�w��*�Y<����ƐBc5�v�'�8޴���r�|�]}�4�KoJ|Q#!����!~�~�E2�H{�kD)����wI�1fB]T��V��%���2�$zT����E$�>����s�v&<���b-�њ-j��I{"��hZ`�3�H]���,�z��y@���0��f���'�hZX��s�@�"K��3}��|�ك��m
v9�a��a;���9n�X[@3�!ZSS�f��u����ⰵJ�C5D��ҫ1�XCHP�8�b, r���*ҍH4,�E��СTPϚ�cWy(�ٿ�[�E�N f�]i��h��#Ғ�l,�	�wX�i�$좿���f�/?�����W��>?��_����J�J.kqW��ޕ��u�?��� RoJE���mD�P�:��v�sr�wx�H�.�n3�6�����đX��'�Y��:N�q�]$~W�Un�9��f+	�Z����^����\�5���AӴ�傜�K<�z6EǖTQ�\z������' �{m~.w~��{��5/_TTHYj��T�b��n�քY�������#�{u��;��xJ�á!��Gw����7YGkm$C���@�Ƅ�ؚ�j`ݯ
:�d�6`D����Q"J���m�@{j�Z�j)�k��e�Ţ�2U�.sx���7RO��R�s��RbqD�X�n��y�| ��
A#����F�0�k7R_C��8���uE?Bf�q���h�ӣ�z��M�`��yP;ŝ7�'��~Mߣ.3O���ڭk�={(w�p�0���y���(�w�r�
��3���AC��z6�3��N���M`�S�'��r��W&~���b�lS����'���B�ʫ��*��a����y�Y�~���S���1 �`b_�`�n�5���g�$f9�H=���B�$^������ڃQx\����hUQqm.��gs���csb����:,����$[�����[`�۫uM���̓Dr?p�]��k \����B�jl�X��$�w�+�S63��W�e7�%^�b	#Y���p�qpB�kU��ӷ?�� ���8�~��ZK���y޻|�������/�����7s��-�>��١�A���F�2)����]��.>2��K�'[�t�Q��u6!��<C�5�.9�2���-�C�&f�{�2�;���M��փ�%^�.yi�@��P�*��SE��E�R�f!���~� �A��E���O'��߁ͼ"�h>aȬ-�|���^[~�.�m�)��(Ě�ɿ��SVZKف���*�Wy�J;��ɥ9��ex�d�T�G�6��P6m��8m@и>�.���pH�ޗe��������0����2 �t�5+|4:1gmEVS�J��l�ı�S��J�W����%zWl�"a�88�zp�*�ԁ�;���{�y��B��FV��@�H�u>Pk��);�}������4Wa��K�d�Ǉ0�G��]�´�x���2�@����eJT;�'f��ڑ�����8�D�6ѣ�����O�G��|K�B�T?NN���*%jU	�%0t
��u.��X���oV%W͸0���_����\�EA{#�����O"��u�Uֆ����������R�ł^�.��.����!xg�[�l�a�6W�uZ�?�
��@�ݩ�����36s��WY���|H�I��Ǉ�Rq�Lĸ6y�vL!�\9xwr]zh)ظ{B>-m��W�k��y=�f䥏c�S��hL�|�-�\%�by؏�[�&H4|I��u������Ō�k7	E�	U*A|�ws�gyES�̵rHe՜bH����Z���!_i>s��I!_�{y�vs��&5�����#!3h�J�9�0���Z 7���-FXjY��UT�{��:�D%� ��p��:��
�oW�8HT�x:���Ȋ�^��4�iwI�6�5��`'p�Q�<J�����̈́;��|�y�7D��1MO]��X���B��寰=DP)�]�n�Y�Oj�]V�/j�ck ��LV�@���ăAB�:ӳ���s6^�p
����]��`�F(���N����s�{p9ۢH���-F�xv�}z�$�t�����;��%�a�W�?.��-p�_
�v�I�7mM�]�I��@:�X�Z4�4&�l![^��v�Gh;�^aY�BV�ֶ�P� F2���!�Z~]�e�q��w���#�Ļ0��M��3��"�w�2ڒW��aM;Ӣ f�`Qi�f�Sݘ~���v*M�<��}�ͦ�~�����\����	�-�vxDIR�=��A.<�S�l���,���aP�|p;~�=LC]������u�k���%A��|����+�N�.��e%�ɦe���븏�,ا 6��K
��w+	���Ù��a{욯z߃���0�0�LQ�׌o ��_|t�l�t�c�	�3g:#*n�C�R���1|ߔ�AL���Y3ձ�V��Dג�@�d��q{��7�a&�F�y��!.��z&g�k�G�40��#������
h�"Y�%�Լ��pS����]Ǡ�
o&�[jl#�N@$����
�Y.�gJ�d�+�r��-gs"=Ic�"Z��ڮ��v����sP�l��:S�	J��zcNE�Օ��Ar���3�͝M�$�*�"?T��$�B�o^02�3/.'?�3��תj}�Ffo��ZTc��٥��w]x�Is4����5k��7Y��[�e�{Aa��)� J�Ȯ�²f��9�j�.X�6��'���m���xC�q��~J}���Y;���`m�z2���gpy����iu�=���+3WR�[������[X���*A�ǃŅ�:�d��ʲ�f���2wlSO��(���M��"G�����q���
6�D�.Qc��Ũ
��T���,D��T��`� �m����_{I ,��u�P6K�M��:t\+RM="e�������D�eL��*��[S�|r"��"�1MH������<잛2KB�p��_����-�mW[t+���Z삉 ����}��w�@@H�l�:&���>=�q�����@J�����3*j�|�Ge�T�������?��GȂ3/�s�7NZ��8O�>8 ��N���;��sn8�
�љR���A;E\����S��=�:̪��=ܸ�k�b�k�*������tzM�!4`�<���ʙ��5��7*�\���nE1���K+�
�3t�n�DJA0=��������s�*[è����!��F������9�Ƨ;ike���q#�o�F3I��y��w��n�E��<,����6$S#�-°&C��*�+���Gl~�I�8��*VB]l��k�']���+⡞rp��ܩ߇�=EY+K����V�w��7�ՙ����J�w��%�jS���Ѫ�/I�193�^��}��"�$#3�����L�M7���%� �iz�l��l���ѕ�Z^0��[��562���\��1�,<.�?Z����Ğ��HDi�E�ߺ��$���<7��w� v��T�`�C|��O�6�l�hv������+E�Z���b��i9�%�40ݗs"� E�ך>:Tm�Xi�m�U@$9X�,K�|���u�lz}Ћ�{N�14��eP�$� ]3"��kU�Yڨ��� ̡�9�a'μ&��W��X��D��:��3��j_�%��ܥ
���'�!�+���J��o�,�}qQ�4�Ҝ|]=�#G�OG��r�r퀣$bB����Z"!O䊄���tUa?�bS�ܡ��A.��mG��&�!��E+4�OA��F��^���؃�I`�|5X���S��Ρq�}9��f�{�1"�*��8�@+��J�2̈́W��l_F�GGY�/%@u�5T��x�p�X�QM.��Ӣ9|�N�p���=���"6 �gB�Z��'�5��f��]_y\��Nd���D���,���m�G8�=@|W	t,�tf~QdvP���%Gw��k�t�u���Gp���JhF5�J G�m�����N��Ko�e��Ň��!�Æ�z� gټYS>��9sb�b���S�	_�ذ��~la��ܪ��C�G"�>�Y�:S}PLq���&a(1����Fu��:*Z�E�cA9��e�,�87~�������6�nOV^H����/��	H��	!x���׋>b͹y��G �_k�J˦Q�t%A5	������ -�9���,QSH�q!O������Y��㔤ez��dF��Ld�� �e�}[R�a�3NL.i���Ђ叏#<'�s[LG�;�w
�zOtzK�"�#��pXkNH��(�I��ɯ�tʽ��t+�l!sтذ�[�Ā��v9t��o����P��k�b��F
7��}<[���~M�/~�U��*��:�e0��&�����6SCVO�`;���\\���d1Ь���K������s�9�ZRxI�j^�I��B9!�Yz�����_qݚN]}�)���V�^9b�A#���$_�~?M�)'�w(9���|���L�4��k�U����	�̑��\T�<h/a

Y�]�U�ד�`r=��5
D�\������� �V/J�)�>����J��!b�!js�NJ�;�Ra�n!8C���w��/��������r�,�%���@\���\IEe�EƟ^�_�$F��V���f�b����� ,�=C.r�%>wG���b��6kV�NF�k�;�Ƕ� [0�\��0[���X���B����\G��ҕ�s��_eRJ
2�h�l��d���T��5��X�����=8a���Ҩ6��oP���F�h�k���FD�E��z��P�ڻ��D���f�8`����s$��XdQ�=�á�D������C��ފ��b�<�G���h?յڻ�I18�oc��~=95��Pf�$�0F�[Ox�p��*�cm�X����TMSj+~�o�.���������IT2 �-jD+���;k(h�/[�H|B�=��b�\�ɺ�����pCw�f�&B>_�xo|�	�V�8�^���k��7+�����pI�)E����ݽ,�K�sT���(���3Wr���37^9�J)"O�?��{/O�:W�GF4zq8��b�J�z����u�6�t	�G=G����&����4�!��7���_�Z�l��C���\cº>�&ǉ��A�E�6$��JN,���:��Lt��to�0��V��VR~O!��p��B0��&biX:WLΏZ���}R���L��O����tj�?�f��� ���7.G�l�t,n�֐r�Ҡ1��j�.O���6߲tw�(�%�t`-�p'l�H�SLnDz�*���G�|��}�M"=^�v�|�oʋ��i&���L-����:u��e�LE����s��2/�q�q3��(�����rP��)s��3p�]���^xp����	���+�7DwQ��Л�_A�-����H�U�4/
[������+u6ύ�p�b�p�f����t�½o�-�� [��n��i��q��d��㱑�l�gF��`����Bo̩`�!��������n�i�l^ٽ��=LCHת�)�����ͮj���|>�4Ȕ@��j������W���>�e�?���p�XC��k����.�C��Z͚l��������sl�"q#$yR�3�Z�Rz�(/7����Ɓ�C�"�	�rb���3S���s���?���f�\�����}�s�:R����WR���-�E®�QX�g�)Ha�r,T�Q�!��&�N��~!څ���?!Uf�S以���W��o^m�?ʚ�"h�*j���v������M&Dc�[Q��M~��ϯdM|,�_��\V��"�CD�2��,D�.��y&	zv��P�@��L��,�K=��zT�VB�����DS=o#�M��gDn=[��bS���~jm���zKۊjU��Ü��b��\�=�B�6�!��r�(�z>�,��K�l)3>�ط�$�?�����*���1d���`�������='4PӦ��n+�WQ�H�J%�!ڪ2h�Vle[f��8�g�&�5�JqE�^g�{��a22U�RB��0{/�ȇ�F�o�ֈ��'��p���?��.:������� ��u.�$nu��3/�&�N�x����_�� ��g�$M���_�g�y�n��e3q�h$�Q+�0?(��9��AC���H�	��Ɇ������=/ ����j�?cCgMq�B����)��NdD�%\���>k9��-��Ɩ���a��y�U�>�y�w�h�$VZ��n����{Y"�`����U�!:�[�j�9���7a.q3XpK��Oj����F�Hu�����5k�6���.�����a�UFJ��Yh��Mvޯ��V��\KZ��=V�4�`�na��B���s�����x��ؒ+���Jno�й�xzt�|�26�-U���##9��6��,�ln֧rʌ��#�X���ev��CA�ۤuH1�X}"���k�Y�k;�Q�r�:+O��y����L(m����wT��r�=1n��(��P��-�7���`HEx�0� ���	v#g�� +d���_��x~ 4;�`�S��J/g��.���}�zX���/玃�z����97�弩�|�q��ߥ}���n�K˾[����}(�[* /������������o��~��]�Ϲ����U��	[���,?i���ܐ��U Y�;|I�G�SD�����td����V���3��6�g��XI
\Lh�6��f��,Qu�2�i�����D�X�&��@�k=�H.=�s����"M)���a+��R�Gm�Ҷ�`&���]��ן(F��dmڍ e*E	���%��Z�.3���~{C�F���Vq������ISƥ,c0{�m��c�x�o�,;����VaaB�|��G�͒YW?��J���Z'+��h�іZ>�#�s�Z`�N��v��s}���E3����[)�H�IŅ��/�HV��H�;)����qm��d���'�R��o"PȠzc�gX��E!�cI�}��s"�:�hYu�W��z�~	� �N����ՌƎ�:U��/��,FR��y�oJ��I�4:fO8������Y��~o�\��9��|���)hf_�T���3ҝ3n�Ռ��+�4-�k�h�9�/�l�܆����}��3\����a���~2[Vp(+������i\���f����J���[R�eW�,��P���f��jVޚL����ˢI>����a�K,�9>��36����e{�e�u�B�L�Tޥ΀��
��dl��(���
�\~��Ę}���x�V�<�!Y�X�@R̷�f��Q��<�o���ZQ�I+�`Kd�yH�l��
�E{�R�>;/�.��K��8x�Z ��c,�cR�Ox���|�w�����Ԣ�\h��wz��P�6�]O��|_#�H@��V �3��v�O6x��Lp)7�[x�,ۋ��
jg���^(t�C��&���ߩ(K�G�0�Ԧ���}��y��g;ٺ#�5j���q� ���	1��Aa����`eAJ|_�ֆ��t2q�֧h�`$Z�sB�*L��a~��_<O�^�$�v�V__E�W�f������uF�;�ʙZ��"��a���rwz�h_�O`oaQ�F�;?�c�%;3W�A!Z�Hڟ&�5O�+�@GP2 6x�מ�f������:	���^�~%]���ϐ;�@A%�|�w����S\��3��w����GF��-T��)yZ��� ;���4��� d��y� ���JV��K�C�j��*��,��!�K��w9��.=(2����p�*�,�P�Z�O�OIr����3nH�� ����.�	�'w����#�.�}
�����]4;@�����NH�Y� Z�%�	jV��c�-��ٹ�H����DH�DZ���eWĩ�Ro��a ��9n��!~[����XdE,�t�}1,�)�`ˡ|��)��G�?-
TT yo �2q˵]�ſ'\�.f����z�[y��3$Eɪ��w�"�p�V�l(��Ǆ`*����R'K|��<��ѱe�Y)����Z6R�l�ū��.{�� �k�I�b�����q�
F��2f�A���̀�9��į'�i(�f���o�?J5��8<�e� f��˞W���Oa:���r�%���#�NFJ�O~����3�=��W+��Vb��̕����� )��.���q�~~���V(,#��Eoﰠ۸�
b�\� ]n�=ƹ��!K��N�Af��Wx����'��CDl1�4���иow.������a��I��;[�8�|�P�禘���`'�Y3�7��Û���>	���2�O6����#�ń�K#���#�T�d�M&�����%בF'o;�Q<��{^��у��)u�j��D�	@�~5���vU<#�
^wHDZ�h˲�]�+���R�j���Z�yF���zL�,��	���ƺ�N$IL{��s�De���
�0j}�4Y����۵��s'#!�=����r8��~�[=���;�z2�Nt��� ��'��O��C(����w/)�^��q�	��:G *Ҭ�&���T����I�|~Hv��0�P����s��|�D�b��}�l���o'���q�ٳ�(b������=�2����0��^}�̔TZ�w �]ܾg��Ձ*�Ͽ�'�2*�S=Ce�J�)7�l��}J�vK�����h��@*�F�J?R?�,��S�6T1M��kE��67�� u�m9Ay*1�"���m��tD᾽Ϫ.H�D����~��x�H�?�I���N��%����.bnO*�S�����2UOx�	s��`�0^�iO%�-	���Co������,8k���BZt^ꀌ p�ϨH
�U��{�
�b/I�䥠��̶�1z��������0M�Ex���D����$쭳y<��ct֑�Ǩ�Cު�d�s��ZR�n&���$���
��N����|������%wP^
W�h�6���a�^�F��la��(�CP�_͑<�Ѥ�^��#����gM.����ŴE�x3<'`�j�(��ާ� Ud�il��i���F�"�"o�.ݶR#�2J��H��^������v��͕���f4=棸�@��-x�[��B�)�V��ʫ�����t�˹ς5)�+�@'YJ4n�X��Om�fX�����v��[��/���^^�?S.{7Ś���hs���:NUpp�wn2�w饛\N�u�:��C���gE�IH7���۽Ň����FrC`Zq5,�<�6���MWN�b&_X�n�ȬF�p�(.<�P��=�^TB�ΐ/�(��a6����ңu�.T�(��)�Ķ����Z��x�@�?@e��4��������Aۧcč9�%��K�|�ki�^���mPnA%��WC6�E�45�Mp��*����ؚ��Ď���\1=�����q�=`��E!HsNDwL�M/�Y���6/d��D0���jX�^�O+ϕ��T�Y�J������K{���&�k=��-���|�q�ؾ�<������w;syQ;TE�q�s�H�rN����֩��j�z��&�m���|<E#wƹ���c,�7����3L�lK���Go'g�+S��;o��9'��є�}H�ree��L,���<��Qa����� 5B�}�`���J��<�rHd�g�j
�SH�=��l&aSV���Y�(�kڔ{�j�ą��F�Y��O�{�|����bӨ�.�?a�(䈺	Ԟ�Udwo�P��QJ���>���V�KSgd�]q!�ԺJ�n����J]@B7���`γ# EIJ��@���v��
Ю����k]՟�P��,aB(���hO-�#9f0	6f���,�]k-�W4�Tw����k�X � ������,Ӳ��G�C��HeV�-����'�Ց�_*9K/�<�M����z?�4���ESR����̎5�$� Q�)�j�9�)_��̂������u�(�����k�~�:���?�1]�c��ዧJ\��4[�8~�X�R����`�zq�V�q�|��/8�>�>8��� �;�^��}M�W|�Ӏ��X��Lhd]7�In3���ȼ���o쿳���An�6N��=��Sߵ���֟u/���
9A��Aʽ~�~�Ǹ�DA��<�2&� �Ʀ�����Λr}�;��(�����{@�P�#+��:���{��O5_���(����<�`Ζ����R+|jϛVuf�0������K��js���%G�!�r���&V�r�Om�p�p�_~�ψx��C�C�(���:\o9;r����4��V���Ϥ�`2�4 ,y��͚���+��l�[�t~����n$�YZ:�7��y�L�<��rl�/rl�v����z��Y$�'Pabg��q�f����;���>=�%`�r�k�s�v̉^�Q����ԁk4q��i�I0�(!���՘�u���%!�%\���n�܎��L�}˯@+�j��Δ�b�*S��^��j� ���I�����7���^�����$�U�#L�R��+b~�1mh����1�(vPJ�>�/�J�P����z�H���x�|,5n�a� Wi�\D���7�4j�� K@N|��9D[�s��g��°��˔K��_(~�oGB �#�V�$X|z��E�l���
W�|m��R*��F��N W�SuG�f3�.����`�Ř���Z
n8�$qMb�J�e�;�ܝ��tts�]�c�Pk�E�-�׺���t��[٬o<�\�K�S�8o���d�!&@5CCp?����dtGdd��_�}��ɡdc%N��3f���P��
�n��x�V����<a�z)
���"�X��%0�+�:=m�n���{����L��/�������,�)j��f��6F�hO�[�t{�)s1l�(��na�C��:4���ȸ3pv�JV�"�et�OS��ao
�e<�����u����v���9�:7T�a�$\�P)3S�4O`<�D����=ɒ-�l��R/��y~l�����?~>w�Q��}{�2 ��h�8��;�P���|*�iqv�,�Asj�ZM՗��n'��|.�Do����n�g�[�`6p�Cϴ��[Vsl&m	�r`,���A;Lc�)��5l$�I�}�n�[�50��_�AԴ�?�9i�7�+�:r�ے�j����R=�TN�C�\|1{�B{%��d�T��0��J����|� ����U�(��![����f��)�d����o�G��_������������=�_��t�n��z ߛ*��]f�D)1Wh)��|����?�ڻ!=����9�j�{�p�U��K.��+��c��Ҏ���R�7|�%����_�L<��=�Aņ�O�a7Q�����q-��x#gN��8����gs
����#�j��f&��(�B�PNŢG�K��b>"k�2� ;Ѽ�k�k��d�G�@5i�/z-]���DP��L���Xc���������gB��{DN�[�<: u��H���U�����}	�&���ȣs�-:�gO�FY��9�1�Yg���~FeqK ���?�G�DV��}Z�#���R����׷0�v�r�i�wf,��N�� �s��N]�~�s��8�ײc�E6���X!oK�)�U��U����"��n����,Uʑ��Q&�G�*�PN� B�wr"� �ɴb�H�n>������g�*i�"�d���bM}�Bc�Ir�>q�<�/�4��v�[xV��G���i��:��qB��ȋE+��B��,�^$�1�_�U#����t,�>�f�_F�"��Bܩ����O�AT�x�1g-{'���_��<埅�4�ԽQV�)�<iyxOO;��+�H`�f�;��;�4-𖭶!�v�a�_�7:X��u1�%�۴pM���idcXғ�bfI0��l_1-���X����Iq(�h��	>�Z�$�t �5ry���@����/��D�a�ӿ�֦WR?��\�r&�p<����4�
6���y����l�4r��u&��
M�x�c��0�\Ekb�JNc�_{����%ϧ���Zq���Wzw�#ő�ڽ�Sa�Q
l�0�\���E�t`~�	�Z`Ay�b��0�jR�8!^�F�L��%4VͿ^�a:��р\Qb��Q����=���'�m1��\i��iIZݡ��1^M�X+B��sCKd9#�́�i쾦�z�u�1;ɭ� �05j���2CW��X+Q�l2�/�U�� *�q����*����%�*�xc����k�pu�'��o�;��o޻Q��ܒ�-��HPт(Oq;1;_���h����F/�(�Ir�{���k�<byIEV�Ir���g�u)�|�Q>����zH9E�1V>-�v�-&��Qm
��E�W�
��drT��3�>Ʈ�-�2����j��
��U�hn%�z�qB�Zާ��^��M���<�5[�����cx
��E�m�{b�tݹ|J�y)��}�~����p٣%/�"�%L*l���r �NՊ~��ޜ�(<z�a��S�&�(���T7��HCj��⊒��A���L���l�
'���P�����&R���=�E�� U���(o�˥Y}��eHt�o���2�g}���/�ls�H�4ߚ%��2"���WY�/��V<م �8�Dm��~y��P���w�Н�G����G#�/�{���u5�!-�_��Q����.��?���kAc]zǖ�7�r(���?��|q
RV����oW��_���FPR�Ȃ�%����S�(�5���s� �Օ��xG����Im������K:St��*�QGts�O)���wv�÷?l?���l;Li� �bV�x�H�F�l��	�7?�/�s&}�'��Z������
�!:8QII"��f����oE�&#�El�J+Ћ���G�!҈y���� ���]te���v��)�"�۪�C>KC�#z����*S���։�y
�D��SkMU�0!�Ymv
�-<t��2��$�\Q��
y���}�T�J���N�>/xùT~��.f�Jƃ�*0��x1�svhi�ٞ}~/��g�M��+�G� �]��3\�z������J0/I^-��>bʂUB�|6��PXTQ���B��O�Qkojٞ����2
ݡ��E��*)��$sJ�N}�	Aعvĝ�oCWX��j�aa��t쬍��a�>��)���*�Ρ���ם8�S��,E�[DZ���9iR�{�
����D-�4�ۀr�VTw�P-�;/uZĪ�/�3��1s/Qh�����#��>	�u��\z�d����%�Y7�R;Ls�:����/��z��9�1�ĘRm���yw�2��s�_������))v�LR:��3�Jqam�9<#I�d��$���=U�(Bm��[.}��ϲ_��FZ: ˌ�;Le���K~!p�G,�$��6������MD���?��J!X�b�zLIUyb7��ېב5M�<+967��� |�N��{a��N���Ƕ=���Z�������~�K���ub-2·~h��/��]�v������QU�iQ�%1�+P�KH�_vD�ew�`����Н���������=j>:�s����1rTՏj�������ı��&��[�J˚*��]�s�M��2Ru�^�e]��@���dc#+
0���A�c�d�f�ie��H��yU�_n(rm���<ef��4$PN�e)��W�w��ԡis�S^�F�Y��Z�$٘�QL�;���6�A�8���1�`4e;}�zjc=E9U�N5A�{����9WJ��n�B�Xc�����t������/��9� ��Y�^��[�8���(ghyX"��,����V@4��x���q�.����Y��{V��ҙ�'�F~VW�*|��R��e����to�н!a�T�
?�� jn{����6�C��n��`���ILx�ĥ��nJ*�Rݷ1�Di������nZ���^N��qky d�d�O�&�hSu�5��.�z��\*���MU�rX�%���Qܙ��z��pO}:�/7�aM���y�>���t��?;\�F� Z�L���u�${���gd�
&�ܱN��� �6_�*���|��=�+rO˳em;ޏ6�0m�|��+�ʆc"��7�ˌe��~7�m����d���'���c�_Dv�`�9����@�
��,�� ��Pw���b�y���zp��h��jĽh�P(�K9j��W�`6�<�t{*��_��$t�V��}�>���g��3o󺨝��j�K(C�����	���S�IB"�V�n�)Sb®&N�܏�̢��8��Uq�g!ǗE�*sļH�z +�2�X���7k@~\$�\<�h
.r~cy�����&��]kR�n��BPr���[�fAkLrET#�+I�;<Ӗo�&hcЉ6���[P�'�����o@o����uB����.� ^_G<�g@4��ٙ��gD�2I�������CYj5�Μ�ׄ 編���P�W�憛�;���z�S��C���8xh��3��b��k�S��C�Ɖ�n�x�L��������>ళYV�;&'(ȧ_�b�3H�ߵbݦ'��k �es��	H	U�I�5	 J�õ\&���'dǭ&h]�o��3>K�#�@Mb�� �V��_A�-��<�;����ѿ���*f�����,�[�Awf�s��ԁ����t%�~��Dw����oԯJI�[�E"b��mX��Μ�y!�p��U�Z{�tu*�F���UL����������$ �u|G!�����)������[��wX����+�^,�� ��B��c�y�8��	d��F�j��{��+�M����f��/���N���)��A wZR�O��P���b��q�Ŝ���h��)5<�z�7��yY���|���~e;P]��Sax��� ����(��iB/�=9�$��w\��=�o/!z'��]���H��F�.@��'���q�)���Fxd��������<<�MU܍ɤ������lD?tWn����-��0I�h,	�B��N�8�ċjER �X
�z�15#.�np�f/Mu�-�f˔k:�û���
q�[��<�j/��\>-��uȾl�X�Sa����.�=]�SQ�+0~#��QA'7Bƈ��;���'����-�	��s�E�U�������U��7�6.ǲy"�&��'�/�Cm �{��W3�6�F:�C{���� qoX]=��gj��P�Jǩ~O�Z�ri�>	�� ge �׎�,40����2���T�E  1�M���k�`�S�ƶ�B��>�܉�r�F��,t
&��er��l[[Re�veu���h��n�J��x�I!�"W�#�I�*@��e�"��/'��%aa2��-\l�nQ����ؔ��0�$\�	�l?sD��T>���*<yy����|"�Im��Os  ,`����H,��<xRL�?[&���Q�R�I���ʥx�̟���Hx_�ﱅ�����b2]}MÊ��� �<�KWS6y1�)=��+�	�t��������+;�a��ۄu�۟�T������C�e�w���KN��>��O���p�6ѷ���m�'�2Q�'İ@�ԑE�v-Gcں�?7;� `��p���톴?���k�4e�vŎ�x����ey2��I?�&P)Vi@]��nC����ܡҩ��x���cX��3yy)�ۆ�����zs��T�дbm��o��Ɔr٣Y���$��+�yسZ Q�y){�eM���5�rs��v*�3�U`3�CT�y�8�@�NA\4�ԵRc7��+X��x�ʝ�È�Cl*�N5���E�J������Fm��ќ�p�T*�� �)ɰ�Q���%�<����~���%K�����(	�"���FL]�o|��y�=V��}I0yl�U��o��_�*��r�4�@�������q:�Bc��榼���z>�QC�f��$���マ��7�("���7h�F�Z0
f�͘�gԔ`vdx0��z�\A�^dc��>����B�&ݷ�	{:x�C��o�jЋ��,"���j�R1�>P�$[��uO7�}u���q��)hQa�R��y�$�2��h����2}��| ���K�	��b����A� bd�|�*%d3���,���u��O{F\�m���ĪS��(� �۟�ޘ��ᙡ8�hAVkh��=��ٔ�-�r:i�|Z9E��eB�(G�#U��93݄`�C)�k]�3J2�B���V��չ�]G�(�s8��TR��b��!�i7 ����	Ўn�H�؜g֩��TVt�VE�O<Ȭ��Q�v�.�Ѳ7����!/���C�y�Ss��\X��RO��7x�FK�Y�F�#R�`CmA�|��+��G�ȁl��+C�(o(���W�H�*F%w��&�[�E�l�^ȟ�_"V��7r�]�T/�8��Q�j0�Oe�I������6tЗZ0�R2��Pgc��}����ֵ�8�Y��l�v>4�/CJ��&�΃]��vm'�5Yb��l��w����X}���	���a;��&B"���YW3������bݛrc��`Q!��G�BY��$�G�b�ڂԧ�UШ���!�u�H���m��,��Z�k4��`��w�X����j:1+~���S�Ϋ�L_���*�B��w����)��7��UT7�H7=(�C'
��e�p'�������i����}�/�ɧǛJ��?L/8�!�Rя�c5�"Rλ黠�D�܀/s�ő(t��E�?t�j���oY_��*��f���p��[pM[�-�(��B\"Q��Y��q�$r�IF���}��@�"svBL�(���I7;�pp���X�h݃�8�oۘo���K@��I� f�݁�X'K^o]<���mi�Q]�XH(��g3�U�-�-�R~�,�/�,K��C5	���>�٥Y!��Z� �;��qJ�J�ك���/%#��υ���@��הH��B5 1
s�=ȤV=B�`W]k���1d,�G
���`�F;�{K�k#�5�?J�!��H�����̕����Z�κV�:�~�sծ��=�feY���\x����gl֙�Թ��-a:�H�x~2�f�T5���ǐ�����=0��y*%19.��9�0X��T��"07l�eKl^P�J�X���P�)�k<�-����:祾���&O�U�_р+^������GMY�)�Z��?R<pא^o:��gG��!xc"�woL���Z3KȇA�W�V�������ɋr�:�bZ˴2L�0V�OTZ f���v���dEv���+"�:U�ՙFZ��8�Î|���QhK�4b0���eW�U���gG.���1E�P�lWe�A������>FoF1���@�e�:뻾g�ѡ$ân{v����H�-�Л��y�~'��T_��>)��Ěki�I�|X���5|M\[��û���a�?�;i���R=rR�׬b3���}aUQ�	F(�5����d�2:y���1�yI�0��n�(eI�U������X�Yv&��4��t;պy��"�Mat��_ ��+&q��Sd<�!A��ય͞b+h���ꛌS�L�am�yk�~�*l�<I�������m��7y��I��u+,5ێ�&A̣�N�(���_�E��v�~���EM�B�o2�n�c���̿l��sCm�_7�/Ӛ���Q,��ԫ�Y�n��i��NI"�{����+���"���PT۝Ht~A�ڥk��f5�k����J�p��O��~�s��YVv�FY0	&���^�ͧzyEh�L��D{�*�r�K[JlY"c��W�6.�#���/C=�	��#�mz+��u����:�m@>��g��ټ�G�X��1�7�yX\��O;�z��ғ]��C�&������0��g��TD�D��G�� K0i8��PP:_w���/������<$���b�f�Do[�0�Q�P0��-��o,�?���m���C��� Vu���3e����	���憻b��&��i�a�5Mu�S��B�c�M��T�~�����kq�ڔe���!��:��=�V~u)�,kW�����^2���}?�FJ���L��y�Z{1�,£��bU�jh�����?��r��J%
�f�����W�����H��"̺߱�o8���Ki�3�De(��;,���	��X`��8�f�l���:�ĮO[j7�ܕ�����u~j~N����-�rVKt�Z�́L�1g/f����L5��� 3KU����b���7��d��1���4���r<V`�=�d������>��3��Sh�ٌ��*�Tg���xm?��5�B��K��w�twg=�-��?"�gVގ���sl.��s�b[
�W��ƣ�j���?s?��'�8�ǅWyc�EL���|�N��ʓs0����<�a��Z\��z$Ds��V==U}��tDG���?r��(Cv>��b<��o{;,��n��OŦ��/?�$.�����3`�$t��j t���ku�����D�
�-��$�B%JO��Ɀnr����`�Jl'��v��+�L�)J\Ո�gBp(�ޑNݘЮ��.�N�(�l�����1>�"n��5��i\�ݼt�[8��u����,�B�%�<����3�J�����[Le�A/�+�]� ��|��K�N� 4y����c���C
���[L=ߡڔ�)9��ex���h��'�����q��]k�)�!�Ëx��9������~v�ǅH�m�ˌ�F������P���Ͼ8*�
�E� ��,J�,<����G)+H��p�T��;��Z�bVyNQ��y1�7X����}��Q3�#�n����7vEwkT�ѡ�̎��X�Ŕ��6�
���0�4^�av]�RSW�!�?+G�A����R�ZT7�s�^,��N�$S=g��uC�)|��Xk���uH�Q�97���3f��
��[�����T3�-�L(|'��U9��afR�#�N���>���a�� �c�p%e$�Hl�n�Z ��F��V�;'L:B��V2�3�8���̡��Y����<���`��n��,JF�����G��j, 
e2����� ���тyfl0_Y�;��}x�FB'Gf��3C���Ks�[��α彁�R�C��A+�W��<J�"S^������(��/��&-�ࡨZ@�3�� -,�T	ځT,�(o.a��[��J�^�Xs���j�l���t#~�g ������~�>�/�+��m-�!��弽Q�
���?q�G�te���[r����	��|���G�?�Un�# wK���1#��B�����T�n��P�������5��v+8�4�Q�R�꼭g�=���g%ݶ�a�B5d�x�3J�%�)��W�c���c�:H���	������G�iMM8p�o��ǵ�Fx�k�2R�����p���"z\r��w� ���Ɨ1�E���k2��th��옊��>J� F<)�pL��SˌRi���~YD���_�o�?���غR�g!%��=4
�W9K��k	��q�Pyk��E��9��}�!D:�V��m�y��,�y�~�'��EiY~G�^��r��?q{��.��P��X{������u�]0
�u6�C����:�Q��TA�3��̿����g!]��zȃ�͒��J�\a���{��O�k�|�'1eB:I�#��
)@|��YP}����y�ꆠW����_2�r��ﱪNq��v���P`>x�5i`��T0=��ɋH����L�Ub]��P09��$����z7�A��L쭧u�.��''Q73�6RH3c{_ȷ��8~ƶᑷ2lYf�I�Ӕ �˶�h`1tEp�J\���/??�w�"n�]�+_�^��<7�u�Zn�>e����ᬅ���廠�+z:����g"Or�u� ߔV�dtRO���Dj'�ݜ�p�j^�5����	� T#Φ�����]���l��_-t�M��E��Z�s�y,ӭyO(x-����>�o ;L�r!WBkЧi�X��Џ�W����4����P�5�����4i4�h��PR��Q�?K�\�
�o�:ӫ\ۆ�����˄ �>z��ڽ��S�v�ʙ��"�l	�@�tP�m*z��(�6ؗ��^F�飚�7}IS�#�"�a[X����up�El~7'�DO�d�x�sJ��H�����G �oc�ʉ���<h�;�d�5�uv�+��6ۇ� �,t�"4��ﴭ��r�]c'xh��z�g
u�r���8���#���x7ؘ�}IU��E��&�L7vnU����
mn$V�����h�n�O�j�Y�uQ�z�,��J���!������DM�ls���hAel�8V���ĳ&O*�m/;i��O�(}��Z��ZfxF��_wh/���quR{j�v3r���EPnK��]^y"��g�_f�^M����|A>Er�~;��x���8*�Eo�G�*����B.�l�� \�y�4T���b��j�4Fc�;	��z��S� s'��Fh�Y��)]"�Z����3m�&χ+q����A��"�p�����:V�q��Ϙ8޿�����t�p�*r�7���A~ވj
�Rx����7q��@W��K�(;D��3�
���i7��)ﾅ�!���VP�p��#�ŵ��sj�?|�O�n�9��`tjngU6㕨4�%�+K�	�M=_A+����I��q����B&�.W�e��j�um)��ӗ0�x�~�t�Ϲ�4٪9�h���'�j@x%n�M^� 
��B�qو`�q��H�>'�JH���L~.�����ܜCs�`
���N(�[���p�6x���P.&z�K$�c~��<�h���L�1>�)M�EW��&}2�,��G0�JȚ��ldO>2�ia���'@�&h�\�3�M�[נFM�*�����I6�o�~=��$�f�P'��_'�Zwiw�cq,�`���S�St��NS�wv�B�*R�گ/f�9_3����nF�����_�7��6>��S\LN-B���\����0qE��,b��"���b8�m�Tl��X��՟Rq+��M��M�p���A����o]	`
�+�c7|{T�A���'4��b.\T5��W1΁��Pn'~��=!Lx�z�xN{��g�x�=ݩ�t?�o��Ƴ[z�=���mk9x�́J2��Ů\e14Z�5mr�m|�X�@�{�Z)�eH��W��_�Q�w2�%���!,{����w�b�/���a����a)�Ȭ	��DVR���si��'��G>����p��v�G�Z:�lu�@�^��i�Z8��m��8-�?���Z��Qt���p'���� udG�*�B
W��������h �$z/�Q��gSq�����G�wP�^!R�i ���|����ًe�y+�Wԝ=�r9۾Bp3��uOH�EC����He/��^<�i���T����^�8D2�A�>��!F����}X����N�K��\bղ�?kH���QA'��t2�չO��/�=gR�K�zHnw}��&扷BW�C�dL�-]2FZ����)�_�!6y1��M)lz�ȗ�V�vV������l�r9�b3���$�Ma�}=Y�z���KQ�&��]��ИD�$,��V�>���Q���!��l1����q��%�P���(�L�sFq���4�84���d�R�x9u��&���>�dcI�H��ԑ"� 5k�vg�lȱ3�U�t�~� `d�<��˰Y�Q{�!��9��-��l;����Հ���������~u�b@�k�A ���|��9b�1y,�P�^F�66m��B���o������_w��k�󺗑#�V-m@�x\�"�@s���=~�*0�X���0?B*s(<��s�k������#<!(������ZV�J6fgX$#� {6D��io���~�s.��E�ų��Ǽm"�aH,nS�(h��r�Mԯ�_?T�Sa�X)"���C=k�(7�h9��3��І`W��\�D0+�� �#��d�����Jx�k�-�m^T6���uX��v�ͅЗ���3v��9�z��Xߙ\�T�0S2Μ �Q6roS�R��ǻN�w�!�X�%����\q2��&Cw����w���֊2?���{�/�ѨXYUz"��I�Uh���x�q�0�n#J+�H*����Z�7׸bz+�hPE����@+��r��	��;�M�?���kt��:dW��u��aO��TS9�~��Y�f��h-쀹��y��s�=	��	sJB�4�K�Fl�=ߣ�f��=�Y���n����	�)��R�45�d/e!_���JVr,���ԁc�6~�W�P<2�a�epq���J;��b2�i�aO�*�����>��Bq5�뜵�* ŁU�O�>RZ���*ٲ�(^�d��'�-�Up>��`����է=����dUWE��4	���j��8��Z�/�,R��س��$��Mu�}�Hr���}C}K�fD�������Mp���t�v2C�W��{�v�r�;0?|�l�����86��|	f��Һ,ͷ��ؙ-	��`>uw�����>ݐ����:�p�0v ;t0�̻^-s���Ʀ_�q�3�r��$��P�㴞�?��ն�j��� Jf�%� ��cI=�ˑ�������!�$�$���.�2��������݋>9�1,�gYvQ�$ yY��@�m�-s�@�_��_�F�^�/����of �_�g��,�qV�r�1�}��L|�.y5��Y0 H��$�&�G}�0�����it�����t(�I023��7v��ї�/@Rm�N�B	s�ʿ!���ȶ�Xn�F�6��CGD7�C#�B��Ŗm���F�Zda�*`k�c}�M����^��7&oJ{�Ĭќk}[���ӷ��v�4Ҩ0�z��b�O-�
���H�۰2��^�����J��=E~�0G����&�1���@N�����/��R��2���b�XAG9
�,H� ����y�jC��D4�pr�U"((2��r�_�?��f��Vt�=�jG�Q8�Y���A�0	�@8P5(վ�ԑ��gK�2N�\��E��wDXD`cc�V�&��sE	"�xbg��Ћuڐ��۩�X�V��Sӳ��n�m�1ܜ�{��#'��`G%��޼��W��p��(x���c.G�Q��t!����T��ރQ��c�3��ަ��*޴��p8���6V�n����2��jBo�-[6;	�E��.�yBH�{�<ŔX ���8d�<�vf%�t�0$��H�����x ���-'�JĢ����-�k���J�^~I/xe>��9O�.T���8��J4�8A�V/2��֐d����%�L��a������ԩ޵�GA?���ӡpF���}`�,d5;٬ �}�Ӫ �c����ʝ�ĥ���ZLH���ҧ�oe
���8v�	�_�nǬL(�W*��Zȗ�B�	;������5�p��kD1��R��g�| ��~5U���͈F�-��(2%�cR�&H�y�F�+I�����F}�2�ָm醗A��>�������O��is���w�����LU|WW����PA�D�?,N�%�y��+��)h�.|�
�u����� �qg��TP+BT=f�������YU�6��o�6l��XR����J6���o�k\v���w �dg�j� �zUk�R���i]�%OJm�ɴnU�F�]T�b�����<������L�x�<�5IX��;;�f$��޷��T1��n҆��۞8�^�Be���\0¸��C��r�+�'�4�e��%�/���v�P!i������FCe%���:����Dٻ�6$*��R:��1�c���ܰ=�	m!��^H.�Л��E���]���E>E
��1���xa����7=�� 4X:?I)���:�k�~iQTO��;�6ԝ��<iNʭ�ɦ�ĥz�o��N����/UU���[�Jޓ������5	��{Ў��z���c߭ ����(�Q�/���<i��Z���� 7�����%t9�m2�~J��N��؉%���[�٨D��f5�1���������u-�Nn*vBl�������D80��g�jکWv�,����}�Nz�⊘/G�/ AE$A��9�ۜN�\�ءS;_%�f�`���聇�!��G�����Uck��k�7�~���o�q�}�S�L�B��'��_���@��5���ma����+���(VLai���iն�_�9V���x�c�4KƓZ�j�d��DA]��wT�U�3'�>�8��@y^�����4|�W^���l/&6�����5S4#��	�V�ZTHp�LU~k��F�Zٖ�N�X��x>�%��:g����������q�Y��y��(�8��[����ޝ�n�4R7�o�y���6K����~�cc�Y�z�2K�7;���Tn%i�NK�;�Gm\SI����E���.p���f����l��(�)��k���7y���ew������qK�?��dZ�c���@���>�t~���]�W���؝EE�ן�>���(��j��&g����C�����zs<���]^闫�54��t�����b֨�b����hs9@�I�݇�y�1ɬ��1n�̜��a�a�i'r��_� ϭ��^?�Qi����3�䣾�>.��}�a�G��,Ef��Gb�[�����O���cME� �Z�r��#ۿ4+��H̚=8�Hh�i��\�+�����Ƨ�`�����gBC��i1I1<�����8-?i��[HZ\���kѦ,�V�ur�c��ʂIעMJ=�Y�����������~@��9�O-��H"bC��V��"5�<R(�y�=;���n��;�Yvl�s=B�)�M;3u/��ɒ��xS��|����T-^�@ "=��H���	dVk����2�����0�O�ݒ�nbz:'�,,�o�G���A��D�X�ޟ�	N����Y������!N�hX�`Ã�==�����8�@πb����V���c�sgGc���7A�r�:�*�6�����Λ DKVZ�}͋$ؐ� q� "MhSqfn�ź1�7qK��6^�����2��XHn�����]��� H
Ee���V��b4�s������t3�����Ub�7[�����fv9]B��mi��)�.�����2�M�5d��z۩��Vb�Q�	����R��\��: w���p�2�(;�&�m;��)��H�r<�>NG�mŖyhCZ���f�9A�v_	S�"c�5"N�o��6n.dG�(�Wj��{� ��O�Y\�j����]d�V'�)�?�,K��jlѾ7�����\5������{�]��y���>�$93*�ϗ�&Yk�|�\c:�D�א Q���"�2�v��^9����LZ�N��Wzp�~�(xx瓚��=]o�|�A���7��1hg�X�,�PX/�hfE2�$�[���8��
�H�U�-� #��#��fK/)�&�hS��>R �Yj�P�Ǩy~;�0c��gj�}d�M@��~�/��W�P騮����9.{�4����?6B�3ȈW��b����<�pA��w�dy�;[�%@�H���}�!<(�4V���h�X��/�H]]������@�X� Oh���T���'+�o�|�8̭����!�!@ ��-�Q�6�Mo�˼�}c�:��c�v��ɘ�uS���ĩ�וE�\�K�q�^d�����(�ҡ�E�BFK���S��ӛ��ң5����rlxQ���}w�
N}ΰ2X�U\G��T�myY�LJ��c^�'QQ�u��fa�����*�t˅oG9[���؀�m���V2��nI�������Zu��x�7]֥b�$��/%p�n�ɋy�(D�f�o�f�����{(�٪��x�������{K{���p�v��-�#���\�=Ѣ@|	�uU
��If�e��-��2��B��<��|�j�v���备C�����C _�ʓ1�ɴ�j�]Y�*p���ّJ��=؈툠��"�3A��g���	̜~y9KݼN���ţ��e����Ԫ��bp��xf�h�=�e�5�x[��������'�q���-�r��YX��YrFi�1�d��Á"
�ߩ�}�������� J�nZ2���mM�F��ѽ녪��WyUr�ZQ�=������9�	Q[!���r!���V8���Q���5"�DB ⵎ���yZ*'�{E��{_�-�w�H�sZQ����e�xj�,���7hyJ���DR]�o�T{��{�%JY�{G�I�aH#z�್��D��1��������'<S����MJ�6|���C���B>])��#��w�X��(@}pqω�>��m�<q��'�Ch��v;f�����^�!˅�Uz"�DD\TlhJ>�� a�W�	�JfF���
��D*i%o]ߥE�P��<^܏�0�IW����R�\��q���վ�/c�څ�,�s`��^�iBi�Q��:~�%����ږ�c�徤�����Q���r!�dbI2�<��Mgȓ,�X��J�?^2s�B��vP�h4��$D�Kv[^Z����wm`�a)���,[�:`-�:��,���֜w%�I�#1��d�;G~KO�g �������Iӳ���QK��k���׬��)x��vi�$7l��/[�J}���H^u8]1�/��7��>�W��	�zٶ@B�Y�������L��6rെ���(ؖ��L	�h�oRu��`���#z���_�.u��Zd�%V���O�^��P���b�1ڂ�����V��h�2� �F�0�9� ~+��+5��^@kjZA�4�z���d����/{>B*���nCg��,��3�9V����ds��1�
��;5���-h"aSk[z��ot��G�*b��5�w�,�78h���Δp�	w�~`�޷f���ֶGz��gc�w^)�S���w7�`F�۽��ß�V�k�s�<o\0��\W�bϭR,��O�7��%��ƦSY���ѫOٮ�&�5j��fl��z���=���6����p�;�>d��(�X�p���?]r�üXiK���9x�$�?��-�qС��4�Z�l��J�#��{�)��=��p���]җT��k�*�'���"V:�u#�`~�ы����|^Z�1d��;5���/7�SY�P�̒�?��E�I�˒G�+���7;�_�	���[x�7I�x�1��>�്.�؍FS�6)��k�S�ă_a"2͵��mN"r7��v�ȨG��d��U����j'z�E?���xk���?��B0������U!�sy�a}���j_�����;�Z�w��W+��KuAėx�@�/��V¹�Z��u�ƕ�8t�.2]ӯ\r-'���G�8?hc�Z������V�fCR�G����?�+�H"g'���d����*_�%e[��1ç�d�1���Q��b�����6>x�����ɟ���P�ż��J�޳M'�u���=�,�|�},�&�Hk$�������ո!~h�Y��U�۶H� A-|\'-��n�(��	F*��t�n3ś?h!��3�?{Gu�qb_��n0xfy��M�m���gO�q���t%�V��i��R����z#�2X��n�:d3�Q�_IDN�#}�/�2p>ɱKW�A�R�3/����q֦��F��H�o�@��u�TI�e�1"j镋��	��1����EP�V���$[��k@Ђ;E�J'�%7�08ӕ8ą�$�2OF� �!�w�.ɮ�x��i��t���㡌��0�0�%��;U�92�ޅ'�N�;��h��Y�0�p���lꕆ�0rcpK`�l}Q9O��U|�n�K*�JK��J4K�8v�/Uoނ�
,���Mcv]�蕀g'��
�c�꼏$����>B�ݿ�i��E�j����N4|M��K�u>wl�q��^:ba�q�5/A�����Os�|�x�%mz��N+겹�חd�|׷g	�#l��\	B�5!o}��,�G?��K�>J��r$�B�r�#ň��.��Ԅ���(=�4�?�g]�oL/8=+`���ٝ�j�� �EiXW+D�[n]�RH���2���:��qߵJ�gr���D�������mNb�z�G��D�zE
���� �����p_+#`�2�z�È�U����	���0[M���X�[o��I�''�d�亟�]�A^�c�'ꄍd�p
�І�Lσ��Ϡ�|�i�����4a�)�R)�OASY.�}H,i�e����K	�RN�Ւ����-sg�tW��
�VvF�Wʇ��J[������;������Y��f���w���2��/3�H�N~�'���q�!i����(��O�#�cN���d9` ��G۳�K��4|Ԅ�U�w���ae�v���7�~�>�՟6��}1l�zڜy5����|�~�?���t�����?�{RqQK�Am0�QY^��b=�/aR�ݓ��MZ���d:P'�"3v���E�t
^o�<P���@J޷̓���9w8�OB�ȹ�f��+�䁅*g�
V\~�����R.K<��GQ�B��#G7eY�	W0�!5m��q�,��}aM�į����v냷$mݴ3-��W�Sv�ӊ��%p�&��"�s<Jc�Z4F|ݑ
�{=&�/{^}���ﺁT�L?Φ��mR��]���=`�Ky���`�L{���-X�Mm�����69�̾��wyR�RT��W�ϕ��U�d��4���`�[m�Ec�ʎ�؝(*��oz�c����(���nۄ���ߧ���A���+>a�}uΟ��R�,)�!9u6�z]9�m'���\�	3�(ʏ6�ER�?�Dm��U0�f(H[%�ڠ���Ɵ|i|�0�����u�8�d�ȑ�ʏI[��x��xm*/)[��.^��Ko�l2{�C2��Jӭh+�O��6FVpf��{�&��jr}rfpX^���&|9�!A�b0h`�h�_ň�� _��G���d�)� �]��*�=<tNd�<t0(�a	�eۢ�K��w�w�{O��%�l�x˾��ˇ�Qx%����>�pe�g�����ɾn�V�?WӠ�
s�0�F���֓� �	{��UN�־=lZ�a�;J���:�أG��:��o��:}���Țo��&��s[2���_H�&��l&0o�ilG�Z�
<��:�>H����0ȗ>O�j�����0@���|����9�rC��؂�=���e���c^��3 U���K�:����=<!IY˘H��uͻU6JrG{�O�<��vvG�G�(�V����2���<����s�~�΅ß��ˍs��Xw�s_�+A��n��)��4�(����N�z��M �O�I�0�(��Br;1���O��!�0aBUp��
�&=�c�>$~�yȕ�,B�']M&9�lf�C�� .�;�j�ʟ�?�FzD�<�Et�|g�)\h��!�d��g[��bI/�m.��y�s���Yk�Ւ�1����y�Ŭ���u�����i�¸_�w��\�7�(Ƚ�.���#�dS|6ڽ$e����d�x��[��Ѯ�b�LC�ǫ��";p�ºϔ�G����l#���1Y=̨�أ��XZd�W��_�K&�^3���9%�׺f��t�㞝�1�`M/z��jg�U� �'��fR�F/�a�����A�ܳj�rء�e%�t1���mM%75J�hQ�H�u�}�M �U�'���1�r�3��,�����F�T�|�=ey9"_��_}���m1Ѯ������@`J���3m��-�M_`�����0.7U�+ H��hl�sTi���^�Y��Ak0Q�����N�I��sȰܜ�%/�~@�@Κ� ;E��MH��F�_��4+4n3��OO�(ی��3�8��*9�jŦŜ�8�5,G�]�Oe/'1����z��!��i�L@��!�p�z�`���BJ����ćP.dm�E�#¿iN�����׼W�Ku�.a^Y�;X�5׺�A�����-t5�҅�@��f��^>��d1p����l�a�X�I9s�]�k�����k+6xuȌ�O�Kowձ ���,6J��?�=,�C��f�*����=����h�Fj�ܖ��9����v.���-�`k9c[Ȣ���瀥:��U��\ki�g���M)�o����w���8����� ��-._���&ܩ��*�-f멊y��+N��>�3��:+l����]�l:Z�8��M+���{��4��_W��'�w�7]�����n��6���v��e7+��K������4��Fv$;��U(���kɥ*��ըL;P�>���@x�@�����E[+_ړ��!>,���h�Ϟ};,�ր��v^d���M����kyJ��*+qxn��w�q硥u�V
����[�~�QS�{��q	���`�����x'f��\誻YVˢ��h6�d9_�c��� �'H=5	-Zyk���U�RR�VS�YEG�H�P���QS���\�)�'�iq��7o�#�� º�Ѹ�W��$ң�#Z`�69��%��A՗����Au�=cD�٢��;�fϓ�l�)������*AC\<�rY"�}�2����.0%Tr��]�.lH�9��m�@���}��nPב�?�v���n�U[ᢧ�~�w�x���F�i!��r�#��e��S�%S}�������00�MQ��!�	*dG���Y��=w��k���!Uo&����M������W8�ʾ�=ǲ�9��^�w �.�l'D>gk�Dp��+~�}[F�jB/����S����]�6���G��{98�t��	?�}��Å�>#.�;W����S�ԝ� }�֋�� ����S�� ��Z4��~��66L��z�)���<��m�d`�Y��VRb%z���%ߗPHj��Ĺ��]�v��p�mr�vYxݼ+�A^��oEI�H��7�a��&��7
��>����8�����a)��~Ǎ�L��=]Pg��H>�zJ�\��u��+�����ouO���uK�3/�5N�Rxʟ7�������w�7��������d��]�f�k�mZ�M�$���Z;����:�*{��4�%y��&}!V�eD�~L�Lų�D�cV��.(���x*�ꚿY��!=�9����'^�Sc�C��d��:���J���)�����l�u��Ja�����Y���q�Z�{ �qF�i)#�����ޞQ�T����s+�����n*�v�W���7��sb��=�*ٯ� �-]I����U�'��3������
)w��j����ʮ��D������]H6 w �r�ҳ�dW�]����4�95${=2o;��'r�1�4��n��°aӧ�����n���F)
���!��1��@����#��G(0c���Hs��-M�:�|���WP��
��V�2���������~�Jz!`6�* l2QM��-������e�R�� ��4�ɋvG��<�愑O�4	��et����!�L��{s�j�V�Z�ȕ��݀\��,�61R:�Gh�X?-\�L�t�1��Q��Bm������E���Z:�L�����-,�_�R��h!�(`�i� �ǩ�4sYi�\GP�!D��ӛ���"*�]�V��$�Jm�!-UF6b��,�=�M؟N;�k`D���36��sw�;T�j�W�l��!�50��f��P���1 }�[�ٯE��o��k;f��$C�6�b䮮�w��eE�	���`��E��[f��e��Q�Y4��Ozx@$~��Di��U	Z��o4*� �T���?X�T-�R������ή�뭚4ɿ�����`�*��+:��0�V+̃�����,����fz%I��C�N���'X�jc����U>���y�[��Y�=k|���N"�B9N-*CI��C��]$�,e!-ѱٟ���},3�3D�"-7��p�o�IO����J�-rgF�b�c-���|�?���NKw2����6���.��^���G�Cx�M�X�Y?Y;�3w���NxՁ8y�z��y������d����ث�w}g��Hʑ+t�c�mi����J�m"�P_��;+����гj�l���z	�rV�e�v��՟0H�G���{��ؼ�ɻ�\�ǳ�x��h�0~���,W�&pN�$ى�G�V1�n�6DLcC��N}�&���飌����[���]��2����W�}b�-�i�.��x;�J[F���Ɋj�5ی2	@����ᣗ�%�s�{���,_K�ۧ���n��yAn�b�~�.��K�y6�j�ghϤ.�JH�f��voF"���[U�n�{lf�� ��6�m�2Ȓ�]TbAG7k�/<-�>�)��jh�-�����(�����S�7·��z_��;�E�E3N]3uxR���n��>qe륌HM�m���^�/�H�\�؄,��=���� Hw=m��U0��Y��u�h�Z��īa�e����@��a����L�X�4�[I�Br�����8�+̃ٸ����Or^�}w$��_���!���B��j������5��maH�����T�������f�BU'X��Y%������M�Y�7 04��-��vk�F�W�،��[����ݛ��_�^ �J����f��]���j�$B�Lf/u��G�o��[��}��)��@�bS�;m��l��ʚM���FF��z�8�w����聁��/+�V��H���x�{��jLN��2��b��.@���,�e�wdd��K����Oٱ�CD�g���e�����KE�g�x�*~Pl�1�$�4K>z��u�
��q6�lZE8���9���[-=M��d!��7Ş�lRVYM��� ϗ�"���.�xhy}4o /�����b�8"�åw��,K?�8�*��i�L\Q������� ,gh�S�e��Wgx��W������^�mK�q ��֩6��\A�7xx[��m?��a3�c�,�-�����dR�\_L��9E�Y�*^�lO�������n�R�m���l¿��!�6%��s���I&�}���P��i��ŪI�<C(j��c�۠!M���q��_?�5Xa������ۇ�ɍ�﨣����Lh�LR#-��]��W�u���aU;���'0��J'��VC-��a̶����vY?5n��B�䷷������z�ZH�1 .k�I���>�k8
Ճ�>t�gw|�j\�Wk8��R[�� /�f��L*��IW��!9SC��:םu�<i	�"9* 1惂����5��h��R ��w^�S���mPgz:����@����� ��{�B�zh�.&�)vNܭ��w�B^��K_��@#��ސ�yI���N�"b����E��i�#�T,��b��:|݄���'�)g��ٌ�gc���B��� yxCeh�1������L���ݷ��c�h���-�#4��d���oU�����q��(��Ad���e��b�ה �9���v�p��G�r���ҕ*���X�̗\�'����:`�4���	��镂��V�f����{i����U��ե�F,��y���Y�S�4�A���9וX�"��O���:���Բ�;nD�9&�����_J��hQ}���Ν���GЮr�.�뎙=`^j��r�ŗ���,�Q��Wnt�a؅�bM��6�3N��o�W�-�z_�*�	-��D1D������겿�^���ZV�:^�e�/��߄]�̞�I���.�SYq*�܁HR/ŴI_�t�?��
}�)���Z��E��Z{x�p`����k���8K��������q!����FbP�alb`q����kp� ��ټ�x�5�'w����Q��<�h&i�����>*�Լ���T(ս!_;?������߸zN�X|���J�U� *E�M���3���U�7�%��D��pP�����p�kG�:�|�Y]k6ɼ������8������fڮm$�F|�Ҳ����g�3������9�[��վ�s��q7a���Q'��B[�9ٴ�5��HI�e�"�>���`�{�e�$GW��y��&;hEН����aJ��{;\� �oY�q=�>i`��d�
��@c�
+�Qa�%2�D�0�j}��P��,舘��xH�<y\s�A%5����k9E�0��������<|7��2QR���Lz+����ҟ�ڗM� 8�V���wƥ8�~��P"�A����7�0��)��X:t>�o>Uŷ�f�{i���X��N�aYE���Z�Vƿ���Z�b���|�}�D����g��@�)�<���Yb��I�-O2��}M�c���1vG�Z������^I�F-Y�V"(*�'@�g�/����_�sŏ�0@,b����̖)��MB	(9��]1���v*y'�5+]\d��}�B��l���(t�)_y>��X[)"�N}>i�K�آp�U��w�o�j��׈\W�o��9���ט�͊�^֮$;<��Nj�"�0VT��$*���̣�'6q���aLi�Ό�U��	����eF�߷���ܣ��c,�0f��~�{P$�5;s���_�����rC�;f.PRc2�J����5-��0��+�@m_����*�x�í�E� ����>>ku�u�!辚�e�����@�]#����,�u����_1��f昨y���b�Ši�-QH��Fa@���2�3�H�G��͐#N]HE����(���ou2�A���6�>O��ǜ-A��k1�D��P]!�h���q�0���΂�o�j0�E��pV�hnޢ)�V���]�u��
��w���B��TI���& h�CbT�����u,��HB�|�t�a6Y2��m7I�(�{֪5���Ņ������B����=v�*T��eis���q����o�HEjN��"���'��^W�>4�' �`�T��N���^�j�{�q��9���ˤ"_2�[�*�%+�K�a/�>�Z7C�	����y��g�gˋ�Yo$~f~}TW�%� ��>�Av�)"{�!fU �h��/5��O 8���⿪M`+���=Z��{*�y #۬��V��dh�Cd�R�EL_B1uP�O��<!����]K�C�����
z�8�¡{��:��<��6�+�e59����$���YW�IY�8tT��P���ow�����I��o��1w�*�<jN^�Wm�<m"���!�j��(��L@�	�ݹ
����-��4�T�GV��x��RT0S�z�n�U���,�	m���^\-uYx��Z���ͬ���6�Z�7�=t��f`��$�h�>9���'�0j��RLr+���S|�n(����?��1�I���"��4������Y�d:9���Ee�S�8��Bƪ��@�m�B���>�oC[?&s
���s���۰m���A���u���n0���h-���k�}�0/�w0�zkL<�8�q��a���CPrΊ4Ie�?.�Ma�e�-��}<���҂2��ҍ�ԹǨ6����2I'v9h I]s�1bi���ә%'���Q$�}%�å��XLu����P �x�J���
�`���~H4b>��Oc�����\V�Tw�*��6m����nƿv(ά�+t�3�_O �%וS,F�8r��*�_H������s���G\�D�9`\	k��2f��k���F�x<�H�L�x��f�]ߺ�Պ,_���>�`��Py�zg� �E�TΎ�w���M�e�%B�F܈���DXLְ�ХUF��AFP�H�����>��ObU$(l��?ˆ���u@tr�^�Y<2_̕d�m�X�O˾��]z��m@/���fjT��2X� Q��~#o[?^"u���0p��e���&�����ԙn��2� ��(��4�㗞H���3�1L�mf`�DbE	���G�[���<tE"��[��W� ����3����~��P|�k����(�c8:���rONy����1e�ﾁ��(����y�j�^�J�� �X�vq"�J�����N�C��M��JY��tS��C��j�5��_���9�V)�a�v�)��E��)��.m|��T6Cc����7F7O���%E'A!�EϞ�x�j��i�@̮یC�,F�i��3d.z����
�ч���Y�7�f��S>s��S�3&��Jke�im��Ƚ��G����;g���,�;|������"�� �f���H��NxԐr&�C� x;U�i*E/����iU6��	=��W�^�J�W#�����ٰ���Y��ᶬG��!��p�{W?��Ϯ�
�� ț�IY6A�tϬ������V��7�Mm�5A�U��+�(P�n�z�z!�=���恐I�Y,͜�8e��ӊW���uYz����W��&"��:E�8�)�����O��!7(�+�:͍�=�Q��ߋ�@B�E(p�;>*��
�@�LVG�1M���ck�[�l�r\���p!����?,G�\���[�*����	�5�M�������&�Ɖr�dԑ'
�B.|����8��	�D��b+\��#�0�^����=��Ӹc�0�7��a��Ţ��-�+����M�,�ه0EU_�t7�4Kr��������#�$돎gkA~"��ɹ�Z&��PK)aDaW%��m��� �E�0��gT���yNM�|�p���$CΠfHE�5^-�}[��cL��N@�u��Y~�1�LL�O��g�M61W�`$+59<ǶWs���5Y���4�ƕꬿ?�)c��v�����eJ%�(9�3�}9��Nt�ȱ��C��}�����׫�ˠ�mЇ�G�/��։���w���6?2�%��J�'vpk �?�O�V��jñ���mY6�F�������􀐹4z�|��h[�p��ۯI��Y~5�S���&�bmā�a̕�gEݰ�t�ch(�${sF{���K]��{��c�(ѭd �����wF��p]s��"�g�����ۢH��E�A ӪO���2��ܜnN[=��v�1t�@O�Q�r�t���Y���b�
�{?����ȋ,�����A�y�Ě62�`i�S^`�?����UFi�uஸ��h�9�~��$��w�=i�AYᲲ╉L�&�ܼ��������h���P��qJ��t�P
���#��N�'�g�H��k
'�4����a�
�[�"�R]�/��$ u�ۚ��N
�t�"�ڷW�w�� �#�����+�
�-"q*��b��ᚣ�����q�9�	'��h�_���sg�U�,;,�40p���]���2��H���ߏ-o�t��mR�c*C���y�0��[��
�M4�q�6,���%�wp��4��FA�(~m���}w�%I�]I�r���~���F��q��Z|F���ڝ¦������Z"Ԓa����+��S�����5=5��!������rt�Jm����Ą6kC�����:.��%��rR�W��e��[C>��~�'@�Z�eN��Me�J�#�K��Ր bW �B���9A�iMZa���ǐM�>�|���a��S�&��b��b$
8'�����N����(�
'�J��P�c1��o�#xg�Nn+v�śf9�ڇP��;w�H�I2�e�4d3��w08&G�d�����	勝dcg����*f��"	���"�]��7��.��=ԧ~�T�e(�BRZ~Τ����E�{���k0��������#KL��/L�Pv�O����k�����L���N�H��ڷ�����ﰗ�#RDv�c��S,k6!ѨK�*>�jw_��7v_�Pvo�J�5��������0|YÒ�.���lx_�f"a���*�5	(Œ�F��������*�@�����2��Ao���:���ur�{�h�eb��]�+��Q-+Qc��ܵx-��ٴ�J�'ֺ��
�, jk36v�������䔍*�y1A�Z��@o</]Jʪ|���ҡkh�8Y����gx���f7��~�n�Xy��i2s���7�}n/����h���Ix))�|i���J���EN�f��>Gh��!���iu��)'?ֿd(�h�O#�����Z$�V0桧��+�0w�8�X������e%j�'��Ķ���`
X4#�Ɏ@֌�Y���1�(�Z�{�Tނ�eަቘ�;�����1�[�G��c{����u�R.1�R'�$�R�*2���iG�������؃�9b�t�82���壌jb�NL��$u<k1P/�}�H��,�p5��Bh��[ �.��k!K�4��L ��"4O�9FŎ��۔[e��#�r����& k�ZiD\��:����s��5e+�E�����Б�r[`�fҲ?��(G[�
�*�NR��B�|6�hc9~x��@p�D��e��W�$E����Qj��ݷBJ�g�~��欉��΋�"�*�},HپW�1��&�xPI��OЌ"�$��u������ϳ��x�8pa}�;x�\'�ʪ��?&���[i�3�$�,�|$�p� ��5�Ӕr#��M�@΄��s���\���َ��"��3��W0v<��Y87 �Mz\c�4���~ag�����:n���Lܽ5)��f�I�-6�0E�{��k����a^R��U�*�%g�0ㅟ?�w����?;7��Kȇ��m�5�Mt��|���Ot@�b�<m�VU�-\n�rVBV߶��IL�l	ͬ<��������ƨ́ϓ��E૯��0���W��\�H�]����NOF��L󌝮��V�#�slV7^�z$�}e?��K`��Ua�ݷ����~Υ�DdZ��w���`���f?��Mtd�t�cW<E������S�0�cYƠ����!��J�ܮ�~c�����w]#�41C~��i������R�HynK��E�r� #[�Eæo�>�rSJ��#p�Zũ�WK���'D�V��A��k�H�LA(UV+��;$�fEK�? �c,�|6�E�)������5��X���|�����{��X�p�-�'�p�����.�+�{��h��s��댕�b���R��w5J�"|�4F��>�x��T�ađd���=,?\�&�.�p�#+�����@^i�-���$��`�J����S9��$�<*$�tz�
�
i\����WhZޗ���p㯲a��R�Iqd���۹�X@ �h�c��A��:�bT �SN�r�`r+:б)+X�����*��EjՐ��{(xuq��Y^ܧ�!C�PE.���$�l@�	���N�mܙ����i�l�s�	Z\���|U�X���K�5��V��_�m�}u敊.n��>�:�ի��H��B��e��C���O����3�0.�UE-�5�{�-6��-39�؉��^ۗ�r�=��>�eq9��ڹ�J����D��
�tުi\���"�@8ajn���\(V�	��^]�EΆ�Ga���ɸY(?:g��֪�"�Dߵ��̗տ�˸�����})"�e� e�a�w�� TW���0�\ߴJ��*b�_C��1h\
�����"/�S�Ê������Y2aQS����_I�	=��lO_w�����݇1>0�T�O]��5Zӻ�Ą`6ک��V�'�>�=��҈R�*9�pW8�d�8cC
L��I�t�?޷���j��]RDo�R�0uČ�]��]4ŧ:*�#�J5����5�=�|�_����h"@���/ki3�I�lӜ����Z�W|�g��
-��]�&��0-eR�OZ��O���Yn���n�9{q7�<z�򏼃c��*kN���%�V�Q��2���Z�8 @*��F�*c�PH�e��R:���B�I،h7u>l��ȣ��-�݉�J����V�C Q�'@��+M����H�@�y�g����S������YjT��6��i<fS�I7|!�k�\����boBR����W4TzFr}�^��j�L�Bq��T�k;ۯםf�VP^'TN�����?ܷ�6p��B!��؅~;H���F�"��>���pf�����TT̲��0�v-R�l,�#E6_����M� >���b�n���J�ҋd\�:1x-��#���xʇ�J��x/ �N<YqMn�y�cw{�%���Y���eW�M-����l��-����|�@�(��l`� ^��,}��0�����Y1��y6�q���z���L\%��4|+C�����?�{�Ca<�_�x(�a	�?�;B���Jڐ���/ɨ��>���@��ը������D3*�X�o}�@����d�7HF-|����a�[J	u�E���#���+��|���,m�׸�/��9��G�EZnT�.8��@�#�i
Wޭ���Zu~��W/ő�]Ҽ�wa�/4i-�X4�M�_���8��U}M�%Q�%�H�\6y��n�w�#@m�I�	���k�l�h=�Kw�Y���~��cT��I�j'�=�j�	3�c���=݈�Nz+��W>�EJ��c!��[ANL�S�!��^b��Dd�z��F͘�u����:!��L7-���A�9I�H6��0�[�2֋�a=^�;`��QO�&8i��Pg�❧�:<?�k��c����To׆�=c�ө �p��^$�G	@��<`��2y1�Gj���}���#L��d1�&��S�q��B
<�:�I�?șβ	UL/>kᑑ��XZ8�m��]O:���["��j�X.J�������f}��O��\��R24'�s40����B&�˱��7��/=~y^�/�HT~�"��z�m���g�.�P��4��rC?�DL������Q����c-�3ƻ�/�6��_	������-�3S{�	��9�7O?��,��ܬ�ÎF�#K��3.�h���c����&�(gN2�c�P�xl�$���s`��~��^��97��^�3�X�X��jBbe=X�+�Ί0'�ub�O{�|�mA��MX?c��G�j60�����}�EZ@ʪ~3��P���r����Zˑ�5(��#h�aZN����rЊ�j{`F�6�,u�DNn���up䲊(�d
�:���-�,#�W�by2����t�ݹш
yD>�=3q$�yK����4�Y�F�4��L�&��J1ȁ�'W~�p1�3�r��d���]��*�G�&��RI��
3�,+��Ϫ�ůZ�;N:������̝���u�MH'J��GF�Ɠ��P��V�c�uhXFK'L|c�n���g����G���:�.^P��}:Q��[�A�W\�-\Q��-͟�Y*�����~����0@K��]&���)*W#�UE����D��¦ԂXђ'b�d{�'�m���0l=����m�VX�}|�Γd6�L
�J��E�Гz˷�=����yD.�P���E��!:�/��k��o�Ҧ�m�1�$�,:&Ț|̠�j���dp%<��zP��b۠oF�&�a�)E�)%-��C~�$�2�F�j�v��DeE�j���kB�����@�K����ZJ�k	�"��a�Sc�#`i2h�L�h��E������7vi��g��ę���K���	���e�l�71�f@���,	�]��V����<�� �n�7�2SB��$�dd@���r�5�>6��3���v�8J�{��V���V"DR$?K��y�+�G�b�����8"���������&r2�|�0m 㬅o�]Q�'{�L\RT<q���Ƥ*ZMZ��H��*�-��d^�m��ן'6�T����fL��9�W�;�����)_�Ǎ���0�	H՟��;X��	�i���"	'r�<rf�,��H��~��1޽nC���fʑ�;^�X���
�N���$�Jl�_�%�9-jQjؿ~��(=��i�2�SF�.騡����%��@Q��z�CH6�"7AF�R[υ�~�ZN������g�l�*n��T������]a�ӽz���j�4OM���Z1��X�Ԍ�������`�/U���$?۞}ã�����G�g�7:�Btｇ�Sr�5��%��v�c�Y��X0q���(]�_ Ih�'�.w)0�d&�YZ�4�^5�����T�#��I�L�"�� �;3��$��CDt� �jo�*�Wn�/��m舔=�DL�~���jBĸ�'y�Y��C2.�X�����.��NM��h�͒J�\0�\K�vH�9b`.x�Q��`nV��zn��1������a�ٍjS��ͤr�� /6����#sڇs;�����e<��׃ժ΢?)�n�����t$s��k5F ���&������
x�~����2 �����z�X�>H��i���ԙ��L��V@V�-�mp�J�?\����K�Pjw)BC��q���}�;A�V�2;f�$�V�'����b�����,���NZų��wͦ��eq$�Y�-��꺨Y��שyT���I�uY18�5��k@p�E>�c�.�N���=�n�q�&:���EJ�5"Ɋ0R�I����o�7&,�k��W�P�:kDգ��㏠�ڧId~���a��	���u��]�I��0@�����+?]weX��@4�C��¸����Xc�>\���uKu�@\�'>�j�Z��p��h�n3��na�y%&~���� ��M>e�������ц���/4�����)7|�mM�Y5��|㊸xi��:7�H�qJ)O���z��Uٗ����LY��(��Z����䪡�ᢨR�4?����[�Q�tG�3A}E���R�*���2�[f���MV˃��\@>��V�̝3q�J5��hf�V�3�~x�ôʬ	�����b��cv��,��Q�H����\����P�� ���������^��H@UМl��/�.�~tJ�\:�2�nSC9@4V�Ұ�u�� �8jgv��62�[\@�X���Lj�b9TA��G�iJ�_��AR��������ǼFm6� D,�-@��;��m�u�}��-SK����X�A3An~m�z�׿�2莈��~�֜y� ���2L���⯺D*�)ny[��c9�a�	 m�&=���js��Tx�Z$-���>�>)���lE�K\o@�S�.c�sI�2)κ8�K�[H�`a�]%E�򧸲j�5V��ޓ"�I���d'7�s	ER�Q�6�ˢw������l����Z6����ӂ�#�6���oʩL+*r]dOͰ�1������g�1���o���X�b`���/��πb/^ퟴ����`Q�e�k����'�Z*��%d�;�%�G�m������Lt�6XO��c�)Nx$�%��J��5�h:����&�#�rrr�=�NXB`r�!L��3�	o��):�IY�3gQ�D�)�w�Y�!�g-� S(�z��W�r�~U�o�p��@�������2��	`��1�d��V?(�f�\��O�Ͱ:�)J�(�L�<�BT�fnI��N�7�Jɷ<0͸�uO�&cc����RVx�k���[N)���H�,�<�x-�0�m&e[4VG��i.�����q�?�s!Eu�gu�4�NH���ȁ?��f|��~ׅ��HY��΄�a�Bg�zw"�tbQz}ل�߾�y��D?�"�|A�Ԝ�ͤpM�8�qӑ�4�7\�Wv��Y�]��q�@${%��Z�L�:q�9q�����
?�ܘ������D`��鷖�W	��q�b��K�k+'f�'�������'AA��_����Գ`���|[sȢ�"kj����93�8�ֆ��Mz邒�$bs��r֢�1!�ECV̠Z|�^f�K��ͬ�b���?�ζ��� 0�<�%��3-e���x��l��ެ����b�(�h��Qf�!Q^����3�����z�;�.�� C�i�oM���<<��|��$�F�H,��|�f[S��-�%��`�l��t&�o��(��^	iYv+)��$_����A[���bM/~�o��ө�b�/�d��#�t�{��\G"��{U*t~0\ώo�+O��Υ�� �[����	v>=p늹}o�������Tq,/�d�C�d��Ve��ns�dz[F�F@�jS�k"�_�ICH ��o��ض����9�T#ީű��0!	���\�s�r$1�*�nk+Z��}|��C�EςY�9 ^���-ˢO�+v���)z���S�E6�Ҥ�	-�y��[�Ϩ�=�$���[T]YB
Z���Z�>�_����s�iQ����W��j�K=(г��B/��t����*��]��'K0�ˇ���`0�"O�j��󪙾e���a+���)o��M�k[�w=S��etK[@ȗ��F��V8n�N�6�[���P���}ju�����-�����尊�?w�jZ&Eӎ+��Ay���@�fi����P��]z]nFH�NNa'�m0�L��� �ܠ���d���q�IľCV�9ZMX�[	��{�l����~�0�O)|,v�����I[�dd�P���AX
r*�%��n�'����9E�y�ƙ��X�N�@�����z
�G���*g���N�z��qښ#��0d��N�;�Y����������&Kr�џ�:�ќ��Q��w�����幯ĥ�<�E(�$%iO���5|=6\z� ��6/�����Ue6���N���$N>��jcKZ�K�4;-��e������>�f��ϲ�3�7 %�7�Ud�f����O�paQ�e�s�ژng��O�҃sQ|6�5�$��Z���	@>\���'�|^N꯬�\�sSJJ�'7�hr�lH/R�Q�r�'Ĩ�g��_t��ŅŞagȒ~ds�w�X��Fxj��B~���%H��`m��de�w�̨L�g�hf�q]�Xo���:��z��_����i��0'��qiY�[�!�>P(A�b�𪀉�D��ͼɣ���Y�v(@!�YE��~���$0����V�G���9��a��@ ɸW�:g�� �nv��5ʧ}*�.�A�!
|����5�)���^���3I=�z�nQZG�%�K-�[A�J��;�N�/r"�~���p� ڈ{��#���w$���*�o�Ͳ�Yn~p��Y������g+@��ga�a"���{4\�u��@m�pi�.��y蕏|��p��1W+e����f1!�VPd�pcEQ_�����X�K�^g5 ��ӕa9ʱ�(��֡x��&
�� o����+v펫cm���j}5����)�� ���	�����x��&S��0���v(��A4"tA��%������[-V�<�B@)�N��\/��:����J��љ�y�&Q�	��\��4�^���b�u�G]�pZ?��=5��M���-b�]��]�ο/R�Kx}VS��f3���W�17�P��{pFQ����~x>:#�6�#�c��t�>�L����1���:�q�T.L+IA����yB!Ls͘X�~�A<��p&4�_^�+�W��ˑ���j��&�0���G�gف����4?i����G��@}��|1;���w�8����W��{k�0]B;�Yi]���1~��e"�<9�v��r�nz��-qww3?��/�e^�ⶳ֦4��Tꗻ�NuŦl�@$��x`���ZH�O�8�s��u{&0��C��AM�����G`= k,��	|[֦�h��=���x���H�����c��
��l/�3�PZaI�����pq�?�J.��k�,9�9���à�f\�_i>f:�u��L[T��9�a�̪�gQ��\���{�7l���G&
��3�*ϑ��r��v<�F�%������fa���x��3&�[}�k��|2Hj5�F�b��Fq��A�s9&k�L�����`�0����H����Ɨ!�?�Z6�(a>�:�@ݬ {W�sm9Ơ��XX�6�ȠH�T0��h�n����W_T�ABn%��^�&� ���d������ zz��9�g�� :w�1B�{]Fu���T.��uW c�	��ia�=������}�h�>�a��/#ѕLI4��BM���O��b�ଟ+H�n��|���c]?�ɠu��[�ۊ�D��O�/�[΋A�GMs��C���n�M#��4�T�����	�w���C�� E')���Yu�ҠB
]J��4<�����e//�wߐ�J��U7g������9����.�%+K�����Ņ�C�qDp��2<"y�.R��9���Hs:�T��j�@��f�v����c������_v�h��1�(
�T$]Ne)]�e���c����q�B<+��H��|\RI�3��m9�&�}�Ld��wj�/��,�uHy��-���8��߃���������5+�~^�֎Xm������W��� �x��Di~��Q6�ER}����`��*�^���J��>ݬ�u�sZc�p�rqTvGJ���5�K��}���Zv��n���S�Q`E�'�ȼ�K�lLO3>��	����n�z��τ�fW��p7��ͩt�$�Y��l0/J3��6��۷z�P����]�v%&4�%A�8������}1=�~]�$�"����d�w���m�}��D�X�#3�^�H�P�����FY�$p��x�dMB~/��V	Ҭ��̹��oGk��b`��&.�"9�ظ�h��W ^��y1������8��Ӡ�u�ǹ��	)�Vu���	�ߖ�H��;)=��h82�iϙ���wh#<G�ظ�Y�;9�T�O8'|��C�H���pv����Ь��������i�u�?�3�N�5{?�s.E��KN��
G��a?u7{5
�"�
�;�˗�m��m�p^�Q�����>�l���}ұ\7r�X)ɈM��V�����aű������9ݘ(r�����]&r8�y��M��.9��*�`�T�*�����U��W�srE>F/��b����+Gj�J�L�/���P�i�9�	�Њ�U��q=�&Q������Δ��R�;����,�SK��o1��P�/	S��vHNCwE��
�&�vBk�gO��k�ϯ}�1��6�]����X�[�p�ƃ��h�
�03���A��/�M�5L�%��[�\�k��~m���B�G W���G*���?&���!�/yg����C��qJ�ȑOM ��#U��/H���Ʈ���o��>[a%k��NL�q���Cy�h���l�Y?��f�c�:��EbJ�ၓ�f�
D=��.m����%ȍ�tH���¶��yܮ(	�q���>��0�+�r��El�dS5�����i:�����?�vx�S���	Ǟ�:��	��&S��J�D����X�0����e�Rv�0��KO�6W���N�ܱ~İ+V�QlH����9t	���$.l��6��x@�v
�����]����ֻ�rq���h�����m9)�!PcHI�d~�u��x�����TZYE��&��'3�t���!f�Rd�n�ͳ�{޹�*-�:�Ԉ���MY{	P�a��ߘx{ӊ5�%W���E�Y�i"�D ��"iZJ��Γ��CL>�j|��[��k	Q��)@��bhB��1W�{
:[�SK�(F�K��`1ӠI4�+�7ˍ��Ƽ��\��Q�Q�Q��^3&"y|�Mc��VG<W�a��x^�^����i����ϐ�$��˘Wʰ 
.�ȕ�=4$��\��&Ʊ���Al"ݚu����Sr[8\V�P!��Y�����8�.XJ�!�Ԭ(�Ķ#q�ǩ+B��a)$@�ߎ����p��F��ҜR6�������e����쟨w��n��f�U:Zۭ�P:���鍶uW�����������f�л}����Yr� 2�OL�v�n=}5j�ZIo�I@M�@������PӚ�ƣ쪗��P�;
�Un���^��.�z�v聲�6gv6�W����&��7��޼,�9!,�1%ɤSY�|�'�:jW��8Jۢ~��%?��N�4�"a����d � ��\�s��J���Cɛ��;��|Mk�ľ��l����m>A8պ��
d�Ma�]4�<,]AMy��m��x�.O�"v�^�����'��)�� �ag�^�;�p��='� �/�S�5g�vy|�7�.�ؾ'_��7�\Q��Z��h[&��pU�!��O�`8�� ��!��E$�ZR(��iI�� ��S��B���ޓ����*��
8�%|k׷�y���U�`9���ξ�?�����Uw�!��EgC��7:Qh�!垀7g%˃f��b�������˱���@m��K%�?R�t�;�i44?����0�|%�?ɑ֨br�� mb��1�ðO+"a�<p�z�7��^ %�3�~|�kiM,`u�	j��������2�ؐ[GW��p	o�R5��Z6>4A�	���G7Ht����K)q��N��a�6=M�|WǑ����(�K܁)���gߴ��`U���ພW�c=By�	��]>��R����k;W�*��sI4�C�\E ѹ7����CX���X��\�>�I��m\04�Z�$3w���6��|���y¹��gC]ՠd��e���/�Ay]�EER���-�z��N���N\�1�5YR���H��hs�i�1o1嚦�A���=�K��pIBf��u����}��(���hrc�Ϙ���@�vƬ����ߣe�ޜ���,^����@�G%6��K��gO��f.�V�����+Yd��/�m�w�M�x�Z7a���@/c���qT�Z�o*=�J݀����

�h�����\k��j��0n�'���E=�����2��9l�'�dR��h?�:_)YT��-��:R�ډ}�-�T���J�щ��%�#��I+��xe��O�u�h /�v�P���>�\��
�T3���%ͻ��uUh���$��լ��`��-�\�x̩�+Y�J��[!C�?E�P�Dͻ�&�A.h2��|��L��|��f�:Ul~倮������`��7�nn�p�HGj�(Z��\�9��t[>�	d�p� C�S�j��^�d�f��,�r�z&F��o�~Hܦ`T�9b��h��(r�f+�����h���⫵E���).���.؏�U�o�Ż&��P�5�~�D��;�Mn y���~> �3L˩8�C�	0�g��.��x_;�Am���%P���<�t�U�7T\u��iӬ֩p�Uǯ�cJ2Xq-�.\��Mt��0��D�m�twM�go��Ϻ��_nT�3_�*�願J[��'�A[��-�K�x�Z����w�Yy��$���9P�Cӝ�o��xV�F��y��	�����"K�x��Ո���q1�AY��_h��k�	ǩΈT��j�_��`:��^�A�G�:�OV2���t�ǘ�U��Q����k�3l�+t �W�XQ˶Lԡ�47h�O@/׻�q�]~��ݰ:"�@%�u]��ڋ!���F���B�V�X�U'�;�j}��h%3A]��+ R~�L������jAapw����<o1�,f�5�B��Y�D�+��]��{A��T���M����}~륣��jŅ���?�w_2�H�	�/�N^�b/��f���[+��?n������7���.M˖�a(��h'b�GP��:7���c�2Y�Fu��ɇ#� ���:�Q�M7��Z�� :*[>�K�g=8V�V�����
㲷�4���Ɠ4{ٺ���d�p�^?���f��J$�Е�*��(�7�߸G<����$���ۆ��X�5en����R���;J/
*m��`�e�'2(�1��e�!u�I��1rh&!g!U�}	>Q�-�{�,���	�	7�5_�b��S͎���-8V���%�y<36��p@'dc�����	�u�{�rN?l�K�Hc���ȔE
���/A��hO�ʗ挫�>��5�c���@]:���:9F5ta��o/�8HJT�OAz	xP�D�ˆJr��4u}5?y{��_3Lt�[�&����/�}��T�]�q|y�q,��p�մ򔖭��|{ �T���+ ~����|�l���fF��)\������?�}���R+cf2��'��\�������U	�!��Yl}?�}ջ�8�g��ӥJ"�,������p�7��D��8��^p\L�˾w<��A?8�"a�����n��?R	G��{�	��%Ĩ���� �	L�ݦ"n�`R�.�<@} �Q	�p!��t∪e��2�	i�b�\�<吐kZ0ɛ�;�:D�I�h�� `�?�e��c���@4�<7!�'1�ѳ]��@k�DCxl��2�������y��͌��(�!tm��b-���N��.B�f)E�Ƹ�Ď(�n�~�}#���x�3^�aO/婁�Y�X�լ���`�D��/;E>ƞ�2���'%y�L�8 ,kP.X��{O�E��X.V�$�f��zom(~_6�y"�in�8RZ
���z�C�OP^��x�1KԸ���2�m��k�_ۼ��*F�#��2�������;ÿߗ�J�V�±|�-�:��մ{5s�s5K��Vg�W=h����R��J�`ҥ��Xk�fѥ7�����Y�Qg���,�)�D�
 ]��h^rHn��h����~r���CWߩ���h%���+�/�t���'U���*���;����˜a��6nU}W۞j~�i��o�2V����
�����SOϾ�X��"�e�c�$_��w���3��^�[��0]�Y H�1r��	zא�Eu�����O<��� [��~�kxn#CfC!j��ZbQ�cN�Y潊Ͳ�ѓ�kT(R������:�,����v�eJ	�3�~�Va�� z�����Β) ����a����0�uj'Ϸ��M�f�Yu�"�k'��l��8�Q,ҕW��%H���Dv���wp��u`b�G����YUE��%�X��zϸ�ҁW~�2 s�4f;�lF=�$�{��z1�3�J�|���g}�0���M����}��w:����ܴ���%�����_�SM��S����V���5��Zy�D���X�:t� �%Pb�n�ոU�)���+^j��jA񎔫���\��I!T�(.����d_��Y���}g]n���~�xר�D��^�r��s5S�Ә2h�/��ma�L�󔌑��ϙ����0�Kp�����7��=d8����^C���lIT��%��M�ȭ!����7P�����AM�m�dQ�:Vd�%E����@����K�~��?F��p�4j��F-=H��E�
�s�6����K�ᗿ�}������ �&����)}x������%��4ȸЊ�x��
���I�����_ ����p��o�i|����?��ޙ���%0OMf칱� �n������P[}h����3�vp�G|4}u2����P�Û�gh�#KRG��!-�pY1�w�<��aM�Q�1��d����X�+�?qv=��(�
�8��Q2���丰"��B�����)�M� ��㨁9�?8t��`�b6.����#>�8�N1k���Z��#J�e���B�n�� v�-?����gJx	�b��K|�	*[�qiV}��܎)�{�A�H�`���|^j��nӗ_n��Xl,öx^k2�򧋻G��1#/=	�!se�W�aY/�D5���kJ�u�1������͗S�'H��*��֪/D�OvY�.��jF6*��������z`P�Pa�yL��
�^ �7�DD�f4���
�����`� 5!,L2%ED����}��D=��fa��"����gp�F���Ҹ���e���S~�gd��r�̵����
0�lF[��]iz<\�	A���Z%h!<S&��!��`��������`UGos?�y�k����� PjA�_�}�0{.���s��R���������]�_Śq���Վ�Wɕ2��[+[�N݇������}�Nbye�ǝ����J�i���~������Lq��?pw�:dQ(��9�eɾ{Gv1��H��R)z)�И,�����v�Jk��LYo��x_ɝ�r3�KFB�6b����6� ���î%<:����[�,jN&��&����;�^���#���e�Z�N6Þ�3��h�S���e= �qn�VsS@(�}s���Q	TP�r��#e;x�?�:�xi��|�h�ތu�}�����]_a
V��Mu5~���e6�������'�uԹf���Cpт��)t.
��[뭚��	|�x��&�]z���DX�����ڈT[�mF21�mwI娓�`�QW��)w�bQ��H����{�M�!<o�O�L,��ǳv���pY�B�U����U5�U��Y[4ˡ�W3^#3i���u��=��*�0-�-���w~�^۝jE���!r8�g�S�:x80�]D��uѲ���.��4y��W���E
z��J]�����R��������mG*^l��,S(B�$h�PS�� C�q`�R�W}�L���.� ��<7?h��Όʵh]�h��jI�8�J�+�B�r�\��,���g��s���CѦ[v�iU��So�J�1�[b�L�5�.v�Y���Y#ʔl��w��3�@ēq��2�)9-�������.ԈXKg ��=A���(
m%�����k렉�����O̩��E�"Q6��i�{m��n6r�����o%���m p5'�uLau��Q~�x�:�R,pͮ��I/�v�Ҵ0�-�%�-�fB�����iL�!$/�b>�l��|0�����d� n)%�G����!�$
���I��4i�_{��T�M	�׊sa`p��dчF ��v�
����D�[Crն��uNi�����Ľ9Cs*�#��-1:��N^�|z�������D-����Z��u��PG	�VXV/_s�����F�Y�xf�+F"�kȅ�����ѽ�8�/n)y8�mC,^�f��'|��	�*L}	,5_�� ��l�)�{�h
4OE0��׽\��=XK�_�ar�Ț�R5��c�������6u���f��5Cɚ���sfW�B�oq��;V��G�-+*�	$A�bb�Ӕ��T7��ME�_�t�}k�x�"8�D�MAݨ��#��$��
R����������G�}��!LE�Q�!���F`�<��c�Jw��Y�ʧM�E"4V���_�F��4�k�­("��IǼ�R���C�E\�-4��64�L�AUn���¦�d��"3`�r;�7�� �@s��kG���G��k�Dڰ/��jZ��d:�5�`�ώ.�t��}'�V�I���I3�n#OhB��8lJ>g&���ʤ��ź6�*~��x���мn��dJB��a0��H��5H���M$ﰷZn��i~*>��b?c����X�ǫ�n(���?����|�37���}�����r&��e;���G���ʫ��E�0�mP�.��m�A�F(������UJ��.M�gu\\�MaK��D�t���#/W\�^�bPo��/(�I�	��P;��ʦW�`���+�0r�tԸr�&�xvݮ��$xn�w�aYb� ���ՙ�99""�-(��r J��|�ЋX�n�O����dBj�m��_	LJ^��	l8,���<O�����@.LC�߃#����>�	cT<3j{����b��5�G(�-����f��7��9�9`��_1���Y��6[�_���< � p5�
6ȇV��#ٚ��yQ���9?��K3�sոV��Zs������A�̊$ �e�Z��9�J[;�S^� �u=��+u9~��-��2�*5�`��&�6Wػ#wF�9KL�6*�+�j��<e��C����mR&L+C�j�Y�2"��g���0(��e2�������UD�5e���=P�E��'�=i���ƪ�5��[h!a(�=e�"�|^ħf�V���SKqx��O�[��]�)�R���`�o�l�$�K9���A�m7&!�+<&"�0
ˈRr��P�4\��2��L<I��U,��\&�M3Ѯ����=� Ȭ|d"y2�8c-��5`r�f߼E0���b�&�k,>�n�CI%�X0"�"Q�����S9��>��~����_є�)��9WGU ���Z@R
�Qn������6�����{�:9�}izXr��P*k����6�L=���h�L��JP�/��1����m��b��q�� V���[�;a�.x�Q�R��7N�MnN�n��yh*��~�{&��C��
�6	k�W5?�g�`���T��w�h��.C��	ż��.ݢ�I�].�bq�w�t��^��_Q�8�)	�j�$�"�]�n��?H��ƴ�9}��f��X>QL1���I�>oh���h�rWzn0�1k.�:x�}D��7\!P�A���c�P��oe\�:f����ԮU���i�7puovZ�ϻ, Yk4�*n����o���o�R��j�N� ���)�a=�QՊGR��L&����u$^�	R_d�D������Zr�f�6�H��J|�Êё�x�@�/��9���	�rWֿd68���y~j9�~j��&/oo�q��Ӄ�hqv�c��20-*���ƈT��c@w|�Z�QzS�5įr�p�cw%�qѣ\����d{��ԅ��|�V>=��J7�i�ޭ T���!���V���}���a�z9�%��*A�RX��e��|'�Yy�bUs����MY���2���!BƼ��,A�uqtk1?~���+����v.����j��ԥh��U꺞�5mc��:Pf*�Q2'd��b9��(B��ʅ�R�W�s��	/�����Q�m����Y�h�za��ꢩ��X2��V=:oӕHv�_Д0gi���!#�H���p_�x���g�s\�Ǵ��9�L_�*�y��x�]Kt>����N,1*���G� #��X
�g
Lv�a�]�q��I�����1�S����AW*���h�Jnz��r�'�:M��&��>�(�j�[�W�l�^���vAp5���K�ڐ��X9$��3�Al%K��J{ȯ� G����8i:��?�@�����>'A�'�/s����.�#�u��ϝ@����;�;��JUBi[�O����bkD�/����CL�mc��<�<W~�RC�������+��pm�Z#S1�q=/<b"|���s]�&LS�U=�-�)�6B�Q`M�N�����ZQ��c�~$��)ˋ��l4)���Vi�0�kW��&��B<A��Ŗvri�^p���}u�A�N��X�%u煬����NT;=�\���e������^����Y�cJ�W�v믇rcC����F�r�|�exl������m�c�Q;��Qܪgfs�A)�{0�Z�̗;�XV�G����+�D�f��r����=�t��݌�����z[���]3S���LE�qɵQ=)q2��è�+�hd�6�w0&Qkf}>�3��Z+�!�=�?j{z�TdׇH�c��I���m_�9�9Zd	��0�t[-Uu�XfǞ�%���0����X���c��H;$�`�ߩ�L1m�H}:�[����@��
� �{�pwm�I�G�MD�ζB�ޘ��񻕊�^W����K�B˱�i���vs�|u���"�:\������4�W������&!�X�˥wm�D�j�{�L������_QpY�Q�"�x�'���d�4ϓq!J�P���B�fG��"W�,`>h��{�&�|O��(�^��f��`��L���L>H��:z����1�P�ޣ�FR;�7�;���t�a_RN��r��4B���o9	�~�RT�!�zK����J�j&��W7�v��^�q|?�s��gO��2Lڷ�	$FXH�����������^�;��&���<�&�
󦡲��Ǘ����nm��U_����#q%��ͨ����vyt2���
�Z��PRY�=���k��O:��5ĞK�k����״�XS����<-�k�haofK�R�@K�AʕcT�tA�2�2�h�?sە�\�9p����
Z������z�Z��6-�O�ݽ��6��hoz6�.����_�����_�'�7�P,��!�|�"�ĊP�>��I��5�C��`hsP��vܗ����p$Z�����)�����&
4��h���2Ln�%w�^���t)K�T��-V>��H�ت�@����#PѨ ���?b���5b'�c����oGv@b�������ڿ�<=;���_3�������ܞ�Џ�����1}i�ݝ�6-���@Q�TS�z���@z���j���(뜎u�������I� ���a�K��z`�zl�к_���quS�k���ǲx�E �W����Wh���1j i5�zV^�>8�4r�@�܆�3N+`�ɱ��(�Kv��ʮϜ�1��7��� 5�-���f; [��-=1N�I ��e/d9%��g�\�(���0�{���/�1��* ������
	�����7��X�&��R��;8(�RyBb8L�������A�]
�n����wL����i����$�ˉ09<��Et�R&%���B�����k���gaAR�s:_m�1fr1��˕��U"7KGL�*��_%����aѡ��P�+O[&}t!� yWT2,��o��(1^e�Sl#ә�ˋ�R�P�Df�P�#��~�6��o�6�6��v���&��,���w��du�[oe1���&���ڟ# �"I�7vh��/��yge�����n�*`h�D �/�j۬D9m�uWmZ'�,�E��ZDPk�� RLh��U�E6p�EX�Cw�-9�p��Y��݂��"Fqb���)��,���m��K'���%�] ��èFq��$c����{/����q�A���-�f�����HG�!�Z����'&�|��$ͭ�	����R�f�+��� �z1"�F�3i�w�Zj�r.�&�#!Qgm�y�@��=�oŴQ�;ߖIN_��j�,�!،i�{����V����ߕ�wOSD��9�ה<�ZD��Ĝ�֙�� ����i7�7!��[u�����`�
%U��m���'�J�>���Ij��q-i�؉�t���U{ӡ�uQ������͓��-�K^\jC����6m��TMDL�%�
���z9Cs��3�h�u[Z}��h��A�"��©*���du݇+C],��Q�s(׺	6?t�F}�m�8w���]!���B|��t l��u�C�	yf6�ٴ� ���e�2﩮�%<�Yy���*H����4���̺M�Z:��?>Z��m-T�����$,9��L!q��7� @Û�P�����iDq���B�̬���;6��y�#�ƈ@�i,�O��!48	�īP���$��PH{��; Wj�u_8ODg�!�د�Y����H�уR��� �h�:���%)�	����ƞ3�=�Tk�R�g�g�7��O�0��ñ�Q��"8�E3K&��5}?�[�J�F�-�u��TJD�����5������Wc�]��	6Jm���&�"
���=T:^�5)�W��w����%��G��a_c�7���k����^6>5�{���r���<��竁�EkX��Qe����}��Q(�S�T�Z67���lJ�ΑKh Ц���3+/�L��B��|��ߡoԇ�ڣ���I~j𒷞�$Uo�p�#:���z/����̼�����G��$^�����oy�A�ߐ!����c["Ӻm!�U[�?�X��A-��@BH���EG
��k�cL(�� �;p��4(P��k�v�;m>4������D�|a�#vȈ�Cl���y�/n֏�7� " �8��v�_����'8��lz���y&��j�<�ϸ����b��N���f�z;�" cA�d�JZ'��k�A��f��_��+�^��w�Tx2޵~"��wp
�4�Ń����z�hS�
���Y� ��3����;ZF��j2t\[!~��mZV
0yJ��%5Q�[�4s�%��=�'�>HnW(K�����=v��@;���f6VW�M����,.	�)�-3��~�>�j��KՕ�,������%�Ð���%�0yJږ��Ac9)}�A�[�.��Q.���7��7d�Kw�=̭H��Y�ᒁ�S it/�B��T7zL��=|��}cس"פ�r�J`!��+�%MxF?�ZZߜT �W&{c,\?v��r|J�P{��{���kO\��N	�>��>%M�Q��#�wb��هG�8`��I�r����!"�b��}s�P��)���S���q����y�]ն*��V�����;�NdP�#7E7{_Jh4Kw؟�jF�C}�2������Sh�Z�+�sjV��3�� 	��w��-�8Η8y�l���[�/jq+*t d���۾}�?��v@��o2��9�C�W3�?���꯺(�g7�Qy�!�}r�$��D�F�'M���;�����Kᗬ�'W�S�(y�2�D�V����.�	�/0o3���uS�ut����M%�#J��X`��)�B�^��˺������]���}��͂pm�D��3�� �.T�5zeq]\�"�bI6ҏD�:�$՟��z�{Oq�e��}S������k;j���Y>L8o�7����T����r���n �yN�?��Z`�]>�Jq��/���=�X'槆�^��h,SޚE7z��8c��kD0��4���y�%ka'��� �.u�V�g?�����5���;��jꌖ%�qG�__��������Ѣ�R�JGZ�����8{^1E�=v��pI�e��id��Gd�h!��� eo$�a}M��UmNmCg�@2�M�Fr��۸�3��m<:Lm"��r��@�L18��|<�x��^|Y%+�`�GD��_��Ce��U�9�<�؂�����}3Fw<WAD�T��u�m��%䔛p�B�DL�w
{�~?�;'E��>�"�ħ�s��n�"�Q�;��P��zE>ب�Q�5a��*�j{��U7���|�~�Aݤ#m�8?��J[������d���]o�1�~�F۱�Ƒ���'��z����3�d����)�2�=HS��O�[H�	|��+�|�|��~j�Vx���T�p��b�""�ě����|���B���Ф�?��Q��TU�z	��N��E��u�-)�րQJ�������ܹ.9đ�+����oM'?l����N�D|du0T���w@�{;� ��$=�*O��Ax�&s(}�����l4�+\`�ҋ������vgAÿ��3��s:�W�{����;���
��LV��<:�H4���{����CV�E�U��Hhw�Ч⽵&�����) )�ۍY��)
���G㐲i��1�@��r���k��}���^���x�P��˒��+[���Q��X���FX�<
 ������W��8;|���T�k�\2�"n��7�gYr�5;6�4�q�����ę ЖQ��ɋ��|Gh˄*�8;�����0C3ѳ{����ujߎ��>�1Ǵ;P蹬����8��Hp�S�D�>|�e(o��� "����&{k�zk�7sM2�?՟�\uulx��i��ܪD�q�W��\�c7��'f���_�-�q��q���Uv ��~���՟����iG82KA�6�b�<�V�AUoN�l9��19n��A��%Z(�__��M?׭I���U~��B��h2�T�.{�h��	v~��b�	�
H�����?��oK���l�g�0����V8s��i�
@2��v�ߺ@kM���y�}_��۟��vM1�S�bm��6���BmмU�d�����������S���L5��0�E.ճ�����xYV��3��m�)����y��!�tf0��}H����WR+�+�C�]�:�b@��~A���"��"H�0Xt_��4�V�k�΅��$=�����*c�4m�[A��f�J)��7O�v�8>`��rrW{C����a4�}H683�hnz?���d�����į6[Х����C��Ń���WU�8��ՅȑK�Yv�Z�KǡǺ9�,��|��S����Uc�3J����R��+9�5ˀ3��7\�Xwήm�oE��G�da~<���|Q�@��6.�UI�'�E޶&V�˼��$�vNe6jR��N4o5W�k���:�!L;o�οT9��	^�<c{�\7��;{N���  ˜�<��(Eم�Yw ��a�x��h�[>����*�� Bd���~�ʅnU@^��B{��v�T��%�����HS���F:�8f�!�_�(�������tW��I��56]�
"3:����;��0�3�]ϝ��F����x�N����6^-K�v4�?㶑Ӂӭ��܀Y>�&�.�K��d�����l��+��g;E�SS,d�8���ܫ7��jv��uUD..5c�D�į���E�\?hh���*^��qY� W�	�!��%�D�D	�6�#��dK(�z"%jBbU�85�KT1Gt��sVq�[�� YO�Y��jsZ�nOm|�.G���fa�yŕ��М�-&��YX�q�	׽�] \��Y�߸���|�,}3��@��rFp��q���1���fO�3�-��XLJR�`3']����|� �����������8�|�Y|!-�����%6qC2RȌ�E��t?<UGKi����Z@�9��/|�L]���"Tdv!L����	l6�����b8W�����	^�^���To���!%���"���/h�ң��7��z�0=�2b��]�e��ث�d���1�l`:1�^��s����AI��p��ރO߄��y$��U����Ъ;u�C� %��"`����)U���ߺ�����#�D��`y��RF��v_�#��<B����֖㝦K69g��cV�G� �.v:G+��2)t�=��ۈ;L7Kc��;���4�l��P!u�:)�޶
��;m���<U�t�"@Iׄ���oޡ��(��Ze3 ����k�y���%��� �<V�:��OA:��p�s�gщ��e���S!R�BR�%����K 9'oL��EV���}i{c�1�1= �Y�Z��=�G���tqO�i���Ӻm�H�Ff�D��O1�&����cو:��a	0V=_�������a5�O'3��KC�}/�C�:�Y��C�s�d"��c_�	څ��/F ���φ#ќ2�]cY�d��Y_eZ�!m�Y���|������&���|�3o��[�*�"��bԡܸ����������T܁��_�>affdy�m��,i�De/��p���{9V_0��=�W���Z���<���>�~m�-�O\�h%P#�S�v	x������{��?�]��1-��uM��l<�悕��؃A�s��+����������u*@�Z�3~CǶ*ݚ���l�AO�ߤ�&�r�y��(2|aq&ޡ��X/U�b�[ ����"زV��k<Dg|�AQHٛ�XQ�3=�%�yO
mG�{glC�.H���� ��]�@�7�g2 m�+;Rq+�<�����p�t=�dB�ɋQe%�}����Aj8̾3A�t���1m������ŇS=d6&ogx�k�Ά	�XF���c4��g������@���G�&�Q,�mH����qp���b�g���5�S�{
�#e�-��'%qF��<�'���
�+�b��4kƭ���dH�p�z�g8��W`�SJ������xw��T��nޛwK��1�7d�=f�����%z;��,b��K6nuA�z��9��G�{1׊@Nܠ�/�6��Ā�e�(�E9�&��U����CO��a��F�8�h��x��]F& '���!
�F��-��˓�j�Т�9��\z�D׈�0H�i�3-���
�*�ѫ�ǳ�r'+A��j�͊�����|��+HV�y���9ە���d�rM�p\.)�rr��c�E0ٳ��q�#�G���;e9��kKr��o���!��pR*�����?��y��kK�I���57�s�;�����A'6�j{׆\+�E&v�6\~`��j����cyM�F��9vݻ��M��`�Y�n��V �I��B� �2!k����W��^��'�}���8�r�lc��X��q@>��ݢ� Z8�y�e�g��2��p0��7�ēۄ�С��/�����v<ȯ��m�nKT�
0��4�5��w�Dk\�e���;���.wotE����TYf	A9tw�weae��k�퀚(�V遱��?a��tvu*�#��-��A�w��l[bk����K�a�	U�+��A���b\v��Y��J�n-��C������C[_�1c����,N)��cLK-<t�`�٠\9=@��\��@cJB#�r�@�ѡ_�i�i=Wc��;V��fe8�fB��n)iM�/�Dϗ���~�7��Ə�N>��=����'m(���L��� �F��=��O�x�2���`4r��%�^Z5���+����;��i͐���	��_h0���_�bǞA�����������{b�}:9*Ȩ���Dc�ר�FS��f��]��>�Y9a6��ŭqf�맲��
^zȪ��NAVD�򠲬��c��m���4\&��iu@�u��<�sU/�aK>o�µE��A�]K	(�����/��C5([ѡ�%]]w�E�̗V���ƕ_�ץdh_s!����J� `�8���_#�A�ڶ}�&�>��0����c�y�5���Bk�#�~�]2�.��0s��T�yͻ��8��O�>��U6�\�N̿�Du@�e@��چqj��p&' pӗIk�ͮ7����:��Y,J<Ɵ��b������n�Ė:�L7>�P�~@�ܩ;�!<����N��u%CR�˞���'/u���J���I��"�תU�v�+X�!/�'ķ��Ve�b#�6n�y�P��&j�Sd#�!��>�:;�rn���{�n�@ԉ���]���?���mñjrF��X&6�����~,�4׈�J_B��cn���BM�U=P����R~{x٪-���<�z�Ofgd7��� o9Ct�B�H�aD]�#!� .8�U�v
z���*��oG��%v���M�+%�Cq� �[�iW ��8��չI�X��� �q�G��������a��<H�͆;��t��uWѣ�V$���+�zxEq��F���l��Y�� ��=3O:H���$���*N���9�ם�|S5���i�Z`����^�L��^H�����ݰ�����e"��hS�R�u(r/�U M ���0�+ ���+Z>�?K��y����ۮ甚�Q>P/���NH��CK����e!|�$L��l�|�Xj������ְѱK��d�+A��
a ����ݔ]�)- ��֧dW�����r,����^JK�>k�/o/�x��li~M�4����U��������@F �i������V�h��f�T`�ݤ5�Yc�)%��U/�oΗ���V����[�$+/�1�	�6>l�t�Sg��;|�",Z|`Iz����d���S�^<?�㻽���t_���n-��,7�Q%��� j��{	�!ly �4��'"8�Eh|�&�jƓb_lASu�CZYak�r3X�hىFO�P|�Iyk�k[x��cS�����TP����Q�L�
�"yv�f���\���V��`IP-���Nx���Kw��8�A��ɣl_�e��N�V���&�E@�:��l����J�� @Jh�#{s^�?D�՝��?�(u���E� WQR�������
�"��H�����R��<Ƞ^7pY�aA^�-�j��K��-���U��ҡV��*�a'yf &�#bp!_r��B:@�}�_�j����6�ܮI�~дDՏSs�XfK�	�
��xPQ�>�)��w<�y\60³��dv�+i!S�Oea�Ȃ���1JX��ں��(��x�'�E&��OratY�s�m�p�^�T�S��|y�nB�3���+�k�y��g��Z��`�/!��u��~=V2Z���}7�ʙa41y+*���?b����H��X�(}ъ-��@	��Q	�lLN��9�j����zu%-��tSb�6Ƶ.����]O�-i@-����@޵)��<��uڋ���0W:�l3r���ȹ�x��[W�O
E����_�hx:;ǟN58&�
ٯBHXہ��TŨ�r����{`�w߷˖6�6��â��/�x�(;"�n�nm��^��=�cS����6��G����q}"T3NC]h*��DHkn�	5�E����#�(�x�`�f7��K#X)z5o t��e��95��K�8Ͷب���5����c.S*c/��dH�pq�ٴ+#IB��c�k���6�l���z}pz7�vW��)L�Y�oНo���#HO%�t���pO�ORD
�����awM=�g��t�vk�ʈ�`�|kO������1ޞ�?���B�����`V;7�潖��϶��"Q#ܼ_%���u�K ���cn0$�7zM��9�aq���V���ԇ�&o3���]%�Ŭ��ʖ��Z����s���t@g����T� �����M�L�iP�Ix!�u�2[�x6N��a!����i��cdUV���e��;�sߘ�"g��fh����ͫ�b��˩���`�"���<��m���ş��P�g5�QИA�P*Zc�Gj/���6�b�m��K���=!&��]Й��x�(�1'�T;�98�[;�|2�E�������IsW$�8��!]�:��
Gߍ|[$A�@��V$ޭ����� s9��!?v5�@����Y�� P���B�hCQ\�*��F**��f0n�up#(D��H��,��֋���
o��q>�q,+m���pK')�(Ki�td��u����FKs[����&h6VJ�t�f�OG,�|��K9��d�E�D�N��jDv�/Ur�b��d�MX�+o�3�[�4PJ��K�w-�w�	]ͽ�����ju��G�^�94���߁���8p��tZ�.�*ĳǌ�0������E�Кָ��w��G�ח����.Tb��6cX:�u�|�A㈥��bU�\\������m�	(gs�0��VoE�����P�r��2qY~�,$ �"�բ
�k�E������1�Yha}3[��?B~K�w�k��6���(�x��.�ᇁЯːsƅIv�]W�
�sT�g����� M]�\8ʊg,�V:�P��n�����z@J��Z�+^̈>�gx�51݆sZ?�r�8j�%+5����"[�#3�ŖrI�Е�.^�"4I���1�"/hls��8���@d4;B%�8[��/�{����!6^��~;a�6��C)��\�..r�}?.�P�N;�h�������@?UQxU��ѻ>b!*>�P���L�|B����iɶ��M+}�0�~���s�F�YO�y�_�0"���gVHM\�#����Z�M�)��G+�r'8s|�8����~k�X�5�A��vy1
k��~����jG���u�ӉD�^x��b0~�<��̛��!��'$$�<u�3�\�].g�u����鞙
�28�M���^�?�|�Z!�y�ސ�dHoH��ⴅ��7~���I�F�Ĝ�D�����wB�p�_TU��i%g�[
�ݼ�:�o�^�?\��5/\���h���*��
@|>�w.W���i��3�F�:��<WB泑1��9훀aފ}����G�v�Rz�w�Vc�^�]�ؿa6u6��`�8#a8�'m~Et�RW��r߿#�&�z'̐�ϸ���_<�Z�w�'P�������8R��])���L��U�O��E�n�iHu��0$�pՇy^r���8j�^)���jqq����@u ˑZO�$���h�pG��S߁�\�J����6������.I/ 6����.���HI�¬S�~f������L	?+�:~TV�?�Sc�GHo�U�V��m��aH���6�j�)%o����� ���s����_��b�u݊�Mp~M�2@}p��7��z7���?5����w���1Wf��a����c�G|��FX��vB��' ;lP�o.PQ#������q�M�܍���H��£�bc��}�.J��AZ��d!����c�����H��t�P��	����Y�V[N$Fl�A�W��뤐�h�F�W����>9�G�/��1"]E?���N��3�D(֎����|��:�.�[�rsI����|��E��1�Y�7�%�w�_�"%����T.E$��,|�5����Lp)���O�J����n�g�z��C��I�6Z�}i��
Sl��������4�~J�JĮ�� �sCR}�&4c�Vջ�*�^%<�7�!r�Gu����(x1��vzL�hj�Wk=h���0������!1��ܣ�uV�0��Hޣ�^"��a�g$7�� um0���+t'	6��W�f�ǦݯĤǖx2O�w���)�����D��}���Uq�i�g�g}`:��Z�)�Ԡ)0��:�cҸ��(�T�so��z\0�D
�K�[��E)��y�%�.��r�NNn�u,p&��SN����!�q�'�Ҳ�K�i��0Ɇ����l��VJW�A�z2�/����~�+Zy���_4O�^0_�Ǽ-���X�ۯ���I��
n��݆�gV�ꗗ�3���^�pV~	��\c��&u y�r�&B+�=�o�%
����-��}=l[��d�H����یms�����J]6�J�ۥ�P��5�g�� y ��`��A%]�wJy�@k�&�1L����n9���
���7����-�[濫u�7�r�@�h���mf����7Jz&�&K��	e�X�/�V+���Wu�Ʀ���ђ��nn�����Y���Wǣ��d#h��Rc�F&�}�n�v�f_��%���N��uюD�8�%�WI�00�p�F5���޵*|@��mЏ;1gr�M���<�}@��Ocف �����V�,���_q�4.����;e�`zo���H2�Hʕ�7.���$��/;;l�9���<�Yv"h��c���8���2�"����F$��è���OG����6Z%)�DO<?��)1@C��&�M���ph����&�zd��%pv�J�;�*D<�W���ǹ�dQy��a§*�V7<v��e����??�Ŗ���d�_����6̓�t[��8�ߙ�^���%�7��&�~�=��w\�wUT7NG���bWk*�e�'��ǲ��m
��7K@2�$f�TBVA���LF�wt����x�$3�(��u�Ҏ��Ġrh'�~��C��3� M�F��'	�]B�!	�����54���u���'���o�I�T�:D�,�؜��!�H54�s쟥p�t�NP<�3K�Q0��%3c��$1,c�i���nt�L��yM}^�:��'�ܬ��X��A"8��^K	��λ��4\Z��w~8���:eDA����������'I�_�@�U�U)vUx��8K<�<r�[���l�t"�/ؚ>�'��_u��K�0A����ȓ�Dd�[���{��$jh�Z۽kS��_,��ꆏ�8�A�ܫ��7���<f
�u�^,�xiUM&��x�1be��B1�F�׉7*�:*�@W��6d��/Y6Ͷ��\�Ǒ��ߵ�U�"��Ig��m>�Ɵ�M��,u�(w8��xO��,wl�l�lzn�k�����S��enW�CZ�ɰ:�����g	 �q�4z�PѝFhO؉�A���R�+p�F��al��
S �S��Jk�>�F�	�|����s,����������;�L�1LԈqB(�����ßu��S���c���$��R��}*�"	ֻm��P@;o��J>?s5��O�
Q*�մ�B.,�X�m?�,:��9�ɖ��?W��R��]��8�:��Z�Ѱ�t���wmХR9�CU�s�4y� K�_9'5��n٢� 9�C'a&=ⳣ�8e����Z!yŝ:d�V~�s(Sjj��Y���	0	����t��s����nK(���$��Z�a���Ļ"�ДAO�+��҃ED�����qW��)����L�A1���+��P��ND�������:9'k��<��4,J��:s��醴�P�k�J��.�k�-��+Ff���E�aA�HfR�/�
���VJ���&%�o���˽�@�m[Fd�GYο�t~�����ܺy�b���l�u"Ȑ:Z�~"�y2��?ME.з|� wg�G�}sF_�`� G���?�Z���v�r���������_Z�Tq�����!]nsG�~}�$�A�-�g�|�ܔZ�ƚ���?4nA&U��ˊ�m�⨂���uk��k�������I�&'�a�L�:h�+��*� ���ի��z���xy�w�*��}�7]����DdP/���jOX�`�����V�i���"_`�N^@�=Qv��@���1�">:�}�Wv�;A��&�n#h.�E�L��3i��}}��	}��D��զ�U#i�F��_�)w��;�mBT0�H6� ���+S�i��+���
B�����d�T$�M�u�Z@���+��V�W�*���-���i�s�?G�D���F�hp�s���Œ!��Kk�l��4�N˺L�ב��Ȫ?�������$�5 ��FN��J����e�C��$��W����'_q�Fx�D���&�ӾX�H��Z�pt<��滛�a15�:���J/w~�_�n��ĥ�����& Y6R�Q!��Мƕ���ǅ�tcgT+��beP�h=E�~J,U�2M8*�p���_{@�[���jI�����T<a�$5|eN��U8gY�9'�؝(��}v 2%(�P�G�a���+�V�7�΢�ڋ-�����L���PV\	� įu�LJ����Iۆ��ُ�\9�������`��A���nd����o$�ḛocQ-Z(n_��i}�s��~}	~��S�LI"f�t)�-��޹������.���������A�ֵƎ���d��[����o$z����1P?�Y�oҦ��Q���.��vIP�j7��5L8HVC���J����q�W[c�!Xh+���ؤE���Q>����=�\h	��u�D��r?����Wܕ_ڇ� O�'��<�zīg(;�7������R!�\�D=Dt'u���q+e`��IH�7�I�}�:z����/����YP&���򎢁��6I����w��Q"F��6�$�������f��YEK'�U���ׂ�k/�8���J=lb���������F� �&xo�Ϧ���_�\�&�F$���l.W�(z|�?Tye���'��J@��ʃt�Z��Q��b�h|�)�QvYA��v��؏5S�s����r�Ec��1Ćq�R��j�J���|f�d��>�#aN�}�V�@ ���!�_�o�Q݃��FAO�&Z�����ɂ�+ɟ�ї����(.gOWP�G�d��ӱ�(o.�Ό�+��	R��kΎ�X�k4��9}���E%.3m�����#_\���yP�椇t�~"hL������Yga!���1��� 9���q6��m���,縡;�*b)A(�P'[:>�����Tz���cM '`K�
�b��4C��}��#�Պ앾x�eZ��;r��D	��l]�_Qq__����U$<��!�<zr"+���?�����>��3��"3�`o���ؑ��}���J��j �z ^�fgZ��!M"�Y����������巭=���b���t�4�//����-0cx�UQ��2����P�(P_��I㱫A�(7��Av��z�zSºIs����Ō(�7h|I���fnl����9��|�':NC�t�
v*�1�~�`�Y��XxA���x�y�2C�z^U�'� s�lD�^"{���/�Q{�����#�Ȕ-��0��S�l���i�_�kr9XK�*R�l_���nf���ӹ�X�`�Mn����@ȴ0�h�虥XF�zj�t�\%?�~wR�E��)�� .��7vB�a���@�R��1w\:���[լ���E}	I�M��-�"·�]I��4.��T^@S�hE�26�L*)hh�;NEV�>�/�MG�b�A���Ṛ|�-�3�ёGt��4�9T�#`(�i��H�xM���Aļ�`��J�^����H�ZlqQ�ɿė~[6`{�Ҧ��Y��5"W7���qP�Sy�8���΂�����8c�y0=U����[�Q�ںF�v��Ԟ��m�R�祶$�Go+���_9&a]���2�ov@�zf��=�0Z�a�rN�R��U��/Z�������\Q{!lj��,\ނ�}Ӂ~��r3N�J����y������d�'��v�Z5}���A[��=北�$ �r\y)6/�����gȁج�8_63z��(�C4�K�Cʪ�s������#��Ԣ�0䊟@�bLх�`>�4ߴs'�ƨ��� =�ri�V�.x���Y�#+o���c���VI�;o�q%�( ��8�.hɚ�>�P'A|*��yjG#V�4��|ߊ�!�6��p�u�55���aC�T�at�
���M9�ꌕ�}\hL�>��.�o�8�Q �n��wgb&H�(�����Uy%�v@Rh�va�����Z���Bز+�Lk>�3��&���"K�m˻E=5a�rŰ8̘�����!Ux�E�i���:+�i�Uy
�1���D��^#R�p�n���ۊHz��� ��b�Eo�@NW�0<�/�%�����L`���f����g�N��J$��
<�-
���P!~[����VԽ��gRp�O������X�Z�A���R�4�	�\4$)d�����<���ϗ|-�|$2�_k�	{��-&I4�d�Vs	Ȍ�2�s��t��ޥ8a������pD�[|=���1?����g�a��3��}5����=�}̭����\�UrdS�8������9�OoT���]Mq�77�)�g��T��@6��D_�EB��!r����M�%�p����7�u�&���QNazԄL�kD�:A#�g�v]}�k��Z�f3�F:��2a��+�M�>�npBe�-2���3��a"s�7������/5,^2z��tdkǌ��Dt���%�@�%���w��TEoe;�.C��	�@*�#������yY�"p�d���
�!�{C�Woi�ؒW�����P�����Ts0�D�m3��e�<E�']��[`���ꀑe�5�H�=�82R��G��j����`�P-hNݑ��(���C�~E��?Z#����7HE���m�+�n�?b	J/Mc�<&C�z���O��Պu��9+�*0�w�Js@���&^�^��մ�$����9+�����[�@6�����B-3uG,��o���¨�=� �K�؇)o^���x9���s���;)������*ܝ]CF�v|5�`-�r�q:duE[d+��	�@�o{&_	)�	�{_�����f��H ���h�����(1))���S=C��Ƣ;�q�i.��	��i�UJ�p����EI� b�ث=\��u�-������E��۩��C_z�H�5P}B�˓DN��>ۯ3:����r;Ri�����FF�W7%�s�r+�M2"��Y5B��w��W�.y����l� V�1�'5v5��A/�֢JE�$�~o���	
7dȰ��A�+�4��?�)�o�aةM��?Y!	w�g$�9��|�N|��P5�Z���̫���S�&XZā�L�T1]�^[��Z%�w0Z��X��~��X�`�L0q2
��)X�}�j����b5UzC�d	_(�F�(W
j�q�"����'	P�K��.���ȉm_ -Cs�+(uc�\p�"���@q�F�q�R���Y���Ρť�AU�,�CEE�얖�!|-�U�ߖ=��ѭJ ���D����3Ŀ������)�������-Υ��+�;&�$j�РC�!w� �S;��}��Z���"����Ҝ���M�i��Qu�B�5��|'��n]�F�Iű���Է����&)p�e��E�2 �R߃��[�g��`+lԾ�2�������}�����t�8���|�yS�]"x>qH�>��D�����ďG<&xH�"���}EoA���*�(cko͂�ֿ@E�<(./X�.����^	���� ��76mCД�cޙ����o�W���|v},��r��pO���Xa-��%-� ��u�,�筷�x߽��D)�(ZI]U�/Ez��
sC��.�\��$��lu���*��3������%�4�xv������Iɏ;x�8���>��~L_� ��@=am蹾�O���	�k.H���圖m+�)T�yJ��f������nm��l�?��Q����wA��o�N�2�])�(���o�9>E�I�gU+�g�vw��ʼ��t��I��=�!/��k}=�6�(�ڄS1���;�jG�5||
9�[�	���]�t��-.�ʜ��Z>�&RE�i�zr����6L�O�5�ؠr���$S9^��gz��5!��D�˂�&�y|���$YT7���X��+�V���Cdp�M/�þ��qJ�}ǩy���|\�aJ�Rieg(0\z��w��(0����1��%��ӆ�3�����Uܯ����0GiZ9c���J����/_&�Q�[L'-:Uq�92YenXtPBHt�\ת�LqA�o��p�f�O�q���M��R_y�|7�a,j-�h<u�ղ#KvD!����ey��Z�/�ò�����z��(���V�>��i���м�:���+ꡭoAB��P~AR������AlvΡ|}�R�g�K(����p!xǧw����;�L�K���>� �T?�^rnʞ���mQ;�G�'y��Ϗg �&m�WL�j>F�.�r���h� ����`���[���W��/)���7EdZ���kR�?����_�t9O����\qbV����\���0�U�qm�~,4�X�u�o�d�sg���ya��7�P�`�mI8�П;l�8�OJ����V���^��"OL7���?�`������G��
Z|D��g#��ϳ�G����u��ϧ�x�~*c|Q��se�~խ�lFy��#�^��V�b����af	+|Ծb=��y!��cpN��H-�%�Y���A��}�� (�r�"��@VS���ŷ�nGr?[6U4��S�ϸU��j]H �j������֊ѿ����6ٞ�P�\K۸C��I�����5
����uL��9w�x�K�n�n����C�J��vŔ��+V�f�t9�L�\��{�3�8[2�c��zg��x)q2�®�����0;��PB�����
�E B0�q��O��L#�:/�]�PH<F���7Lv�Q(�
Z�Ђ��8��WO���:'=aS<�B�Їz��*
C���u���*t�ϖ[��zO��䤱�.�:���H�6O90K�[,����jZ;((�:�Lr�X���-S5���+h���`���W���ֶ>A�`$��Y��8�#���s?��~��/�pQ�˔7����Js�ə
s�&?���gmK&�i,0�<-[��b��#���	>�[�D"D�f(7=;�fPH�C*�ee�ދc�M���P�=�=��@C"u���o���
���u���	�j����5� 5���u%�=h�֩�KrԸc�L����皤�G�px^u�7� q��;i�#�h��&M5�ӵ�W.Ө�y�3������N(+�)�6+�5(����w����\�U�@��5t���V��QḔC"��8�.�:������_�>ٳǽ.v	�XЍ��9ꘜ�p	��������+C��t �Xk�5�Ӂ5�v����sԩ^�Pذ,�P�OȻ�߈�� ���mU�mIa����ʢ&��|�簞l�vuP��Y��:3��KjbO�Sl������$jz�����_����8(�P%�,�����0�n��p�:kĹ��};����)[�j��-Bu�
sZ�z�(��ݑ�hI��su��4o�^��`D�����? �F��#u���BM}DX�:�fnr����#u��_17!���N7#�w�3�U7�ܾچxb�̷�0�f2����D�\x3��(0��e˶E�\�~(�y�=�B��BP�r{d�h�3=Z,^���i"�0��8={ ��Iq.��l#�P�"�������T��V6 @lEi���機�V�\λ]���ǣ���a�Ķ����[I�xWD�%��H�����6�����{������
:M6W�m���wk���5������٥}4�J_�z�v�d�ɻ�`��_�N+]���pQh��O>��p��md��[�j����E������r�/ʲ��i���ٓ�s�<��������ٿbZP��(��)�����BMz���n���vh�m����S��/����"' �^<����lo����)���Ԍ ���A��7�F{xs��!?�I���4?�����յ�" k�4`M������EƶFW[q��ᴔ�Wp��HY���+6w��ʅ�O]��t	oe�PL�u�7�oT�L�L��0��P�.L�v�-����-VUL�,/��d��m`�]+�i7�&MV`󡅳�n��_���?�!�υ/��?��J��B�&�w���y�R��"�Za��7�D
���Uw�k��N�� L
Us�y��M�v��\>�f:Ug�Ro�,�NG�ܞX�<<�2��i��Q���3Aꉂ(���Y�I9������N�/�F݅Wĸi���O���6SR;A�O��}��
%�~����������n6��x�3-Hqr��R��mIkoe$M�בh�X�r��/��[�y.����vY�D�ҹ�ε�ݣ%��m`�Z;y��L�N'?���0=�G�}m �g�\{SY ��H]�B���T:�Vb���:zduI%�06Vf����@������W�c+1��=[b=�P�q�X���
��}�V�I�n<5\����c�N}k�l��`�Ő�;H������o�q��H�������ⷣdﷳZ�{��=��#]�#�����OY��x���!�,!�/"�
��}���͝����缞�Ϣ;�m���[�!�E��p�mͅ�R���&�`�K�զ}�l��P�H)��1u&���.6ΪᣵbfPX- 
���y���nu��+}��&�������(O|�˄{u
��*=4<�>�Ѣ|n�W�Imf���ۦ���q`��nhClI�[���Oh�+^�v:�� �~G7Kv̀y�i�G�^��/a2p?	�a.'��ɏz˹Sqv��x��؀�HeF|�Ɂ��М�~�>V:�d�,4�K�\�KЭՑ��2i��k�F`�(��+:y� �2�45���U@������'�8�{'Y���tS�Y9�#�@��<��k�����L�XqAP6ZL���#�m���kh��
W-��WyZ����ݎ�3d/݌���>�Ws]bQ��2�K�������=e�hݐ�j|3}y��ksq �k�`��gmF�G����F�Ƥ#j���+�W��f�E����B���ig��^#��B�	?~��u�,�8x�e]�]ۼ�<
��������$&��#��b�S���iF������25�s�bj�
��y�9])��ɫ�!����9�����/���A�!�<��[����y:4 "4��m_A+	؅��i�*�#� H�����F�1�M��� %�����hh�_̜Oc[�^6|�����\��&�>�K�j�j��V� �Zh�Y��[�R���r�k lG�it-�FO{�數S�������AT����Tp�_�:�a�߅j&��nZ^ѽ/�
���m�@bI�끇ڪ��Kw�
��'�r����J ��;Aw�����I+˃H��Y&%aO�WQ:VYwg]g03�7�7�e8���O��UYB�D03�Tsj�βC����[	��f߳���Z���H��HK���;D�!Љ��mYÄ�f����3D�U?D�[Su7�ڞ��Z����I
��LᒤVUr昋��Y�Æ�SƲ�=n�%y��i��=!�`�Z�[���̹?���e�qT� ��)q�@ʹַ.V���t,l�k.J�%�8��(o�_,c �mȎu\c֭��e�F1����0��ԳΘ6?\��ჼ!@)��9F�p�FQJ��7O�bf9ּ q+�pԽ}��烓	��k0�@�o 0��	�}�R����'��N��A��a&[�gP�����:�Z4k��R��9Q_��+����0�n��6��]G�у_�s�x��]���O��H��>�������98��V7�,�M�4��(l����H���`�̂Χ��!q���Vm �S��Q�`Q�Y3�<zh�����?/�ql������s7����9vp�n^�
m�V�V�����?T�&@}iᚙ�+p�=�Y{�:�����Ԝ�+Y��p�pc_�g��6�1�]�!D_k��oI1�sį�Գt���BMmy��p��9�Ny,o��l?H�B�¾�G��l�RY���L��2�P�d^��� lt
�����p�tS�W7$�L|@��\��sM!P\������C���d�(~M�E�U��h^�)��J�����:A�R��F����M�f�2H~�m�r���u[�_���n�ky�����ӶFP�wC���-�_%9�ɟ*A[�Q����ݯˋ@�^��	���Θ�U����I, �@Ϟ���:���y>��g<�������?5�Ҷ�@cW-~qEN&�緥�CR�mz���)%TL�\>T�5���7"/&@�k^���}b~�;b;*�H0*�5�ʑ����ŵ�z�m ���6�̿�D�v[j{�e���pi7�U�$"��&[�W�,��52���J0C^���q,</qD�Q�������8D��U�8PCJ�]B����������ײa;�Rh�!EZe�+������$7��]������R��P}�����L�vE����YrѪ���]i�������(�*����#���A�V�J]n�)HkjI��p��u_�GA�x>	I	Y_S��B��A������	�����ԃ- ��s�������B�;#68^:W���+�^G�	��!�1do�.�c��$cԃ���r�6�h��"z�����\��"A��-��.��mx��D�C@��?�\��=��F�s/
1�m���F��M�ù��ԓ�GN�A��'P1�w+�Q�}&�;B\��1W���_	�QS����L�ҡO��Gr�w#��������b׻��ֻ
�q�+���㒔Pج�x����\2��8��t��|<T!�	�a����9)��-����]$����
��\2bL�A߆6�uA(c��:�Ԉ=�G*2�,�����^��b�����\���c��h�i~��"��ħL�ic}n�ŉDJ�[��G�}dk.0�p��w�$��t�4�9h�<FE�3Ϋ'~�a��W7�QF�r/h?�a�F��֢fL�`��FdKŎ���'sG�s���q[$Y"���}n�в�o.C��՗�z��޴�fO�\�� ֋�{}��2��MA��2����ku�l�l7�u�	Q�o���s��S�*��f�Јqd_5���Q�1���x���ϲ��A�`��ݔ2B��~� +1U@4�u�I��(���4�^�U"�Z��MWL�#��_�ͨѰ*{��]�"}�#�dQ�J�Z� Q"�~_)kn$e�sQ�їG�3����# �@뱅ϳ�?wP�1g�z��o5� �ar��VѰ����T�Du�[.��!��WX���h��r:�m[�l�J���ͦ��I:.$��O%3���<��m0����6��N�����sj�Kȿ
�}Jg�ГLl�
X�d�o"ضum̸F�fy�E8�R"b�'�U� �E�x�ǻ�V�@��ÐTj�G5~��ˌ͋���0�����O�b�+���(�����n=��!��g9�<j �v��'��S)/�,�Զ����"w���V�������i���nq~"ފ�y�<o����+�ֺ8l�$��2f�h���t<s��,d(��ɷb�W���5(��he	��������u��noY�q)����	������0��y�$s1�d�cI�3�o�%���3�x��'*�@�����,{� ����!�f�z�E>
��g!&��[����H���Y�L�/h����):U&�J��(�"��6�;��S��xFƃ�#��2{F��������h���#]��ѕ�FxJ���O vwW�>���h,"gf? ��BQ6=]�_��`9���|Ay3l�	�2�}�KE�B|��W���C�8���ؿ��w�6>ɥd�c�I7V:fR���,���C������5���Q�!���m$G��^�Bk�2cj�ov��r�v�/s����Gp�x*M~Z��|���%��nU�!�/JiA�RE�m{n�.>��Oϙ��d~�&NQ�:0�p0�Rz���!����Aɫ@O����r0�?�>��<���Z+]���e�q�k�.+Uj��Y*}#��L����,���PB�4/�tc�+�Iw�1cH��ASZ���3�Jev���(:W&�,�Kp��f��\rʠ8�,J\C�#G�r#��$��J:V�:���-���\Y_V��T@���U�ۦM !�_�%����ahodIJ�ԥ\v!�>g-H-)�(��5�If���BI���A�:�eR�Yų����C$w��ē��o��hxGa���#���,�4~8HUإa3����E�>��;5d�*��}s��ɗK|iU�Z��P��P���2�S����!I[��ˎ���~�/#�sS�5�q+��		�����}Y�7$駭��qm����2s�������̍{�r ��1����,�<le�"Q	��v�@�5���CT�W/���W�6����L#a�������2U���t7�$\��H)ǭ��Q�\��[���� 
k�2����C�ȃ�^�#���^���c��<?���0���ad�N)"��pwlSl�D]ƄOF��]�Hu��炀����C��W
p�+��'l�J�-o/
��PV���:ko0�Bd��)'X�4�Q�ѕr�m�j�@��Zbu�Ů\�t1��!~h��/��F�!���˾�G��J�`�ɭ�ʊ�G��Hxń���G��+��H@�x]�/��+t��W�ON�4@n�M<�f�VS������"�/J���߫`i������D`9C'�k�#�}�DG�,T�����>�����]�u#y(����~טe�~H��6�E��JY}�Td}���u��|��V�������������+G�Uƭ��_=�cK�uΛ�Q��
�(H::�;�=�,�x��c�=r&E;V���
��)�>�Yc�[��XJ� ��0ӌ��M�z0G�cA��!ePp0\���y0)�P����kY��=��1�H[
�c���؈RulwMhp�`ꧥM�6	��A;�S�����za�TʬR��k���w(����.�W<{�'�&\�GH�C�������ǵ�#ѭ��6-!��$U����w�=/L�۪�f?��R`�}_l9���l)8�ÿ/=�QYA�������]��!��mPu��$e���hv�@*���f���
6:���5B�$T$늍�Oo1Fz���>��4w. �4�[Ԫ��yB|L%��g�J�-��V���Ƹu�t	����QL�&����u�̔����6��W.�@D�Ǫ��$�-AWd]Wh��������?���&���W��h��ָ"�Ư4��gK#���;Al��0�m8[~b�@��:C��}0���A�x�q�{H���^s� �u[E��.�����VJU��0X�z�˗�@p[��	���o�#�����eg�~�Ѽ�2բ�H��v9�ε/Bl����
�?��cc�0;�U�?�-��gg��g��\]p]�%��(B��y�dökq��;Y���)�O9�U�E��	qY�∬�bI%	~�����,��W`���zE����H΍�q�8�pk&k��.3�˿���[xF��&��Z8�YD�À��ˡ�����<Ų�P��p�A�J�|N�~o�qR�f�4) �
1z�)�����e�2�W�\W�e��3�"_	I\[��d�_��f���H�4>��
��%L�a�Ї{�ܘ�7d �� ��;�#��50��g��`��kޫr ��ʗ�L �f�awA���[۽Ih����_(�	�LrPF�l�|�+J�1�: ��`L�mC���'j?���0�2�����l%�����d�U>��j��~K�-]��P��Xkst6��u�=g�o�W`���o�cO�d�l���v��8����HYk�g�ٮ(_f|����#u��r;���7;��>���z����)�0��������"?��ux����J�3oz#6C���|��<9N�#�yT����9�>�x}������F�Fc��+ju���9���B��^���MqDsrC�%c]�<&j�ڥͪA�jo��XF��qI��%�8="�/��(e�p�.�^�G_�w3�v,3�@������羇�L��K���'	$&M���\H�3�H�Ҍ�%��*�nW�����m�B�]?�̹)H�j��&)��c3f���\�:J�=I�U�|��1"B�~5�TZ�a�`�u� ��򆛤B$g����e�[�6E���XQG
��ۼh�r5M��3B!��o8s�+� ����Ôn�ԫ��^�
.e��Τ�C���E�v�.Z�,�]9��(8 ���d0��(���J�i�ۋ!l�O�ćj��#�?$
V��-V�E)EMp��R�I3;ك�&ߪ3�-i�O�a%-�EBK.vˠ��v@���e6�Ma�=5���S����R+R ��lq�ᎆG4�d����&���&sЯx�w%�.��7��N3���1_E��{p�p�7��L$���_b�npՎ�r��n����W`ߴʙg��.

.n����d��]���9�H�[#}�&�F��\�	 �I�
\���Ћ�X��شsY`��J��Zo��!��Q��jSyf�0����e���$��t�QB�_�g�p�~ �����f��@�_�Ȳ������H~�ǆ.�6�<��?@=��Tz���ʤMZ�ŗ�+X\�g��?������
X^%����X?y�J������r ;l����9�a�eU��qd�|�`^k��P�A`m�/ce&�P��o<�#S�g�?�R"���u%m��2�oG��d��h�.��%���ӣ	p���)���v)�;Dg3۱>��� !]�P�UY���H�5C��sYΞg:���%�?�nv��!I�<̈́o
'	�Ɓ! _y^Cż�.�@��[o��j���}��x�9b=~Q��V|�_y�c�=�%�M ����a�$JlB鉘D��3y(ڐ4�ߘ)���4�>�&I��܉yz�����p��J,����c��2��Ee�hr��ׯ��n/t����,~�W�(\;�eWӓsG���d�cYÔ�(�]��b�|U.~����=��z�����W��f�Y�
��-��M�: M�����+S���O�����1�'~��s�G�65��t����\���9�\W �)D<~ƕ��� p��]��)��7
Y2�sʳ��רTŰ�y���˴�c�-�u���f�-�$�C,P�N�	��
)��݇�ś̋s�
R�G��5P$�h�%��-% f�D�?�-�e#�S4M��]�&
����D�*>��8���p2��5��4�>�������9FD�.�M�U��m
n��F|��v��h�|������
�}�g�5;=C~C��D�v�_Zm
�]R{������բ��d�2O�ʥ𚻀w���T���v��7X}�}�~�6��R2W\:��J]>:��ӧC��F�>�qu=W��۝KJ[9��힙z(C��I���>a»盏��l2���Ի��o2 B���ٟ�Y�|$e��9+SwU���$����x+��v��R��]\\����(����1�xni-�rE~U��y$���R����;�Iڞ�s������:���w@M
t�9�:`�'������g�|U �!�Po[��K�$Pؐ�������@sD���,n���tQ�&j��<�ops6<,�%���#�ct@y_u���U4idS�ׅ��<�T9/����}ຯ�<�T���>�����lde��@l)��1�,¤:�E�� ��5گ�����?B)��	�=����1��T�aAO�*�m\�����I�������.s�D�K^�};E�O`H��pr�*4x�ãmt�T�"��d���� vm��Y�/���b�D����J+����'X&j$�4�x#��g��7��[�\J T�y�k3����H��.�j@X�q�ٺ-��!Qe���CGx3�� �rpJO������ ��xɕS��R�fF4�D���=��B��&�JH�膍n�H��ͤ�����?W��q���[����S�p	e�\G�8���-�r;<��YW\�DM�C��� 0 ŔAjB�z��b�L���>Ki4�R�9�a����a�)��w!�K��j��)a�XenP�Р%ޚ"������"��C*�i��p�a��df�!�i�;�.)�WƦ����)b�	��'�i����o��\�
��y`*��꿎�@iSj�Wޘ��c�LxF�#�x�����%tm�����vp�������Ő^����a�6OU���xU�oL�m��?R�ėJ!���"��l,��33�~=�Ba��ad��^�F(}'"�2�A�E��_�c֟�ඵ���&�\_���K����r��>�)|<Z�ě3t~c(B�	t���[%����}��I������c��0��ʉY�(�c��_�?����#PU�� �և�eK�bb�CU�*��������H�����f�d{��M��~���͊K. xg��U�m9T�׋P�*PF�@�	�O�֬�!�>o�?6��֝g ��s���V~���&��_���q;�nS,��tӋ��/���ӯ���	�Q;6sj�"Ls\A��F���&�����������:VmLE,q��t���1!�&~�oRro���0���������K0�D&�tť����V�~�C�vxs�y�r37�u��3���)��7N*^�ah�t��σ2S��H�S��Q�����S
`נK��c�W�e�x~!����J*AજtݸpE����������,>�)�,�,�V~m�M$),��}����t�1f�"�������T��j���U~Y
G����A�-�m	�����S�f:R�F�-tJ�ź�5�����{��Uݚ�k�L���D����]�>İ�ʏi̭2�� �.%O#H��H��WJp�I��k��ୃ���5(�s��!�p�ΈAt���w�,�ŵ�r<�]1��-�k~e���D!n��v��7@���?O��P���^�[��LZy��'E�B+/È�	cQ���¬�f��.�q�czK!���mS�>G��V�������>E�5o���0u+��3�+����`����P��� ��+(ŝY��E��>}�M�\u�obJ��$i��)S-�7@A'��ɗ̹�h�e��y$���P���8��;�D@���R��)ZSb�9�-�J�Mu��1�՘8
� ���5��d[��¡��]VL7��d�g���в�|��$��ە�j�}��Qǋ0OS��ר��.= �"G 9Mq4�*�n"w����y��%�Xw�NMň�2���a��O�e�xr;ޯF,�F���%<|������VM.V�1Pș�����r�S��`O]��pu�����O/�#X�]�'>�Of���[���Ꝏ.��O6젣]�f⮌�aM�V9�d�!�.
GΘl��rM2Tє�ؗ5�&�'3Zm%�`{��S�ql�,6|"2�Y���o��h����}���(a��Pk�e2 �&��P�c\ιb�r2�^LA���1��1�g}HH�Q ��Q�vQ�Ze�a\qM5�gq@��ƈ�������J�'�K�qP�4�c��uUۚ��v�j�g:^��Z�͗�V�(�S�:��n�e�������d��Z?���]��e,��ʡH�_vQ2��[%�V��% �,��:���HStY����um�\� o��Ɣ2��eg��*c ,�e�e��}�,�2J�|9c���ṁ1��w�����Lr�7Z�,uZ;Y�6o��$7�ٟE}��b�8��Ii�DǋQ��ѕ	zTzawT�W@���*~�q!��M�u&����kf�\��0��aa���V�>&�:ޠn9w��=�	�
hJ%������Dɗq�7�읯�y˯�3j�������J�.�Od�~g�c��XL>����p�K�[W(�(�d�2�?R����P;������� �#ga���5���N����x[?`e�Ӆ�>ؤ�W$��tX3��{S�?xr������1��>-s��=\̀Eb���ػe��d�	]�1����壵2�д~�b����낒�R:�!���!$���nC��L�過|2��hG�|1�ْI�/v����bNkD�Ф��Q�б=���y�\�֎�w��%��X�ݲţʘ���g�WR��q}�Ko:��l����_�k���<��`�]5�`=�+��Rѓ���eݟ��^4�r�y�,�t�H���^
?a����(�p�5�o��=���^X/J���i.a��!]�E�M7;Xۏ�«�z�ßв7���;�`��
輫�G�J]�����iAR�2%��D���}uZ��� ���oG��&��V� �3�oe�����P
c�&��%�пO��5��H*>u�;fހĔT��"!�+C�?T���3�A����ʨ�����f{IsLJx���?R�}#�4m�(��X ��3�]�n�g����D��}
zw
�6�˪�a���O;1�K؂�x��ѥ�L�1*�Nb�Lψl�K4�3[@=�����[�'`�7a�0��h)X�"��e.>�AK�9�s�ă"^���;`�8D=F����_��ņ����Dm��0����cnZ0�=k�k}솖�ґ=]L�����¦�7E���v�Wv%h�U n�N���F�'�!�g���6�To�4 v't�YU*�hr!��rDQ�Cn�1|����$��Ĵ`���S�Y�%�R�o�����6��Ȯ�a�<�������Ja�U��?��΀L�	�zi|�A�[^єl��'�ې�uv��Mt�h#�SNȆ����1��DE�do)%b>�3��{a�EM��$
�Z50�Dn{r���<�?fD��u'�>��A��>9�J�s�d���?@g���q�M-%a%G4F�Y�\5]GH :�B�0�D�,�t�*͢��t�p���}�����K��P��s#k�Z�ɞZ,�媻Y�=�����
v��`G� p�,���M����?	�:v��K�<�&f6�§��L0�ڪy����x�-���pU�b�r��/�Nْ������	�Y��x�X�u���r<���յĝZ~�_�[��GT2]Dc+�{�"4�u3Dk%9��y7�`[��_�fF��_ 9F��4��	���=��J�/��
	�'���a9��l�+x�Pk5�vdapٓ_M��c��s���9H�b,pۢ�5�Di�|�4S�= &�%��?{��RA����5��,r�<���.�����:����?&���M=�7|qUe-�������$���������#E(B �-�X[�J5z
�:��1�V�uG%`��}kp��{u�S���^�&��\��z98��`�5D�Pڇ�D°�
���wD��
~OU���R9��
�Ԯ�ǰ��2H���Y�~�xРT$�ԝ����}nzT��64����0U�\�(�߹�eoM�o���f�t��&.�������+y������Ea|��&�u��*<� �{���G�9kI�Wm0��Ĝ}¹W5ԏƷ�6�dU[
��� �^ }s���A�_��g1�+�c��uYMG������N���M�#jj#خ��TC�,6���$pN`���G��ꅋ��>�Xe^�`uwp�/�R���4{�r�'�75mϞ�	��F0�X�Q�G�{�������8���?sR���W�5^��~e�h�j�� �,H�0�<�b&kmG܃\�1��}�g�b51��P]�r.��U�B:��k�Tʊ$��}^�[�2�3�T1�Z�/;��	d׳\�?d�F�9~4d�t��r��Sh����I:	�;�Y��:�.���XN�>P�#e��}��Rm��^��߫����%]NAotτJcx��<P6+Ɂ���7�,�����H@/��A+L��:��t��E��Pt�+*H��[G��
�5�,�/�)�����Q#�0�ӑ�
鯾���^TC٠\9}���Q`3�>����a�?��	��l���{_9ɷL*� �[�Ou�l�$iG�Ex��4��sX��7rU��G�	��}��Dߘ���]WD`��6�׮OT�_ۼ��~࠴�V��ч��Cءc����G�+*���{�j����L���	���$QT���j)�c�H,E��k�Ԅsі}E�o��ׁ��4�S@ۉZ��R���17��ԍ�\�p��}d����vκ!Y���N�-;ً��ûA���`^�o0$S�� n���M""��6߂^I�P���),[�z�GjfTw����'z�YA�Ye
�Y{E��}�q䭡v�Ŝ����;�
m�ڲ��>sI��y���7|���R�áCx�t���H��ȍ?��s�3?�W���2s����84��+<��K�J���r���^E�~����yo�gBN�sc/(8�>i#��*��vA���&t�`��T��)���r7�r�A���F5�f�� ����Ϯ�	?羄4�������RknP +h%���:z���ԗ�I��^�B>$��}�O��q�6]L;�l(�ƪw���m��&$U;!�}����WI<![$���B?!��Dibwl65���j���U؈�d��cT[֕�a�̿�ص#O�#�����ʙ�4�ٜ|����#M����u�ͣ����^�q%�0ړ��p���XS�u%jF2dM�W�˗<�o31��l�2��0A�h��T#�����Y��j�{4ݺ!�~�b>rv�TݚRQ�<8lHGR���ݲ����m� ��l����b%�ةD�F��U�ӱ��j��[k��Ą�u�DY���ac�m^dK�+���ƥ7�.��&�����tVM����!=��{����8˃�a�4��8C�D=G�@�����i$ZD���5��!�Y������E̜��S����I�;x]���*��wQ$?���<�?�g�+���k�aEF��<B!��Ѵ{Ap�IU3�K[���6�Bǫ�kȱd-�.�Y凌�ݱ �w�E2��qB�P���6
�|��l�� ��d���Z|~��v�z�V�7��"�0#W���@��������Y�r���"+ "q�6�Z�L���1̝��R);�A�ac��o1����b�2��x��cT��W�宜��k���[Ѻ�����MǐC�A�s?Z.� ��X�|�b'���*B��~�t��7L���ȗ�S�������9�%�(�������U's;>�ڜ��A�2�V�ADo$ D5�.e
rB~Am<UA���=�X�F7�ֹBD� ��c�-mG,�ٲ�՟H����f&�x�P��`Q��������B��ۃ�wιߏ����9���,�'HP����T���/�4��F�d�aT��v����avK���֑��k�h�Z���
L�>׳�-Ba�;bˇl$b��BU�D~4|��!�o*�arK]'���#Ŗ�F�DDa���%�v��Mq���r9NP_�>-޸��g����ٕ��\6���AT�#.6��ܑ6��AR��g[Ɖ�]�2d�L�B��	�F�����~X��ף��I�Y�o���:LZ�ɶ�E�f=#¥�~Ft����opM}�p!�:�bq�� C&̦d�-�VU����Z�s��ޗ�FG�1���T�k���H�K�ʽd�6޼h?h�Ă��4�E�*7z��R�Ԕ�/�A�j�����7C�
~oϻ���7H��s8��{
V�j��S�#�Nҽ>�Z�b��0�c��L���\q�c9-�kI<���b'20т�lQ*i��m#yݗ�-�q�mh�ؒݭ��ui��e�(h�	��!]�_=��)ǅ-)����BxE�(���%ϵ������C�
-|3mx��B�`������M�e ^ty-���Ib��X��v�����nF�3��X���A�*k 	�1�n|uT-�L�PVM���4��m3N��fc8P�U��-�ؾC���mޭ����E��`*IiGQ��Hy�R�o�w�$�Hv�x�s�~��d<�:r�u�Y���=ty����(��U�Y�rwR��e�]٭���f����Y�@$�vD�Z��@���� ~���NMM��xdʜ������u���{���`��,{e@|������U��o�����f��/���� ���xX�KX?[�E�϶j���3��z&�v@z�U|��T�m�w	��d��[~��$̨5�k��X�_�.����s���͟��.���ܴw�z@�)CD4�|#�$��K��r�;W�{t
���۴N��>�h��ߦ~�1��h�ls2�D9���MԨ�R>�����5vW_#���B��*�����q�����W��dx��1�E�J�Xn�h�ٻ\޽�]�0�RM��B�})�!K�$����E�z�t�5��a��̇ʀ9�|�������r��;E�ã�X3���u�֢��V=#�ᙆ��\���6����Y���A�Jn����+�m08Ɨ`��P!'}�$>0Ӭ>X�˛o���%t߂4��js,Ȥ���h�)&#�,�c�?�6�A5]��2��[u��}��w��d�m��J�Z�C\O���6���4Z�	:q���f�MJ�N�a	�q��m~���'@�k]�U��#��vޖ�}��`��@���y�M�5)�Ge�$�^Z�W"K�K<*�����M���d�:C���u���Ú|n��qHl,�&�U��qon���3�=�G��W�MN<��*f붻:r��}����c�iI���U����ʃÉ�Mɒ[�z��d�'��*4Me_��=����҂�1h�N���tĀ{Ewq�Jw[h>MR{���-r� N�ǭ� +H���EE��q�(��⣞xg�D���R'���̉C�%'�F m%��P�cHe������FV�A]�������kdY`O��/��:�ի��*���_�	)x�����=J��4���0KRx��0)����h����g	�D�6���))�^-�־_�$�frɺy@r6|u�0"P�F��M��a�Ϧ�j�=̿J��!��`#�5U�9�l�����de��/ŵI�:)�@�ɵ��uo��4x��A�hX;NEd�^�޵iL
�&��i��1��DϺ�:SO����jq��UX`��rk�^����ǺH��?
��ܶ�N����Љ�m|����lBٟ	�o"�C���^p�iu�E���Ke�뜶�=h��Y4zV��ӊm
!q��n��g��),�mH��q�QO޽��l���|^��*Ȕ�؇�Jlz�Bhʐ*[�P�GQ�-����נ�0N�{��)�}�	��;�/�r���/I�F�vA�����v+�&[���sv�0V���3��>�VW��T�~rsQ��l-�H���m�W�M��OO�&�ֿ�x��D���k���bp�ҋzS�~��b�W4���#�R�a�������)=!'kʼ���U�!�l�2�Ihdm��w0"-�a�����;g�W���%�.r�f�c���>Ӈ�����W��_q��
�5��"��-�UkS_O��������I�4��o�d  +13(��d8C�R���T�d9�����&#���T�^����?�}KI�q�μ�kC��䄻�� 1���Z�.�v�$�:�t�Cݷ�&ֶo���fw �x��scݤpKbkڑ��@`3���������C��)���(��*���ݡ�H�҃�b6�>�7�f(�Ȍ/����3�e��?i�����Gv��k4*��"�Ѧ�"��X���� N��̶J�L쩗N�Z:ڢ�SQ���'N3�^n2Ta�IPl*�.`e�n�������J���w\����l� �*H]�2+�>�1���$�ta[����H�rv��}�Xr��)gl��-��@��ᳫGHq��!5`�1H��y3;:t"/�2�X��1n�#��S�ݻc��	.f�}������Pw�>,��I��Q�����Z	�
��Q�d��a�Ӆ��C9��">v"��K���`L9PFo7AN�_��Sg��T��?��IPr҅�ʖ�`�>��0�s�_yYL�/]E�Z�.��R�����&C����Gȭ-i	�`��s䄪�Z�W��d����!㛮n�qG�d��gg�(׃����{�'��0�Q:XP�xJ&r�#���2�Ǟ���Ͳf���OU��▱Nt�+�������KӠ�e<?�*���4@����v�Ȫ�S��lq
�jK�y{�䙂�j
�ES�eWm��Ns�jQ�pƓ���)��i�Hs_�N��Nǽa�`9]b��,�CDqi6�Q��B�*��p2������?b�vt�����V���鉯P2��КÖ�2f��>.܁ID4�c��/����o���������Ka	U��K�,T����:jn0����k�������t.���XL����>�ʬ��)�����:[�,�;�_��r�9)�/�=Ϋpu���D?��笥�������Hj�i��Y:����w;��YUg�2jײ���7k]�����\M+�=�*�iL�����;s�6��+J�<�ox F��z�26Ԧ�V\vbX�d�Ҹu���z�6�kFV�	�����(5/v�Fb�~�o5�y��En0	m�_c��!ڸM�f.A�xNӭ� ��'�����`A�YqH���,�W��L�B��FDCW?�̡�FX2��1Y��=�'�W�ߤ+���>v��)��X�f���jK��k�x�<�~i���I�rd��k͓T��eu��UR��Q
�Q�������]�����[���F�6D���s��x/t���9J��xc�s�@P�=��"�_�r^%����@Z�� ��Z��Hre�PA [�� ��TG?ʨ���2��t@e�� ҙV�ἆ�n���vB�ׄ5 ̑����B��iÓ��>~�t����^�J�ǍO�s��C��U���.�~�z[O�H��X�U8ӯ��j�>�R/�_E;��xrJ����iX�ք�Abze�j������n}�=� b4�)໳���F} D�U\[~]��z��s�t��n,#D�|��o�t�-����|Oڷ����/�2O�GC0�$�xd8w�f\����<�ә38cov�z"�PnZq���|t��M�k�8�(ɧ���&5���Y#�AlqI����1�U�^C�Q2X��S�9t>.�S3e��:��Wn�M�K���kA��q�b��	o��%/J�0����?�||�uB�һ^�N}'���4�	@�����z��^�t�e�$�K,��8~�����CN/��n�h =6��:M	��Kwt��b�I[���ٵJ��"��e�2��̬	z�W��C�ֶ��lX��[G�E&#���"�@��B� �S���M��x��Z�d×���������v�֔S�7i`5�
W�V������Ȼp-�Y���"f���i�&�>C�-
kR��2�O�����4%�ѽ�C����f�H��Gs�����bq��S����&!k"b� �Mog�}2���ܷ
���"9���%�(	듌/)�vݼ)�0f��H��5�V`��?����	��k�&�x��I���bQ~'k�7c^ߐ�J'^��q�|N�&���7��Eʖ�3����ױ�(!ϑW�@����JF��'��{��Q<���HՃ����:�1}
_�^.V��v`UA�:LEȘR׌�A��h�%(
���
�(XL+X\����bW�Y���{p#w�|$���(�ў[~���}�xO�^��{d�J-�6���`�l�cqJi�w)��FV)b����2�}��l̏G�RIrB�ݰ�ఒ�|�Ș���{"��<�81����I�X^��4��p)�$��|n�Ax���iyظ/��5;���D��Q%����^w����爮��W%���H�!-��.���\T����7��p�e��2X.
����� t!��_z^�Eѡ���R֠$�`g|�Z��t��Ԑ(�2���Z������_�v:)����DH�p�W؝�O�"ӿ�$<
�:���XǷ��I8��4q~�Ї'}�tH���s��zJt����3��T�@�Z�VaJ�S6����MCZ��3��l�v�TO���`���X��'C�0;ԥ�'ӭ5��ڦ!������#�0YYM�9��:ꁰ���,,F��|/�g[+?�$\�O1�v�B�y"u�ա�-%�$��p�o4�kTt�s���Pg��{]�t�D<�ƳZN���L*}�8$\^� H�w-AX�??������۾}�O��E��n��^#-*K���hV�	 �i'�;E�')��7��Q�O���D��k7���k�3��i��k�-!�""!��Y� �t�{�%���C�H�nU��a �u�b�E���N	=e~���f[�ʳ�@^����v��z8hɠK����"?*d��FS]��Hߥ'W�^�3 r��s2`��La�k����z�JY���8�=$;���Ϭ����忷�6I�G<95%K�Ems%�!�l ���3�{r6����6�}fX7�#�M'��mu��d��5�}�/����h7[}��P8x/��B�MI��k��a ��΀ޮk��E-�a%��ěǷ2<���D�Ǿn|��w�%�]R��R��nԫ�Փ�D\}��96��G%W�oN�t��K��ފU*]�i�^��@8.C��m�+V]�1U�M2�]*�~��z��FV9,�j�ֆ`�X���p=YWH�B�Dl�X�ު~�\]j�M{���P�_<+� 3��<���^ՠQ�E�L�Gb�lu�� h�D6��;�|&�P3���1$Bn+�<̓�MU�@��*�W���D�A�A|Ȳ��þ�o+�f���ZX���"9Iw�A�?c���Ż��ՉF���a2~v� QV�g�r���[�=��,�e䔸����Ȯ&�;�d�n���ּXG/<�]�ވ8B����h^V�����<�3���*�~��%����\�>�#�m֜lsR�׃}1�_+�"��9c�Ìl2b:P����}�#{�1�Z��Ɋ�WsI����IT��)xp!`x7X2�P�2�^��	��3��!2}la��0}��}!#�����NP
OQ���ء�=���U��Uld�`�*F��3S�bq�$�@�DL�T�$8���C�ـ�&?��!n4�����K$�@J��V�Dŝ c�?��sG�y`g�����	�_%�Ѫ|xg�RNy7e޸x�٤1�h�����V��թ_C���{y�=�xpB���<w���E���V�#���Xp�>��ʽ*a#a~Y:\wazTO6Q��w���&25��G��#�T^�
�17\5j<��Ռ3�}A��D�6��z��H��)��%&�Wl�
:5H&Z�_C�t���g*�@gTtԱ�`'r��,�6�M��H�KS�{[;����VC����wm�~�K��3{�`,B�^<�|�j���@�uL��1DD���c�.rl6�������@FF�ø:�����	`��Qtj7���S��)����ږ���ĵ^�6�
�Τ_��z!w�B�#.�w��#aV޷ӏʅ���Ea�dl?y��8���m �7���݆���ߠb>�j�z.�� hi���۬��V��-	;��~������a��ۏ��񏉫[�@����'�Yؕ����
r;K��U!�z�ͥO��4��|�O�5ր>u��kסI�x��OP�pc�)J�0.A���R��;��w���T���s��MoV.JQ��(�l0-瘬��T;+B��w�n)k;e+Ï5��Z�N1�X���uE���
�/�$Ľ�~��I�`aw_�}��͉͋ad׎��]��ٙ�B���t�~?�a�\��x%n �v��g���k?�6F�f/�I���H������soJ�N�EV�D����+�����H�!:�
��wr�@vN�p����i?����9����8p��O�{���Q�TR��ݶiӆ�4+l��̫"�.}:X&�����!=�������-`���� P#���_.ͥ��n���ݾ�������hZP�P����X��䄤��z�\����Xj��҇/�N���8NH�yI/�uM���}4����+�?e��v�[��"_T��--���|"P�m���vS�>��jq�?۹���s���ΎGeb��_���Hu�l�uNG�*3_6�	��1d� �F~-C��3�ܑsꤹ�#0�l�;z=�v��m�<-���:�Z_���M&;�� ?�N��e�q/��Vĸ����a&�Y���B�KA7A4�DH�(S8�J��A^���z��Q��,+O#��u;�ܫ`Dd��3'���JX+��N�����_X-
R��96y��#}���]B�n��3�ޜ��#��S�f��Öl�!X��*�}!��`T%Ĝ�ǖhdOہ�F�OD�gd乗Q��]8��{G���wZ�<Y>�e~f����DҴ���(��x��`;���VP���^����g5�Y��ﾗ4�f�w-�j(E���[B��R�5���DLzW[|�"�b��\�� QR�E�i4����jl�7�L�s`I
�/ٞ�bjC�k�*�Im�/;���,�Ǻ�/�?�gfC�} ��S�+5՗�����Hw��;e��p!�&+�E���!�ғ�7�^f"t%�O���>�N�(<0���I�Y��r=�ga�o�4Ӝ��<mm��o	XtCˇ���5Xd3�����Y3 �L��c��^�²Ӣ�\E�d��I3���ʈܡn�N�UɄl��،��g�Вӊ���{�s���A���D�$J��0��k׻L�JJ��lրY�hُ<[WH*�5B��oI_u���6q�c���.,�`����L/��u��	A	N�4$Ay�Er�@�~ߍ� �5�� �������А? ݹ�#�JFnSȹ*�Ş#��{�D|���Z�����q�s�S�2��1�\(<��0��+�('@�&l�q�B#�e�q�7��R|�9,�S�0�\�_l��a'�{&D��������ޥxW=�׿�<*�8���0j�D��K���KE>1J�mq{Y���c�
2Aө'�#oř^4����|頫N[�c�F}�S���%}3��Ш�ߠ��˲U"G��I�83/Uo~��o�3���A]d���pdQ�h��Ӈ<?�x���	�&���k+-�=���ڟ]�=݀��L�aX!q�s���&�*"6���Yl�3�9R�xg�p�ݾ
��Kg�<�A�緉ynzL|��F�,&=y�$��2_L�=�=3�@6��!1r ��nq�ֺ�Kv��b1ţ����*�Jh���r��3���M�@d�k񽞹���.��l%���iʓz�G�#>���c	����ق�h��G�w�+\�нn�[�Ӽ)7������*nl�HK�įD\=f����DH��W�t�s��KʌzA�Zt�g);-\h�ˮ2����� ���.�I�7��\J�ߚ�*�D�ƱC����� ù� E��R�h'�:�m3���Y�z���`��G_<���WIʡ��)
�E?��́���x��rQDz��쑪۲��p~�xN݂�afP�,0��\�e����3^+`��X�W��f��]��)��1�%D`x�]���-�E_��#V�NZ؁m3e�/��E��I��.�)�-��Q�G<P��A��,��ǧ���p?�N%�w����:���u3��t_��Oi�2jfw���7�5��"�D���I'j���`�Gh�#�x\aW�JD�o8l[�*�Ӏ�Z|���������-��M#溁��:r�,Ȗ7��?��f�$D������L	��=�m޹��8�� h�|�^7��n�4���8���S���]����Sl���%��H����ӑ��A=F�u�C&ב_u#��ư�ٔ�/���都��Y�����f�Œb��-���*a�?��)�3��䂇��!�$*�c�]8u�>�9���b� ��up����h���6��Ȧjk\��=���DK,�j���� �){~u'J`�6���5�H��<���B^`V䑠�\G���B��ү�Ծ���BU���4F	>���an��ƶɡ_��a4p�)�8[�W��R��d]����CkYq�����X��Ȣ1������$[y�D=���#�Ao��)񢳌/A���y�OuI�����Ȋ����?N��i��<o�M�]�< �`Bqܱ�W����Oy�a��8��dzx?W,�Q?U�ՈL���g�}��щY��'|?������F"�C�D+���d֋��a;3&*�/G���c-/��Q�H]�q�p��NuP��iD�B0nY%-L\�ˉ�}�;T�d� 3n �|�
��`��uAl���JZ���M8�b:ŵr5@�l!�� �{iD��T��l��u�O]�s�&��w�L'�V d�Ӳ-ɻ�X�(J�V����߂�9w�Py�80®�4�x���2%��v�t��Z_�!<E/,���+	O.�_�x��yQm)z������iu���j�\z�x=�i�A�H#�k�/��͘���O�6�Q]��$�f-����I�6~`�F"Aj�)�z��B�4�5A��ћ���[LR��^���*O�u��HE)���j"�J9���'�@����M������3�G3!N�;�\:�޹�_v;��͵�`�m�����K9}�����sRY~�G�
j���v��F���i�lz��|��Ya�	�/���iH��t��n�2�.�1��Gn7�䶗�"_�d�g�j��	�D��m�/��LM�[��qh|�7��M*?�V ^�실r�`��*σ�1�0��"yқ�+ջ��'x�p֕.π�#�wk��Đ��H���+�=Ԣ�\[�� XB&a� <�K�#ӱ���]��o"���S��Z)��nd�C�]�9H��ڏ���EY�to����F��.�h��E���E#�*�h9
�y[��J���;;�TnF�S)��:m���Ń���#�V9E�]kVդ�254�j���ҕ����ק�ʕzUU�����y����&���v��!!���C��8�t0��x���
�{FW��, ��r�U�MU��g�^��t^J�kV�����\�ˋ�(�.��9k����F�t��\X����6�<����>\<��ZP�5�P�5:75���j�]�b���n`�;��]��p�2Qwj3�Ͽ���[9��8���5$���:ti`B����ړ���Y	�/U֒�R1r�-��Y{译��8�*
��<����[��
�*舏q�ߜ'��޺�#$>3]h1����-�i'����7�8��[�N����J�r����4�H	A|�1�@b���(y5s�[]y
�-q�I~h��R��X�E���QM������!��v�]e�&�o�[��6��O�x�8����ߏv�m�����d����5U��E�y�[)C������qo��/�!ZJ�7���'DY"�A7"f�Kɏ��=�2���|i�?oJzĊ����`s�mRu��8�M	�=��us2�=Ǥ�Epu;���&�֕�o&�̟Y��cu=�[k�j��,j���	���_���^�����4W�$b[��S��4В�V}�����ˆ��s����RmN����5 ��ƛ�瑣����n	�a�p�?�ء�'�=��e�4��z��\3��G�د�˒�����o��NoG�ٿI�Z�ߜZ$�S#�o6'����GF&��dT�(�τ(�~�i��8�F�p�q^���ͩD����L�Q�Zh�,�^"y��y��t���7�L�[F�5?��ZI,+X2j�~	 ķɍ1��T'�>�`Ռ�.���s2>D����g�@�=�sk�3�6(�/B��2G�˄mj%����
F9�P�)�K�%��(��CU4��(t6��EuѓҺTn�J�a@���3�փZ�*b e��P�M����o��O�+a�V�Xϰ�'�!�O�G�5��Ln���a�n�j�Z����dݦ+/BN���a���!i-R����}X(p>�28mc�6�4�5}oXE�
F˨���s�6 �=��	�>�*c����x�QZ��瑎�Q��4�� ��S� P�	i�q��t���Z���e�&[�Pa8��lyGzsd�F�K����V����*��cà)3`u]��@M�/[Lq;ǹM���Y3����Yb�q���Ӗ�&P��0��F^��qp�ˢ�x���f^�`!�5����3�*z���ny��9�.?̤��>3o���r+S����{�T�e~2������`B���G��~+��{����l�׻�=�E@?$�/����{���ˎ`	��
�2�/O�}k#\aRWn��$�KO~�{F��뫶�>́z5ʢ��T\�>�$0�K� p���?J�	vr�χ����ĲH��F;�C�N�n�!�)A�|�:fi	J����MNB��.'ƿ� �>�/<�J�7v�?�}���xl�����0�U@Z6��%��*zI�eD�}9Pe���wX(�\�Vr���_��w�%/�l��vԮ^��`'��2ѩuOO���P㣑��FQ�+�7����VAc����Z��a��������GM�x�2�@��#������ڜ�\��	��BOai�7���4$�46��J��ժ�n-�;v�a>�I	��}@JFG'Q�r�f��Z��7L�<~��t.������Q�HH�w!e��,CcIn\Gϖ3��]����j����5���[Pn6����x���(6US���+�$i0�8������sz����c*vH)��Su�6h�h^8����+�"		?��W$�k[[J��M�"M����֔*�D�V�;�+5V��dҖ��e��F{�ǂ-D�L�cAQ���!>y�B��`�I�(�]HQ�O����ӯ�)�R�HPF|p>���pUCZ0����$����5x*[�K�#���x�A,Cw7��p�`�ڡr��l3^��de�C&k�|�uEy����.Ȁa��.�q�^fo���Zi�����|V��k���qJ����7��ǸIE�n\�6Tf�\	x���vO�12�㚤.*E�_~��B�W�4�z6�[�W�.�~rIT} c6�d$j�� ^U��l���	f�N�E����Q�
�����췢蹦"��?o}B��y����2��JE���I�a-�s���S����B�,^5֗�-���@20�|,Yi~_��'h�z�&���U	$����b*{��o����n���Ċ+�sV�=߾�8#����z���$1�4=�.4u��3pu�f�-���'ŐB��(Io܅'^2)>+Q	t�@̦��&`Q�r	X��1mK�
�+�W�e�~V;�������uP5;��>,���u�x�O��8��o��l�vԢ-z���i3��͢�	��[Wb�����	I6Yj!j�������eW���i���/i	�IOVg~%���7G���d���P���_��gaA{ð�f��	0l�J9V��K���lŀ� �Ңއr�2���τ9!����Ǵ4ګnS�SB�>�I���*E���|F�ܒc�r��i�"���E�iqE�'~�0�8q���]��.�ȿ.s��@���	��_��V��Ј�Ǽ����8Qp}��\�]:B��]��)9�� �]�u�����ω�2!��/s�IN6He��s���� l��F����*sk����S����Yؿ���*�2"W>�sw���/�N���lgYKF�!�6#:�z9�ߝ��P�����ܿ��e+�D���C�t08�X!À������x�20�
R��K��D���9|D.�T+�{��S=P�9M,�ٴE�;� hj��m�%�L�.�(I<�G7���T.��0������Ī���4�{�\B�����	�б���F^���e>�3�p���
�*���]�V�����#F�m����:�8	$�u)5���i�N~���C�,���� �H�Q�/��y<�h�<�CaҚ���Ђk%��P���5����� ���RC����3e�4dI����j[���t]���G������@J�)l�l6_�Q�A������kF�m�$RJ���U�{�9�(<^���{v�:T��w���t�>cr�	o�f�l�1Ȫ�B����İ&AQ���#5ܣ 	�y�}q���~���1Ӽ=�zA'{R�M�����$K����HH�����9�/9?���F��^�8���j4B�^�eH�����<Q�I޾�z��Ћ29����	u�ұ۬��i��`P��`���	�T���0������$M]�.�S�j~%K�B��$h�u<6��h$���aQ���%;���y"b��F�ݕ�֙'�D�wZ"}Ɂ�v�{ך�LO�3�������H�B�_s轈��{�W�Cpy\��dUr��+���ŝ�G�"I�<b����p��'����l�
�[ީ�q���}����
������`����+�}`��}����*Ca1d�KM��߬U�O�!Q��prj�q�6�x��*��@Ȓ��^EZ��_B{�XVț:&�3Iۙ{�ǳ���GG�N�U��Ѹ,�@N3�u���>�}�
/�Ō�T�y��|�*��JNr=���d6��SF@t��� ��$�B�u�i,�+r���=%t�'���C�k�� M8"����atc��΢ۦ������b�K������<Y^���Ɂ�������PX�ȑPP��"��jvڭ�/��Ȳ�R��Y�o�9k{�sHFy�7�MF�)�ݞ���g�ݻ$v ��&>��׎��N|�tӃ�,����&�
d�>�^^fj6���xR���b��0�%�%nd�Su���R�@j2ukzJ��^��oc����HWD�Ml�rEI�^e�d��2w��Ȧ��.*�'�S��h=_	,%[ʋ���/��t*���"����%h?P쟬�|���ݣ�A]��+��8)t:>��@����Ć�kɴ��,�d�4C�ñ���1�n�&��5M����|}�x�J ;�^��y�ҭ:Hա��{#�b�b\���1�L��C�r���<j[ee��5?,���Է���2�o��9+A��M���h�Y��:9(w��A K�`��~1�)�ݣ����*�{}r_1���>U���#8�/�O��P1|)����FV\�*c�vR|5'�%��O"�B�Ⓑ�������֠���qf=��u64[�x�j� ���^���f��j΁�h���\�=�S���
��w.�܁�$�	͢��M��7���ɾ�7�
�B�v&e~�����}��P��H�QW����7�[�Id�L$��Z>')%�:F�쓯��!�x�B;'�I<�Sw�倶�V}R��D ц�Kg�~��3�~��P�&
TCQ��L�Q��U�����#"
�kv4���y+���q���!�OH�I�g<3�1��)N��F�����<Խ���K���?�1��)������A�Fj�{[kV�@d�h9�	�~�&�����d��n�`��9 b��Q���̺�j|�����t�x���k� jc�ޙ��%u���hkc����""�G�w�C�{�|`�S����ȼ��tC4f�I-�I#_J���)=�Jj��w��{9��ů6��0Xegv�ot@�Y�Fr-���/`��P�hޞK�8�yv3>���}:v���
���kѲ�^#M�%dfC��`�HK0��W��U�7"�9G/�u�.�Ϊ5c��PFO:�d�9y��g�WX_��^{xۀ�,��Q�kK��r��R5�1N�'3VU���g��IۿϮ�ry`���X�J�W���L�i��>�g��1.�$W����џX$8�l\5|���u�t�[W�������y:�J�/�^��fdX-��Q�եұ|�������Kҁ��=W�Y���+U�k��S=ӧ�I�E��q�h�	ra�'ɻ����4��ux�ウ�\fqNs�,��6s$�uVe�hZ��8e.�"��X���
�
(�F�ϴ���>�/�,��.��M�2+�^C�;\��!�w*�l|��k�yE�AN����+���s����-�����?EZ	����;�'�[��1�W`FV
��;��G�/��K�[����G g��/�MC�pY���J�]-B�/`�:����!Z�W����EO��(���,��b|u+/G.��8H����h��ДQ��A��M*�2M�xұ۴D�}2������W=��{E��]�ڣS���}�P��9�L�k[Y@��G1���
'��j�ŚN���Q\�����OQ�K�]��2�D�(��W���n�.��/y��� ��YAH����͘��Cn�&�x�T&f��/ �E]�/a-�6��W����. .|Ϥ$l��A1�l���N�n�Dp��ulW��(�>�;�S[�K���I�Ӻ:�����#����$
�WS&s�;5��-XSk�:gI}�ߑ�<)*Q���BxRd*��:��SJM#�P���~����3Xx	��"��Si�7���D�E�F���'�O9Y�D�A5��x��>|jE������v-��:�<��_������H�g�oK�h�׷�=^Qד��O���̘[�5������9�M�U��Ä(8g��&��[�N؟�Jѱ�Am�4&�6��ktD�ۘ����R*��A���t���a�u��xl���I��\��nYt��rFB�y�� ��y���� ��y�	����C8o�Ƽ�SՅխM�������.v�{��P���_I2�S����Y8��s`�Ula��@������Zkj>���&����t���z��9oP���]N'	
^�5� ��e>�1���:�g��	���|���("6���N9������51R�c���wk��-*�9 �7��M$���?]P��oN�H��G�d���:�Kn�y�pOO�\U1m���j��Yd�����D�Gģ�������!�{�X�-��
!��Ǉ9]h���)��h*�wl1uK�NJhs�����U6��/�Hܺ����i3�+V�����^��Z�o���ʤ֎�|�� �y���2�B5���G_�Z^�lh]c�b6v�����4p����ۼ͉:Рf]_F|ǈ�[ܼ1�Il����5J���@�;��v`�h	�A�OX�G�c Fˉ��՞�$����J�I�,��0|IB����t�r�d�՚26�2`<���}����ηuS�U?���_�l6Jl�����RB$��0ҿx�PbS���q���Ы��*&��`|�� U06 +��q�J��0�-�a��RRg��0�~H��Ҥb�.�%����Q�z;�{���DNR��r�3���}L�-C�^1h��?�Ո���q]$�E� �%�.�{�����A'�S����{}a�Ht� *`��.d�_�,�ga��%V>E׺���2���P��J�ܯ>=����O�^�j�L<�ځ�0��Ϫ���dx7�L|�>�ǻc���hР���m�Gn�Y?���1`e���Eė��s@�`�țԉ9Ć�����f�����+��h(�Ӎ�<��)�W09�&A��d�E)��2�3�����y
?��a�t&s�d��}�}��U����j�������������⛸:/*�Lm@���029"5�r��V��H7W���k�;�Y��Lc��h4�Ĕ-Y����?���unL(��g�HQ����R������Ո�d.��e�"%�,���Ӧ1Z_WZ�_���-�e�� )��f�A ���˭��Q*`��ܖ����aW0��.��<}�BPf�Z4d&�rD����F$S��ގOv�z��:���K'��(�煆��9p2��v8[6c/�X��=o��P�5��Ϳ�ݦ��o�3K%p���ݧ�1�,�ԅ�{��BF����j�#.�]��
dW�B̕�x�� �P\o��V��{RQ[M��9��}��G�~$�3�I̚��TF�tkl�����R���+�Ơ�W�������ߔ�q�$��F�~ڬZ�$�I�?��9�)ҟ֚a�7\�%��iOl�/PS]�7�x�Z�*%�����fF����$�ǆ'P�:���(� �x���^q�Y5�2a�~��b�OV�F��[ƙԞ��D!��g)R�;E�/�Gl>�ɼPA,��)(�Of��\A�?�"W<���3�c����M�%۟�:��h[�6ǩ�:�ҞLfJy��c�u�g>ߡF�]�o|��@�+9�P��<�_��~��{u�_�o�i�=>ҪA�r%�o�6"m�nF*Jn���-��Ⱥ�}�-�\&��'Cp4��:-���Bv����4��k���
���9^y��]y d#�����c���n�J=#��$Xq2L�m?��ѝ�g��Eų�:�/��a����z��g��_���Z�X���Q�z�N�k�MT��T1�	���}i��95l����5O�E�����MCt��O�A�IV�L�PS�t�y	<�H����T��Q%8D��C��u�M^w���]���;p��M����	7��`>ٔ�`w��8�Z	��M��9:����/?�"&�O �"*)���	GOt3�L��}1LY�9��	|�5Hʥ���S䭾����<�\�[�&Z(��b����V;�JS��H"G���n�]��ǖ�������,O�7�~&r*v��fҚo��Q<a�Z}��*�zJ��F?X�5T���'�/�DpB:���i�!1����t�C��d]��h�G�O�#�<K��C�U_��N�}@4�6�>K��L��zr2D��r�^�5N�o=�E*&�4l ��u��b���o�JM���V�����)+a|�p�P޲3c�&=*9�A9ԙ%���g>���{��	�0�J��w ��z '�#q�:f�1U��h���} /U'���7�Qz�5� ��Dee�=�
z;S�d�/�o)����)�ۋGzy
��ľ����foso:}��r_[��Ʒ���W�{��z5���0ȉ>�8D	�;��F�/��G����^�}	��fJ��|����:�4ו�!CA{����� �3U#�.@N,���>��0t�~��[���g�+
����<K?���G��c�G?!fQ�*&Q%`;�@̳��i� ��J2������{Ci�y"�b��$,�����+}�*Y�;3ha��*�L�,{Z�ZH�*�ҿ�ͅ��t ��v���΂�)A�8�h�nQ3K�����O�*���tN��nq����g?��F�5
Ȏ�G��c����Zs�{N�._����:{�T��p��$������%M����BC �}���O[&��r�TB���EƋlL�A��2����o������g�<w�K����6���B^�D/*2��Eq�k�x!��>���[j�T�虇�L:ɤE�uʨ�lu����Q�`��C�HF����=��I�4�D�~:�	(��`УC|�\�r��fn�p�����d�ok=��K����[��K{�N%��䕋���㢼e��H]��\�!��y�%�$W���#�t$Ч���K.�]�vv�����꼊�J�D�`�6b ��'3��Ha#�8N{qĕ�f�)(񈺭�U3��wMķ��l��\��<"�}�ڮd�5��}��t%5*)���y� �:��ۉ�]�%N�z�vV˼[�Ӓ0x1�}�cV=��JЁm)��iMeĺ�X�JK�o[Ԃ �w��q����KX1����ϱn�Ѐo����^d ��䓟D���S ��w��d�ͅ�I"G�ac����j��<����P+��nʬ��'��ܙn���cm>��]�<�����eI��������l.���<b|��<O�t��1��
��~eO�6]�qjWQ=���矶��zq�D�p;�*��i��rjE�jDH*`�l߈T�^ʵu�� ���}�*��H�׎tW��TM�Jևz�ZD��ʋ��(�O}����ǢX�i3�*Mx�V�JB�ɫ&���m/��G��Yp�d{z�X� ���B91�a2��c�2�դO]7�Zs�.�:/��vaOaL6���$��n�Ӗb��&��c��ã('�7�����w�+xk%�z~l
/JEQ�+i���ݍ����!B��h�Rg�����`�D�Ӛ���C�"����|�����PE�uT�xhw}��!KB���`\�YXc�C��w�x�N�b��G6�w��'�}�҂�?cp�Ay�tqb+ǊKёo,�Z�Fl~�DK+��;ng\���c'�ׂg��ITa/e"���#�"���Y��CrZ8���X��"k��FE���і���̓RA��;����@;��:�?Z$��6�d�>\Y{@o����d8"V�W�Z�x��"�@i���U�V�8��e�n� ;*��$�S�,�e��O(�i��������I�O���|����X&���{O��96�x7I�/S�VN�Geo�F�U�*�Y�2Y�8z�WF�.�?�5�8�{ԓҚG��&u��Hrrs �O�4M�P��s�R���TD�[�̞L9�����h'�D�X�i�/�/��z�\
��}/�2��jl��`��h=|ƻ�n������0 �[7�v�(h W��34Lr*8�pOr���Nt����aS1�y
�u;Ұ��Ѷ��:m!�r�R/EOF�;_��,	��A��E4�¾�S��U^}�U
 :-�Q�����񯧹��O���������,$F��Ы������T�E8�E+w��*Y�8�̩B�NZ)�0�\%��r�C�k�>��Kn�^��V6�yo#��,,�}B��AnJ�1'�R�GǻW�35��wY�4��Sa+\��˕��������0�rGfޫ�e���-����w��Gr��
����������D�Ɛ��uZ�[;~��F��}�loH{H�y���
C  ����V�
���c�Fg+�@��y'�����Ip�h�0!_�o�y9$���/��r׻��SP$��bG�����>.����@|��-����+��+>H($�Ê�\$�0�߽����#a���R@d�@IRw�����K��ٕ��S ��P���v�ɼ>`�!�-� ��g�|�R18VJ6 Z�u:�݌-4mƒ��U��"<�����FC��0�Y�#�
�W)��7����r|?)�J�W	Tm���"ة+6�R�$ܲ�4A܅���t�P�e�}���0���S༯�Cl�?���&dI��y#��(Q(![Z#�Wɖ�V�cݫlh��/Q7:Y���X&����vz���HQ�׭����?��KR�N���^�4�S�"w�ާ�&�k��X4K�*:���Jz(���&�aN��������QސY�������Б��C*�������y��$��Љ�X���7�]��XX����)�+�*M�q8�~:�AV�{���cY��(I��]��@�BQJ���q��e��w��S�)>	�eA��ҹеz\�{��RJg���(��N�]Ib]�����{$�	��$@�������ih(.s|t;�� ������,�����R]�V4�:
�(�n��K���7���g��F~�"���|�ƒ�>��"[b\\��-�,k���e����DV\�����1]�@�s���-����^cڱE�O�ǘ"�n��,?3m�ᔈ\�禍!ʓ}�U�R;,�;�_ٵ,��Z���,�?̮0�&zO���6}/��[��+ql�Sb��J]�(�{@�Z+�Q���r��0���\���o��	�U��?&�b��qb�مvlU�>�)"4�����<�_g�^j�Z��O'����O�tf����y�К�x����-zP:h݊���q9dvWHf�u�� �\@C#�d��G�<*#�t���K�'0
��f�3�3���Ò߾0�2b;�蝹�ԙ��Q�0��xqXO`��A�,�����b��Oy(��Nl�Hj��ŰU��)5�K�K���O.����ʠ����$���QB�7t�|�1���y�DzlU'?��wm3�0�b���&:�\d��{\�ͽK���=�+ԇ�r����w�l�������P2o�!�	�ZW��y�(x�R�i��BV!΍[l�r�����ŌQ�g����#N4�R"�-��>Û�?Ǔ�\�uDG����5���w����VF�T )��9 w��ծc���FٍDB�\�"8�:�0�0��&p6m|���u	���z`.ZsA?n�4�JՂ݇r�G��P��G�ʻ����E�0.� ��$\R�b�$���|��3c d�A������4�1���P�$oQP�F��=�d���e=.ty{T�����>8b�О�y�;�#k[v!���J�~�a�$��>.p״��J��.e��~����ݠ��#E�!�%Z[?�D��_�-Vʆ�<q��p="L�������	�sbR� �K�G���2���	���kW>�]�#�L�ÓR�X0����S95d������j;>*\���7�`��eX<�w8~�e�����ۍ��J�$g+�eq�dE����4'ՠ>�F��unT$`��{�Cv-ǄCj�OU�]j�tu��`%B�p	oo!<�ci�����z2�S��{�(��g����ߟcٯ���������B���N��?W�Y�m]D�f�P%*f��0�[g��>�v�ô���c~d��eG����Й�(���n=�ӎ�lF�lQ��~�����έ��8�0;�v�M�6G�}��ic�6.qH+�o#T���!p�������(��r���f��$�cpΙ��n�ΣJ���۠��c�P;���=6C��I�rs��*�j�"����ҭ���Tmd�l�io�����?/���oz�~`� �/�8=��Օ):��^�^;�3 ��ҧg��ͺ�/f�dt��+/9W0�\̜|㬄�
�����c�&t��o��u��")��|B,��$�G�]�����Ԁ��K���?��i�t�{�g�	Xem���C����9����l[�m�d�x{����f��v�yH"�ՠim#�h�L
ٱOsQX��:V��B2.�3�Ҁs:����g�4o�M[)�3a,�V J9zxv�UE�m���9.�/VSyn�T֒��'��B�4
&vV�FA.I[�u9D;�m�|�J�L@����Z�~R��(kfȄF�b�U6׆NE�J�5����#��SM�n�3s�j��dЉ��cŁ�5M����.#���[��b����M ���98���E8P�*i�Dx��Sk��T����uq���� 0y��>��L@�1GDB�T� �CƜ�d;DuZ�Wn`a�����4�i2�����}�K��:�(�V���B������L���F�ҧއ�˯�t��_[��q�V'���1]HsWK&���޿��<N�v��:?&��_5�h�U5����˗�Q�g����<x��Jȣ��2�d|��C&�ǕH2�.��.���N�
����$G5y����l��B����Ԑ�c�o�6�JH���F�7�ٕ9u��F�ɽy�^s3��V�Ե����>H�����.��؄0���a�������K��y��Ӡ6O���96�r�~Qpi+����?vU��tB�f�<�p�>�a6 ��E2� D����2Qo@�@�����ΐ�z�:!=.Ph+�, �p�S����u�l0*�`},��쾄'~d�3��%Iu3��m���u�ؼ��v��e*g���-ş�p�)n�~�z~���f�� {��k����Ж`!:!�l(�x�;��
�za:'��$p���]�a�\Sً'�����>��=�Q�b9�=�{�9���x[� ���-�J�ӧ��vk�Ϗ�j��M�"� ��0�.�ᚱ�نذ����
\�_Na��yS��⹤�8EaQ%�l��S�~��3���0P�����Г<"�l�$���l��	�`yg�<9��
���'�����[�x�=��3��QLV������`���q��K��K�Y WW���[���ǋ��	T�����^����F��L��Y���Lez�8�#�xuz'��C~/����]Σ�f:�E̵�3qV�@֎g�N�UL�0��0�Fi��{I8H�L��"�>���Բq�3����c}wtپu������PCu�K�1��i�//��E���!��Cg��<9T��H�7dTO[����V��ܩ������mؼ�ϙ�1ڀ=<�]��H�s�R��FkY7w��� �U�!p=�]����Ův ��-�LxB����M��l��x�g������ќ�m���q�^X����1'�s��+��N���mVnP���(F�c/~�M�F|����5N���A�v���P7��8ڏ�|F�[#���M��4�|ɢ�,����k�Ѭ�@p��Bl�l3��[!9;u�؍C�]���[�
n��S��w��п։>�Z�$/���L,PF�&D�=
�ߚ�Ta��5,�1���0OS������w��l��xQ"0�j���y(Ĉw�gZ���y�f��	�Y8��m�!0�z� Of?ZA�&��$v.t �>������ǯ��v��%c��hԡ�C1��^Qqj����=p�X��tܸ���';��* P�2O�p�J�!�����u�%k�(
R>�k-mZ;�̌��_N� i��1Н8?��cM4 .�M��;0��+�5sJ�e=�aLW�A$�q���&�HWw�F"rC��jO����p�h�Qs�]��L7ani���<qQ^c���쐄]j�g�uVm得�3��d�O&l4�$V ��K��k�'{:���k��G����kG]JQ,�9 ��@ʊRe�⩏缈� Mu�ed����T�=6��{!��Uq�{F�=��|�;/`r�WoLU�V����Q~9��� M�����{Id���_B{��=���S  �T���6���,��q`JF��""e�gQ#^��C��@�g&cțTy�Qw���ʯ�%��Q�Jt�0_�7��2��j�2�I~��&�7�6��D~�EF���RQ��j����Y�cTK`q�B��߂���zSP��jV ��{��KZK[͏�%����=p�+C��i��%��<�QW]�߾͎������>���E�k�j	��צh�%a�s
г��}���|� ��y8ƣ�b&��26Fp����C�� ��L���6w�Cd5!����Z|�������uiF2&}!�l��o��fG�
�]�����K����J$u��z�'Xʲ�9~�������PF��M;Sq
n�����.�s�8&y(��t����z�C�Ź���-\`%kc�@Obf��$�֡w��ܒާ;v��ҳP�hTRI��O����$���yɿ~�d��M�IP��zAm��M9�j��L�&v��Px�^\CӔϑqU��p��W6��3�Ħ��+o>l����FM+�6SL�f�D�ol�����7��h1��.,��B?�������C\Y�.�����e���c;i�Z�-X�x�jj^�i�2�d�qfSM��-��y qt
h�+!���wў>��Oo�;�7�$��?�K��9J�������L�y`��=��L�ϩ��)�\�63��)�8�!��\tn��	n��Cʂ�\  �I�$j�d��)�h �M����|�v�l�� ��2k���N�g)h6���
����"R�����ݸ�~fR�2 �*��ޘ�-k��w�},ݙw{zIڜ�i�mᷘ�;q�c]��u��*ǰ���Bֵ�V�3Šf}/�ew�a�18����ds�(��I�nw=y{X���;����Wd�������C��Ͳ�`�j�63�a���a�XgR�U���3ȅ����QK_J�}��Bbrx.M��.ᰰ
t㚩�T��W����QO{�����~9^��˦6���/�ٚv)��_}�
fm�UkB�&2z�9k����`y��	Ѧ��E�0Zt�~��u��:������PJ:̢���uacv�
�P'���r��; %ݳ�r�C���il4��Z��1 M������[�]�{_����o���*�*�0z��+��!	��y�<>����^����d��?�+�pA�g�E*#����p Z�g���G&ok}��⮕�����v�,J:�E�!��k������kazs��SBn�X�K��Ҋ�����ԗ�|!����u��xT0�!y��f��G������=�++��vB�i�~�l�k�ڸh����D�\�a谜�{�q�ޒ�E��xP�@�c���/7;�L�tD��@������0z;jkS�%^��U]I���6QZ�_<Xjm41-�N����4+\�_�Ǥ��1���%	iQ�$�AI� � ��13�V͗��Q���I��͛�:�O��yP��`ں��T�̜���<��[�����e������4N�ԙ�Uz��m
����/�ĩ�ݓO0,���`�J���/ ADs�Q%��'�`�ݎڔ|����x��W⮴���d���K�v��B��b�eʊZYՔ��?>.6�=�z�ҕ/k�=������n�B�R�Jӈm�$n��7��W��?�m�i�;�+�-<�W���* �'߰�bU�bӢ3��"�m��b5��k���#�f�q�.(�5��T��e0��r�!�Gu1�L�z�ۉ,٭'�%���{G���o^m11�J�.�"��Ujꦟ"��X�>��<]S����5W{�##Wc��	�V����bXψ+fѸ�u����X���b�I31�	�L��b��b�W�I�k����T5���8`e��,��/��W(�q�ss�*�]�����(��n�8~A���)�����9�!z��/6@$�<�청a3���J��)G��w��ڎ� �z �۫=9���[-�g��k-ݲ�y���rt�X���I�B{Yj�f�]�-�68���cte��Ԕ�B��I�-?�%$c2�bD�(^j<��*��K�	�c?��H[jQD�"�&�	�^18��x�"�
T�˼��G;�-$��tf��������dt�eIfg����4>���"I*�?�XQ�{�&�mM��p4�T�)�|�s��mz 
��p�X�Z+�*�-6�����њ�٣: ���Ϳ���v|���]�*K@p���"7 ��e��ݧJ�1vի�5�"�NX��<q�\�C����p�n՟���)�8�b��:gIV3��3z�%������u����.ȶi��C�n
u5����b�:��%���	�C��� �K/m��[.;;����L��!����_�	���v)�fG�^�����%�¯�˻tS8���%M��g�-C��so�ޔ�z�. פq�"���	];���R��ۏ134�O����J ���Gc�]�t�c�ٲ��P��*}Ru���Z{;�jA�0!�t�����1�õĆ�@�uݗ���Kk$A:N�Ń��U��K���m7b���-�h�,�UG0��Qh�Ye|΁=��ա������li��\������ROE�')G��Us2hҳ��B�2�<��D�0��w�6�ZYG��ۺ�,:�]nґb§ϋ+�%�r���i�Ϲ'{˷�����	��i-ʹ��4G�>��1�lsr�� 0n(�2j%�Ra��� �C��(��m��W�s���(nӏS�6�|�,ڞӝ�ɲЕ�_�;���0(j)8j�Jn��[�
&�M�[5��$�V��c�,��(4�g��-�LM:�'�K>>����9r��Q� f�
��=��������8�9����[N�Gx���*#�1Z�`A��?�KW��1�^���\T�t�D���Jp�ID��pn�A��\����E�z���y������1�E_�� j��&��z<=���c�*$
H鮼�Ez�S��dX���͙�� 9m�&�-N]@[��'p`j��Wc��Iu���/�#r�T*�z(0�Y�&t���ܿɡ��^5�����N��S�w�:�&��?�`@�`T4j9�ݵ��?B� ��(1y���e6��ʐ��K`�'�b:��6|g��i�X$��0{:q����8���_�έ����'�ж�x#���+������o����F��6�>|I ��#X��18� ۙnG�}\5@�:%*J�>}Ch��;jF�$<�-.8��:D�̍�I�p.����$f������#S�"�d�H�ڞ��e]�f{�8�V.f0ڸ�G�v�W�#7k��x/g�����HM�+ڃe/q�K��<2P:A�yrq���-AG���vrЁ �:Z1"�Gͼg�v���;�>R�C=���*��b=��?��L��e8I-�}u�ֺ��P���w:��2���>)���Fb���kq��]���ˁ�<����� �R$m��.D\q�!6�_�'�v�$ؽX/ַ�<�ђ��9�e&$IU,B�N1�޾��D�-�ӼC�X`�	]���o�9�~!�:��`�/+j�[<oЛ�Xw���D�[ʭ�6�
T���?�)�+�7B���a7�[{�D2n��\Y]�=��:Vİ�`>$H��Xߟ�8����f�Ã���&���{�����QQ�,C��Mf����fq@�[C���LJ�n8��Q���m�,!���C>.���?ӴTG��Uxbo�7������x�6��Z�:S�qণ�b�jb��q�e�J^���`T$���ˏ̬<uz¶]HR���R��$ ?�	�+�5oe�׎Kݓsa�k��>2�|c&��=v=!�A�-�����gK��QE/�: [Ĵѹ,����NF��2AeQ�*��c���e,tP�O�TM��4w0@������"�n�n6j6��G+ض7�Vd 1�Ptt����f�AC�IЉ6&ma����2��i�U�c����2�c����TF���7@+���=���|��B���G�fÏd��	I�L_+Ο���
����Ld�c�7�?�����h�����7@k�Rc�DIb�W%ʤ-�S�c��Z5&��g���o���>$�M�Ғk����c1� �1]��l[���p(D�L���2x[�YR��}��z-@t�� K��<_�4ʪ�%Pָ�`����T$'��;f8�m����ˇ�����I���aJ8XE�J�-Ĭy�������ws�O���[��.H;���/��D�pon,DV'�~�~�܎cC���%���2�m4���pXa@G��
�Kp�Ř�:��Ȗ�׶�&м���>~_TmNi1��<���᥶�)EX*T�I�])9������e�-���*��`�̬f�1h����p��i5��{�P� \����z�n������U���`���*�J�]d�֝��/*���[3XOOSR$U�_�w��c�(���N�BA�%�n/����Jg`O���q�`q(�Gpu��i��ZvwsC�ꄲU�����J���9?h���v�j"ތ�.��>i��#P�������ޙ�9~ ooy�/�N{�I|������)���I��{�X�N�n��+���d(v[jg�_�Rc�j�S{o�~�G��y�-9vز����n�El���M�����M�GC3ߡ�Oo���kú�z��[^g�p+5bb"*n�b���CˢM5��Q��ّo�������Ԥ)RF�q����H`���V�-� X�N��#�4�j��#�q���Qm�X��F;�"�� \͗,�#&ƺ�U�ܡ���D�������s!�=��l%7���7�b62qv<@��Q�E�ߠ]����O�O>�>J�@ӧc�B/u�St������5igUv�9��D�q#��FT��X��H�Q��w��|-�>�CʹvL�]�l3�8���)����j���JhF�lr尛�d"+�L5�Cn6�]���,-(�&������βX�~�� �5���Ѻ�����Bc%k��鰲Xb�=��� N��f�Y@��G�=��q�C}d�C��VL7U���Ԍ�Ȃ%��mG3FO��f�^��zaX`�0zrK�H�&��}�L�Ȼ��e���̀q����Z���-���n�v]���\&Pͨ�aی��ܕ����_��I�N4$�/~tK6���d�i4��,���d�s'J|@�����O^D��Lvj��\Zɜ~���[_�Z�n!ӜA�%� ��4����(YL�%���#"�Ւ����y�V��i�`LG�!?Ê�̦&ͅ�Q��ّV�F8��R������V��5��Ϫn"����6WD�]��i�w���M�� ]�$��
�K9ڻ���7��r$�gw��_橞3��^�y������
���ڄ97����IX�� S�r)��)���`:�������̃7�,�:�����~���(����U�����R���+b*��x����D.Ly��L����is"i�#�n������O�!�`��WK�5ST+T���X�O���\�,�&�O6�vf�Wi�����\H1l���A|o&6{�����] "1U�����a�W[����w�r|N�n�K�����1�ҕY�� ��^��ЮT(j�zڃ�A�J��?�*�HLM���
j�$��Y��}h�F0�ZbHE�`3�Z��!D�-w_��<YFag�QH�|Y,����1�+�"�� �,-�5��W�)zaEO�F�wc0~�d`����[	��'&HU'�����涘�X�(t�UT4�� $���Y�r����+�|�w<	
2/�����½#�:(1�D�x4��}�	|�9F~�v���1I��+k?ݫ�k����6f��匾^�0��E��n�㱮�T/~�
A~�A ���le0�s��~���%M�&��RJ�28J@/�:Ԉ�ȼ$����v�ڹQ�Pw�U�r����{A�]��toŮ5�e�P�0�I('�Ȑ��-�oZ�K��l�އ��K⧞���ߓ��XH*W�,�����g��A����/b� 	�|�)k��Jj��V7�ջըDo�q&+�j_,��f[-	%TKH�τA�\�?Z�<Wʰ��-�]�%I�gɴ@�8���|���S��������"bz5�d�A]"����QՇ�g�P� �7R�#�w!Z��e�P�`���6"��q��;*t�:�����!�[z��X��_�N���*72ĉ��.%}Wz>�4�:�8#|7@���$���b�A^���wA�?Hf{������b'
܀�����.K���A�pJ�3O����=y��%0ᓋн���r�a:͜��lE*�*z�{�J���A�M�*��*V�w�M�i��E������q���n�iܶ��_�����˵6�4,���"o���~��azQͪb��������5��e��������N[�uC��m�uv��}t7s�N�8DĜ?P�z�"�P�t���N�;U���#���9���Q[,Y/���{0���އ��0�R3�6[X>�B~��W���qB��O��Yvy�u�	�/�[��ݧԜ��Չ1=g�?:�����m�#�dp�f������EjELka
+R�;�����ֱp�ic6�`�����{8흘-3��B�{M��v��4��%���};B�zXu��A�/��H�S�r�lǟ�X.�mtK����0R��Gy�j�M��
[mp�)�Q�p�Q���gl(���SK�XxD[Q6�(dUpe�Ǔ \���2��"d�5����0۲T���z�P`����N���t�%�r�T�Dq�b�H���9Y.O8D���,9�#s��H=�L���������^�4ur!�BEG��R��6����R��X:�2���Ҭ�R��N��⏍����pl��.R������AZ���p�\������%$UAS|��'�7N뤫(�W�HDA��z��+�
�Ȳ}��iw#T�ّ 3��/8S���<���������86�|��ؗ\l�gö�.P��l�]���t*�VNt�Rٮ4T�r�(=��=-J��q�4�[Sp�<_
��t�*�X�\�߮r�����F:{,���
r�7�����
}C'�T@��컞�A{'ю��	�+�נ�6��NF��9��N�J���o�V�VT�K���A҅x��X.>ϒ�����>�P�����QW��[���\��P:K�����rQ��z����%gfi.	dMU���X����h�4�?�f�tx�Zi�>��q��?L��촙6p�P��������*������8d|��c�9ʱC�|���c�\����b�`���tё�ۀ�|1�I.���<ϞAo��m��3=QE�"N�.����l�:!3�*�G�����s���}��˰����F\V^��W))�3��(��*�W&F�k���tZ��)!��M��1� ���$�8a]qt�?������S������#.�#;+�$8���E�[������cX|�٨����$XO,0R�/������3��Z����F��^̇���P,Bi���������%$�3H�� ��[��Ƴv�Yi|���O�l�m��+�@cM���� �����G�~a�pU|���u�>h����аbwt���í H�7�_ޜ1E�ƌ���῕�+I��y6>��V�{�I���UA�?Leؾ�z;X?���'�| �j�����&E������!όn���~:�	�x,��8�^���(�0����w��w�¹1�E���mJ b�@ u��9#v$�Lks����m��KE�7�
qp��I0b�G�(�B��<�L��-,"�X��\¦O�,^��A�J
���j��;\��\z.����{�+����3���Ż��m�Ӕ��EI�Ϩ�hXMy�6�Yo��C�5�w< $&&dU,�?.��㈬�ϯ�φ�J�4͋f�m-���!��Z��eP�9��;S�C����G,DLY�po��}q���O����z��c�T�NZ閽��ǢwLR�|Z�8���Ւ}�f���ŭA��3���Wg��= �����qߘ�� ���n'��c��h/��B���}�4WR~ǜ����'��߽��_�/���x<�ڿ���SbhA�<�c�Hu砍E���M3��>0���`6�)�ܼ\~H������X�ؗx8#	���ˑ�����ML���4�~j�|F��c�]���@��@S���a��V�<ձ�@��q,���3$��hj��z�*�u�+TG�G�U_lw�m/x��I� �i�c1�2��=�un�z���G�٭��T����[ŎJ��qw�/�$��
6 �+�n�(*�%P���W<nݰ��`���� �7ܼ���oAx�_Q����D�x"s&��f�_p���.g���{�П9�n��|g�l��B�KH�95~M���*(l�p͹ᷲ1�[�0WH͓̉TH9r�8&�r�4ep�Ksgr,2��lm��$M��tK�UI%Mȁ������E��V�G�fMM��()�oH2��f-'�2�#����%iՄ�-��V����L(�T{�xt���I�����➐��b0�J�>BYU�k�s']�����H�LBe�Y�I��A����ҏ�R��<+�YSu����1�ث�/}n��STmn�?.VH�U_g ���&�!݄�?���o���[����5�a��a-N���{u՛s��~Tޏ�%�H����!t�����~R� P`Q�J�3�"�|F�>V��/��-���_����S���3�����G��.+�m�m�����`�ẄL���$�|�5��0Ԣ���pl�!܆�k�̂X�5�1�ZU�i��V��Y^N�Y��B�_~��J<(s)L�E���nL~P����P���Ҽ��h����ܮX�BUz1�q���;r��E�Ђ�o̔��������������Zq&%��{{K���q�M
7�c�1�9��iXט�9
�9�¾�h�$;���-l�g�k���N�$)lӘ�
"��q�4W����F��0���}岉q���d�e�1.*[����\�猔�UV�P�k�6;�0�?BO��>�	(����񊠈�ZW���x����]˞�K��%�P����j*���ν���L�P����:�!o�\��Qd�}z�2�@����ˇ��%`�T,�s�q��Џ#8�,��'��]&�����6�IȲ� F�I�����  �O����� �\,�X��]8)&_��!�
�&<;��а��ҷ3���G��	�l�=��k)�����˔{s���<ʉ�n�˽��N����d������2T
�B��ߐ�ʊ�c�Θ�6iy��������[���Y��Ha������&�
�n��y􋅼��2Q��7��6�b��~w�y	G�U�}� c�T�sH��(3ց��%x�B�/p�T�
��B�7Ç�փ��ۻ�>J��L9��b�({E�k�b[\�T�L�j�I�H�/�9�􀵭�YQ�i�@��m5�eI��y�F��a'f�>r��K#ў�y�'��{���ӥ��'��h�D�*��Y����P	�}��M;�b�'w�w���<� ��ZYo����I�l��B�F������������3 ��\��y���ٶ����u���a�^dYt_5��Og��H	�Z�y;7�Ƈ�[��t|c!4mu#6,]� �S"d���J��7�j�
?�L�>���n�+.��N,�7���,*�E����xp���w=˚�����U)�W��n����f�
s�E�B�^�s~�M��Nة��)M׈��� ���y�e%�5M�n��T�f!���Ep�yk�����Ȳ ���U���C騱�n��"��R����Mj�[L��s���{?g����p�����U'qW��_�	�ҠI1G��ۃ+���"mV�|i������(��?_�l�F\��Ԃ,�?��?�KIX�����w&0�z�l���/7��9�&����ln��k~�
���0�W� ��O-���`�o���Ô{������x^�yj���s{�p�J{�O����L`p�}=Ӿ�c���/Z�X�bTL��b	�tC���O��;R�!%�8�"j�0��HE�֞(Z��%�A�r;�YpOh=q�2�Ǘ�ݍNb�>sz��Nr��-�줝kY �<މ�&�c�T��ڋ*�V�T'�\�;sN���!m�_��6�(���⩔O�X���)ݿoy���$�	�lg
��P��P��P{�[�|�S������N���r�B}rǟ�{��w[txV#��>��*�s�R��ʤ�����j�������F���VV&��zf"$jJ�r<���=�yރp1(EG�`V&1�4R�������m�hX�a�
���d�c�̸^���h���[Be9�?�4��@��j:�{U�L�!ɽ������4c:KŶ���Q�8��G��O�/�����k,��kg�ӛx��I�t�c�h�Mm}�H�Z�!����;��]i��,�*'�+%OyO�>N3?M���7Bʓ�;d�6��%���[��ّ'�f�:<>б�:i^hrc0Wi(OUh��K�\����qEy�m5�T��^��w�4]Zy	*�Y$ۼlSm"|�믫��%d7Py�.��Gk����%�nZJeaLiL�]�5�{�`��*w�]wk�=���v}���b�&�s�`�絲�S8Q�?�w�3tii3���9�}W������K�qe>A��PK�,]����]��p�$�#�b��l�%-f��N:�����H~��KT�&�����8Rs@�Tw�4�]�j|��C��w�c\���N�5aΓr��7�u2mB�ͯ2y�6�?��b���U�A�@�R����Y���b>�Y��0Sʝ=O˒�	k�?��v��{Vָ�V8B8�:�k$+� �-��>T.�R�1.���Ph���mj�K+`*"�4���&�H嶛5D�y��D\t�������!6�t(��E�B6$s�Jd��o��	���l'_�ʤN՝��!���̸ƶ�Dz��Bڸ�%�`��QNC���9��
亮�3*٠^�r��k>(Oʧ����1��=!�*E��vlf�<8"�iz�9��n��Ϝ{����Z��Y,�Q�#N4����˷h+ޮ͠E�_�����}Vd>98쉃լI#_�=���駲�1����6d+�����I���0��S�̯N�����G����Z�9*4��NFy��e��0�4�^�����]򼑺8)m�J�5���P)�.�5����xB7��)�,���!	������X��
��&���a�`MOƌ��}�i3'~X�Os���Y��%�.@��,�EX�ߗC�K��?w<��	
I���/IgK*�%$?ʉ*P�{�F�r�0��&�|(r�w��Q�"9����e4����^[?ڞ�z S܄K�cO.a���`���J+
����tA1�c���6���n-���؃�Y]�>�@���X��pq�=�� �MQ�rʘ��?5%9�I>�Kka�ǖqZ&�E{��}��MaX���?n��]̲� ��	a�d���WMĈ2;��f~���x쳃��y.�R/[7�`�!�K��c�������6�+����
�%{�"d��a�� C���_��O��S��P0b0p~I�8<-u��|��פvdA͉�:�+_��3��{T�;�C!�M��� �4@M˥��TJ�D��0
��Z�Q����s���K����Y����l�l�[�.G����b�?	O�$�>�Y��7������!�j�;�|(�ˠ�(#ܟK�>����!�d�8�O�����m},�fISJus�}��/3���8A�����l��û�������W���Z��&���d\QI�T��Is�Q�f�*5�v��9P��t�Ǚ����(X��5�`�0��gν~W�?������#����ֵJ�jt��$ə]��5��d8�g��0���.v���}�E����ٺ�SF�]wh��OM����{�׍vȔ{�\�̔n�5�jK�B���#w�ٟ�ǰ_�Nm�R�m�/=T�T"�^���+�\��Cd3y���J�1��'�^;�h��R���Z8T�U�̽3�L�
�]��0��$�.�qA�����@zإ����f�{i �d[ ��^�h��|$��IB��1X�-�<Li)g=����ɶ�BLH��֏�Ҫ+� ��{�h�bG���9��tN���?��O��;#��$��A��P��'���4k��V��{���Є�E�n���^�)��v,��]�0�lת0�A���b��TU�DS�ޔ�k��YM#�_����{K2�TyVA���Y��/@��P��J�?n5Dġ�V�^�
~��/j|�8��,��1yW��(��7�3sZ�p(j�Ba��JhL�roE�Ō���n�K ��J�C�CthR2�~iڻ�P����)��e��ޣd":�UBՔsBs�������c:˵%�~GCf�2~����L�,��姕`\5����P�e�j���}0+E�vд�MEAԌ��S�B��Q;K��t���+�A���{cV]J�$<��:ã�ԑ��vQ�{��>�����z�!�]���J�D]�����F8l�k!ҁe&���5a2�x���ހ6�'>���=D|���(�q��5Ҹ-��q�������<�gb�)�n �5p�7A�\"�:�h�?g_Ӈ"]���?+"m[�.=��ג����0��A��[sw�
�ǥP���H�>��5�tFd����h~�3)�����ܷ��2��qa
ٍ��@��S���tm��jNP>K��v��̈`6�ɫ��PV}�_=�IͿ́�1�[D��T]�dR��]LR�u��t�0���QfoJ�}����@��꧌� �QT�Ӷ��]N��d���8������촓`AW�%�'�E������L捤di��r���i�c�dh~ZP���l`Eo�`�}�ʼ\		��s�B��5��ŌBl���g��`P6�V��?4)�_�ChP9'Z�2��0e���� �$dk��8� ��`|��'X`�[b�܎��BFSw[o��dsꗕ�9��4�M!e*i���-���C/%��K��!�U7 ��*��5��k��L*`��%M��2�I���2�I�o@VB8�d#��;~�;��웈,z��?��(_���۶4$��2��.Ԏ��(��@�{�z1���7�����ט�2C�D��R���$Zk+�R�b
!�F_���8��C6��l��UCr���pQg��r�&����t3�vd�[~@�K;��܍iWA���Z�!���"�n� o	������{i�^��kZ0���F�+��7����������WY3�V~j̫w�s+��E� *a���A�9/ ��˻�Th��v[j�M� �h�oxo0�bI�w�<���JQ���}�(=��/Ѐ�E���������<�	+7�������o�fk3UK-YLFpM$R�'f�ѥ�^S�$�{Y��N��r0��[���;"���@i�?i;�*���$*^���U��\�S������\j��H��c�A#akl�L���G5�#]l�QN\H�x�aA>͹Y��$)�������_�S%]y{e��(�/=א������7Y^	�����vEvV�!��xl�n��aCtv�;8nc�Դ�3[@$ZX2����đ�s�*��A"��,�!	��7�q�.�֟2!}�}�"k�p��f
\��Qoi��CO><�)�n�
9���9Vq���Q�P���)���c0J� �@�s�2@qjA<MyDi�K��Mz%#����w��x�P�����w(�aq�*9$�� �_o=�_�D�?J�U!��N*�iR0"3,v8��6����K��P��w���&솕�q�?��m���"I,V	��Țk��e;AD\ԭ G�n�O�VQ%p�afv烘�)f���i�Vl��G�$�$�8ʣ��W(��a�ué�"�/���~�FH����C��M���s���9 !Vt@�U�\��|TsG���bU�Tg�+�eN�j{�k)O����c�?��SB�gQ�1��K�|0�k�l��|��Z����G��H5�8ɪ��v���Yߊd���E��7�R=�3P�ĉ�}��R+A�*�M����W��YLw�g�/%��>O8vN?FC'�T�5�'����rc�-N�BO�a:�[�{�
��N�*NŸ�����r���ш/���P��c�JRփO�U`���j`3*}H	�������-=Lϐ9�p�N�
ϰ��8
�0�5:C�@��c�יּ$��
���nH����*~,a���ʓ��噂]{ԛ_ű!�Ƒ�r�@��/_J$�7��VO�`�c��l����}���a��hP���	�^�`�[�m�7�bu]#�+���F�wT}��_$�eFe��@�딫���(p�ͨ<U���Ts$�����k��. ��?[���;������ 9LCŬ��hr@��Y��..�:�Z�̷�&��l�{�HH�v���@�,e$E�_�nO����pqRU,�����̬���C6���PkEu+Ե)l��#A]���Z��&�������T"$��
7\�YrMN6��)|�sF�/GaD�-�,"�d�+���|MUb<�k�����������W�+�����4�5��%9U�6j1�����z�j��8Hw`;��)�"���[��곂/�]'�s<̌�֍�*C�*O��W��\�~�S�M����z(p�F�-Š���RQj"�!k>��9��եJ4�(��~N(�S}NgČE��LŢ����o�a��0�h!�Z�f�xd%a�K���ͽ��*�9~�9G�6�t��FSdBmF�}�(�z�����p�pq�0�j���ލ���Ň�ܩL�ށ5(c�x�;s����M�̿Gg%rA ��R����j�=�,�*r��r%b|d�����g�)AQ�����4�C�9z���"hc:�X9����3�q����,�����m�V�h��H0[jw@Y��3������i��v�A�T�9q|�s��o���W9��(m����c���Ǉ@��'�s@~u�����(��>�߳p;�Wc����:�z��L�I4�Ly*`�R;�|t�bGk�/�F^��s�l��B�g���\��#8c{ѯ;@�I��������aMg�p@�@`��V�S2���·��ZE8>I�����T���,`�1���6�{�e������E/IB����Q����H ��t;�՝��7N��'Jh�"�y��yN}�D���Uw�S��H+�0�AP��oR�u=;�,�1�G ���<������mWUp�[i4�#55��~W~V�����7~֔`������#���g�)���C���T��������+�O�A�^QN $y�*j<K�S^�u�.�[��ٳ�!�ݑ̫_��=S���\��.afH��u.���1Ӱ�Y�3#,�:֥�����:�B���c����"pl�rs�����snI�C�e0�㎹ǳ���x��\����Cy�J�$o�ſ�R�
�.����{�ٶj*�c=ܑ��{^ �W4(�V�X�J����K��=n9{v��S* �^�A�&F)�0p��O^^\qD�粷���;��H���|C6C��/�_?���z�z
F�B�����X�)<�T�xή:�!�]m#��a��}��{��]�z���r��q���V��у�������4G��A�/�D�=H>�Q�4�k�����)[�{	w}��)j�`��+��rJrcn0�Δ�l��{��p���c,~V�l8O�&�_�؅���({�Z�j:TVً������ל�����v�/�S��v�V�3A�s��������l�\�ۺ����9y`�y�+���)�˚�4)ܯ����@U3��J*a�����Τk�9�(��B'�D��u���3o��?��6�V�9�L��'xۤf�_ T�+�B�h�L�>����#�UK��g(�{X���\9;s;��s1Kn�ّkᒍ͂&&��g+OG��d�Do�_�����#�k�cz�f��dއ�xN����]T8h��C�o�|�hy!:@S+� ���6b�^	Z/�s�i04�a������=L[5K&̖��{]��a�eqk-�~�/�1��l��{�����lrP2 ��ݠ�4���R#K~�$��.��ᒸ���t���8�T䨫ٯ�!GS��"?ԍ"�j�4�.��E������ֵp����S_��)�N�_.�85���W����h(��&+�#���;�[�s�WZ������\9l�@�ݐ����t�Q�J<��J,�^�EX7�뛟�[ ��DY8S�����v	=j��ad(N� 8;z��g��gUwk�%���Q4�L̄�l*V3����F 2k�ꖓ�Ͼnf�ٕ��)1��G�P�X�lZO���tSY��I����N���LY��/]���Q�p����O���1-.x��Y�衵A-1�M	��-��|]'@Ѡ�L��P(_��?�a]�:��Ӳ�9�"���VL�yЁ>����O�������b�(/c?�s�@P!?#C���g�/�gBYʻW�j�^��b`�R��+QJ�[��3#=z�q�Wx�_�uAo�9+�B|4��"���?>�I�q�":>�Y���Ŋ<@B���� C����x��|����ɾ.�͆)j8�7`K%�m�7�3,w�LI�Ñb	�U���Wj�ځΤz���O�����/�Oa���]��%�Z(��@�w���<����
f:��ܹ��?tC�X��M�� nF�q�0K���0Z��Gys�b��b��czU���J�����9��1���UL��k��& �2��+>�PFSyo��ԧ��������Ճ&B`<j��#s�@8��d��l�n�o{�W���;���zW.�����Zm�H���N�,���V����Q�dYA�C��KՉ�yG�gh~���V4����J��)�莁������M�xԙ�K^�P��կ7���Oun��]�7�˟��X����H�`�R��ppX5A@'��53@%Q���C��
�AG�����Oyɯ����Ȫ󥬥E�0 +;�;��$:A��G�F�h�R!+�qR"���B{y�Z�����H�T�'7��ܑ(߳4|m�ķ{A7�zF���g��U����m�Z-�QF`���v3�D+�\}�(�����i\�y�tPx8X�E9�"�����Qwr����U��<D�##�.c�=S�@��b��I܎���v�)�n��v�X��bE�.��}�����dȬ����eB��:�w�y��T����X9{BȄ`���x�`�.[��3dh����H%��������0d���x΢��
S���b�[�T���t��(�F��N4����N4���w�OM<���k=�7��*�8!�g2��B�G2�;��d��
,��ӫ���|l�!�\w��6�����s��yȅ������GK�ţ�'�=Yi ױ��Ʉ������o�_��^�IZE_�*��n�߈6F	�=S���G�#�1C��k� EH���[����c+� �H�:�B�8o�2���{�v�d����`��9o�@�-�R�j��ڃU�16�L(��E�S5|�{�<�~�9ڜ�5�y�,ܞI%�7�b��������5c\����#�4�M�M��#��8���#�@�QMt�^��Y�YZ���a�=��"���ΐj��ȳ�N�*&u��è�|�?�TQـ/�,}��Ŋ��Dm�}[AJ�^�|��D2	���[��w��T�B�~h�0� �_���+H���ѱ��:�KD	����1|�X͇�����t�G]D5�!�L�wj�_�W,�Ѭ� ��j|60�;�Q� :���Lr�Q��i�E�VB�O<����������u�U������#�#��֨Z(��#5տ�C5���������%�~��6#b|z�S�0,z��=��#��ve/5K�����R�Bn(?v�q�7�g_�&��4���tdѥ��$��F���v�� �x��� ?K\����;��n�xV��i1�tm���
��a0��?�P�,W�������M4��
z�w��m����>�hq��g?I���ߩ���>�R`�|^o��=���݊]�L�q���� 2&؊K{���Ko�����V1@�SF�Z<��Љ�3�0�}�~dzz ��H�p����'w��1��Q��s��D柔�ؽ�`~M\��m�,Xce[����{L.��_{I��p�T�̢u�a��$n!w�dIc��ɔ����[u��&�W�~��t#�a,k�G|J���L�� [S%�d6	)ؠ?}�1��/���B,���D$P�y�K���GF�,e;��|�"FX~d������&V��BI��?o	y���_�0��$d�;�OAF��.�H��6�E���#�^2/N����)M�{���]�E I��<��HX��d�o��$�5Ƌ�[4{�~�#*����MS�=�1�5�ޯ��d��)Ovh;;�B�۱��j7>@W�N*�~��H���,xt�r�0��y��o5����-]<�~Y+�6��U����O 
��G�$u.ɘP�k�8c�� %0�&ϒ0��(��w����*ю&��.'���r�k�&6�e��n!g�-n[&5�UZ���<D�1Y��_�/K�=�~�ӹ1���>�d�n��d��vH�^r,�n�)7�$��'�!	i[g�F�ǯ�|�H��~{Ն�H�nqEJ���@[t1�*�,�86Wc;��w%P�9�{F7��|-R�-�Y�w٤� @����E���(�'7R�=��1q��Pȑ'e.�%�ݶ�{
p���)��} �h��!�2v��u�<X}&|��S������O�@�k��2PH�*]�`מ����a�uvDH&J�~����L�/VX���"�e8�;�E��'��>M��݋l(�mY�W��B�A��T�d�/�O�L�kE��;��:K��['��*�1��"Y�'�M|���A��[�bdG�y#�.�F]�uyٱ��$��qj0��Ј ,go�"��]!3}���hPv2�WXK	�y�����=�J�&��s�I��2��A^E'הڹ�f`��y����_�VA��:�bѽ��A�qM5�L��߳�W6��T�ݝYTI��WB����L�bR8\a��.b'	 ���h��a�Uc,Q'�\\ק����灝z�6�,���#��4Th+��oS������~/��ąD�^͍����U�]�3m�8��1����#7fC-��x�N,�Ӱ--��{����l5�>|;�'����yV}�RǺ�� 0����O4q ��x��i��,���Iݡ�"����p#L5����l*���y�$�ˠ(��w/�cB��8˄��D�%q�ġD���C���?j� {�A��qp.a��{[֐����{CZ��N�.%0�
���/�9HlqP��3����cD>k�>�a�BKP����?<|k���	��26UV=6�����C�gɻ'�^�^c#�i�Jt��T�K3�r=��:�,�iz�T�.^~���4�*v>o��i�����^��9�!�Zfgb�Jz�Q�X�LUl�ҳ;�?�/�q'�e�0d��|��j�zɺj�X�u��ʈ�U��D��KEi;������x 9�J�mτ��'� 
p0������cZt��X���!:�Q��3C�ق[�$�M�[�gx��0��na/�;,��"�����_O����a	l��S�]��_�\-��X�u�.���Ĩ0g�j����I������--%z�۱���S!�y<���g�lf1�2i?�Y��Q�NP����v��"�`�	!��ޜ�wƝ}q�����=#��g?ԕ����?Go�� ��${�@*~|{���L�Cj[e��;�|�;�wZks��en��咒�2;��M�p�#ܘ.�u�~�]f���Z�Vs%8�+>��w�2��ZJ�֬aCN��R+��j�Zdy�\����=���q)�]� tU��׈S`=��Y�[��j�t�g����RE�C}fDm{<��+Jb���$�}i��E��Y/��  x/�4XB����+�}���������:ى�̿,�� �3q���:�pr:ࢯh��Q�g��G�DT��P��z�)��ݪL�C���c��L�L�R+��)��j�����������r�)z�%Ͳm,]p�`�&)�פ��?��d	��e��b�ԇp2��`"�j��~W+Ӗ�5R��&#�6�8F���.Ĝ9��Jhŏz��֊�����t�8��'�w�9q^��C��B�;3l�=�K��L���s䖥�\a/6�D��Mg�<u����_Eq� N&����?ԏ�q�QÜ��L����'�SJ�h�KS3��p���AÌb��޾�N[xP��+�6[GI�N��vK�8*b�+��c�_b 4=��́��a	��{!4�H/�e�q0� ·_ڥ�{ސj�5>�3�W�y�'������C)���["��ya�C{zd��?u٢�q�_nr�����
���ɓz:i��׾oQ�{�e�.�i^ �	w���־5�|@����"˩��6:2j= �Ym�5g{V���"�����0���;���:׋�B����#���S�E���ٿ���m�Ӻ���;�*��z��n��2L_Z���|���>�j\<^��$���|�"���G�*	�KY0��\��&�{F�/�p5��<Y��B}6=��?Hi��.�d9)i�Ir�� �Ƙ�eXG�a(�&&,�n^&z��mK@Y\c�gF 0�R�ʽ�^/g�X��Js�ݥ(-ت��e�	�m�<3|�.Q��xI�HPjs�cGuHԢ�d��o�|���T�à���n�QqT: �)�q)ԧ�ӊ����L� �\q|�x+ڑ�u�{PON��TKlyv�j���{�.�p��w?=F�`�Sgf-wSG��P�^WrV�<�O��@P��E� ]�Wh��g=�5J��2�k�#�5m`~zD�403�)1Q��㲆ۜ&č��/ϻ��lpY��'�gLb��u��OyOw��N'�Zӂ9 /@�1��/�{w��)~�rg%7aB{��^�<6���V���
��}��L�Бc4�SAf{��A�Ӯ�?}�yPƂ!ַ���
g5�r??�п���FQ0��\"�&��I�!T7��c�=]�2JE�D�J�g=?-S��c7����E�/���<�����q>yX�Gɡin�p��-�5�y.[��V&�K]��X��a�ڂFP9��kAR�Y�׏�Y0+������n����F���X�yC�ܰ
9|̌������_L1q�����]l�D�<ʠ�(�\=3�M�y��5��ru�r�'�O S\_A`<0*�HyM��ۀ'#��h! �o����^�A�g�`���x�n�,�Rum,����p�i��6Z
AS��@�}���q\�$=�:���TlD�)3�o%���Z��!|�{�0=���Q����9d��^�����mm�	�RU��\!��8��Q��b�����r����,���!�ّx03��V�X���2�Ň��$h}�I���s���TSQ�x�D�@V�nM�z��JcF�p �b���e�#ZO�դ{w�#�v���@˼BJAj�z+2ءu/2��0����]��� �-_3�i��qL��J�`�v��PM%�=���h�˶HJ�A�,-c�3�j9������%��7b<��"]\�_�����*+1��|�q*�cm�^��v��R����w�6|V��۠2�ͥ6}{�h�+��~�)���i�p��q��
��/a�O�^��`���i��g֨t���v�3� ���2W�[h��a���Yo�홴�:j�9�@rb�q���sΆ������@��@�p���A�K3��^�H8��qo�ss�Utt�]����?;�A:�����6�����*`fk�ϒ,W�Ō�b;�)}]�w�Pha��o:�4Y"������'�B|k�iQ!�*�Z�P��C)��:�j�N"�v��o��v����@͢��&6۽wXQE~3�!�����kc����ўY��j]�l{�ihU��E�H:Қ���G�߿�I�k��v��T�����-���nT�x��e�iW���+�6}���@ń���d�V+��<*�[I�����,�sY\s���Gu1 WRka�B���e�����4���%�]S��곐�Ø��Z�R�x�9�'��5��1����8^�{*K:��3��~�ruu�;���N��40��b45�nUͮ����)���iylĶ;��=������{�i�+�������h˗^���'�V7N)�4����X_jw���d��l�����cvJ����m&��|�-���K~�p�{oo���>��+�p.s��`���>"����IbO,Ó��mgr�����!��������f3r��ӫ�`�StO?g��:�
�.��
���Ag3t�X�1����6#���.�1�2��|�}@�z��Ц��2	B��o=�'�W��n׀%��x*WM����~b^<l�M�z�<�+��ߣټrÇzʅ�l#qH�æC�%zg�g�V�iM��"�V(��������L\�����Ż;�T���[���@�>-'��掇�ŭ[��H�,�'�P����9]qvc��Y�z�� ������(W:g�P�dSWO�e�ޥ�J����ؿ}F.���7�
�Ьפ[�,�"�Bt�	��`1qo���V��׶����,u�ߍ��Rӫ�~���0Y2�-�g׀KBɭ��S͗�X"0�\ ���z۷6~�b	,��G�R�_��5���w����I<=�hQ��K�Y�#��`���[�.C��x�J�mE��܆B��`��o6��V��Z:��W|�JHG�0?��H;�3iUrr�Ҽ2h����y�/��=���z�O!^�hT*�*0ˎ\�_T�i��f�
�Rb�VR�bV�A^� �\����đt_�s����*@	�aL���'1c�'cL��,��FW��э�Ȏ�mwI����=�rF�8ơ�ZE(�(tT/�B�yQ��4��ݞ��I�3�tQ�.�4��yf�1?�g�uҴ��}��r�Hepn $��j��>G��e�#��ʀq�u;��*�7����"`���;sU�������;l���&�&��bÛٔ %�?�V%�Z�+�(��eu[5�ʨɇ���������h����kW�9yb��d�n��ЍŴ"��)�I!�T���9<}/3� �2G��c�� 8�Z{����j�G�gk�<hV&�~%���P�ͅ޺��pe��A��U�A)aZǪnn�Nj? ��{�S9@�h�	��_tB�w��D	��,V���&yņp�ey&������",�`[�q���p��u5=N���u�7�%�W���31�����yjv���.��F�H�M8�O�W�*h0H�(�ʕn��oU�1톅����D	of��H���0�o_J��b�D���:T9����T�L��YVJ�,h�����6 �땮;�6��4 ��)Z���6�>��q���X��K�	�Ed0�?"��Ġ�0��F���Ɔ&˨����r�o���Sd�1��X�Wl8[�ڽ1TC<�	KA��ep��"І�N���� x�?;�����r'������M�Zʌ��2�a+.���\�!��p@(�N]wb���W8vP�kc��~�܈Bh���I`��Q����>$��T�ɭ���2F�a<n����j�'x0&,E柨.���m��%[=��q��3�<G-��eᮀ,���y0�6;�A	Q݃ݴB�4��b����x�39���V�|xÚ�o�P�O��5�:M[��C�[f�OO#�������D��^�[�) R�f��F?���n�p�u0��}B��B�7mr<�/�&�����!��'�>����ڥ���:<6�.f�����oZ��CJ⺎�'yZ���b�vPP���Z�@�-�yV���e�̮���u�p���$�e�/��!6x�%�*��<�+�Kc���Z]vp�赮��<h�UZi�8J~f���ћ��: E��8��߇+������_�9(�N2Uc���}�J$�l�P��)��0L�73�
�,�܀B;~㺰%�+V^45>�yK�|����p�e3�Z�G�̸8�~�h�X�9���@t�g	�Q � B��G�		�W����\��d�OS�v
 �'5�3	'��0���ɷ	����/�9��|t��͞��tR�Rx�e��+��Y`�	ߕ��I	L�Vq�/���#��寥>���P�`/W;�;%m����fZ�☍�d>���e\�Pc�m����u�W�8ĩ��ݪ��"ì2�;��>p�YN�s3S�D�A���#7����D� :�(o����<�B���~:um�2��C8,9�[v�(�}�{G�f�o/t4gzg�K:X}΢7��
k�>#2&�@�t�|8%��F�����j� �E.̌�R�(M^N�p!�>��f�ǰjt�����zm
���b5��@&U זM�� ��nI�ʮn�z�C�CT?ÜNGy�y���Y%�\pf)�R	K�M�rCh'i�3oż�&E��tj8�͘��hU(�8F�g�D4dn$_v���B��7�����y�h���ٯ:�� s��l��!�'�Pg���7�f���ĢF�|����hJ�b�捿��S[��PjL峜�C+Ci�ȉ�h�ލ+��j�-8%	t�:n���C)��,?P�lb����0+ܚSOkca��
w��B����:�hC���7ÚN;^�ofx-Q� ��4>g��R��[_���S$�uu�Ix�.s�v�x>MX�G�Q�����9mK������>�W5��Q�޽H3�JV�cCD�A,|��=:�Yٯ-u����2	9�h�"܇��5P+�v�Л�h�l�-t����ѦiH����U�գ��_$"/�>�'�z/:�2@�g��;ET'x�M����lr�$D�l���G��-Qo�l����W���x���r���-kyP�IY]���m�=�ͧ+�B���3V+ ����͞R#���$?DUa����:��fwV6���3B�FV��Ѭ�ȫ������l�O�-�Lov��~� '�DH[����M�����Kop��SL���H=x�k\p�7<F+̄\=�V�/$l�����y��8ˉ���(B���7*ݒV���W1 h�.p�>��xe[�~��$���xjo����f6qK$�p�:��cZ xjKz>�l@�&�@Ջ�4�5Wʐʭd �א}r���Q��q��/��5��8ؔI���z���a����),ܘ�&�D�>C����>J�!�.���z�?T��Hkx�#�u}�����z���	3�?ly��RHVs��$m��_[7�39�.l`�� ���c��D������R�f8춪$�&�B���}��!h�K��̚�'���_^vf�bMN��U/��ִ��v��ݹf%~��6$Ʒ��vL F��|pʸ�+��,Qtw#|me���2.�́7P���{W�hU�6[j�>s�7���Y:ˎ`-�X���"j��ڕ=��?;xn�;5�+��l����c|����Ð�*&[
�y�|���]"�b�&�e����U&_VQ�5���-�E�X,6#��}kV>t�8=��Do{�Gs�Q�Җ��ܾ!WA8���%�}12��/�����X�*�r�/"U���U���M���C	9`�ҕ�\�P	��z��Z�Nu�W�C�[d	:�����j���|*
�ៜ!���*(�J�3t҉�؜��Q������ą���Z��������Ӯ��gb s�6�$�e��C�x]����D	����� 0$�*��)��#����4�%K��&���_sR��-Z����ڴ���1Sl*� ��w�7�z^��c��#���v�uf�<de��9� u�Fس7_ͣ$���I������I;��.�����[�x�Z�
q2rO3`rR�C/:�r҅c��3E>�'I����D�"����z��k�����܂��mYjwd���;Л��z������!��d���Y���t��{1��u�ǖ:��!Q�D�xX ��lW�j�͜g
Z+RW.C�rh���ES�߮�@��=�zߌ����Aqi>�&W$q��I�+��Kg<+��1@v�ƷEE;q���Q��	�����Z�U4� �n6���]D'ǩ�I�������`&5t?EŅ-���HVXU�G7ǲ��{5(Š�����_|���6��>��%�d��p
xn���	a��b�l�G�4H�����/�����ϭ��89|}�C,��K�ݤ?bH�j���B�M��``ƚ����,0qsþY��8�L�1.��_���<���7)+!�3�W�q�,�X�3G���T���0�₲��0텗�Q���c/}9�"�c8ۃ?3��V�ӑP+��}t�_��ouO�Sn������HN��{̮�ޥ�	P�UY�O���}��#+	�w�Ci�>��@����1d�ʨ���%��L#��g���=@���ڇi��
����y��$�R�,�eݲ3���+P 3Ǚ���$��дi}F7��&��F<N�<$��ا����˂i$@V_�~,�< ��H\p�q6�Y�pZj;�r��)��aJ�����R^ɻ������
V�#��;�r ϶�zB�TZ�-�r	�6� >GS��V��2R)ꗗ| �<����ƣ���d	��|��������+%##��5-Fj�)G��jC�`��n��Wg���K���
��� $s�� �&sw��Fh�gO��͑ց^C����J|Ь4DIWݤ�E�)�_/��4�-E\6�.�Siv���2-ߌ��u��$��
��K��a���4�Q�I�ߘ�e�U����1T�	�L��8�;���Q*�w@��Z�q.��D%  	�35��}˺�fZ����	�4"z�sv�k�ͪ:c���3�L� �&�<v.������)�gM��*����#��C��������Ж�R9���K4N������?cY�mP�4�6�9W�E_�gd����$�ݒ%јS0�>�%9�]lSxT�۰���ކl
7�~�x_��a�굕�! �~�d�+���5.��FM0ˡY��~5i|���F����6��CJU݀f��C=5X����#������ʵѱ}��^V�+qRl���C��jҟ�����7D] �7�3�/�"n��H��驛K��y���0�� >!D�>sп2 �ԭ���O��4~����E:�DK�)��I��bH����,e����T���lG<�I�����E�2�����z�}!��S�=����L^Vr+2QU@���k��\���^�q��J����A��@A�7֨G}�13�m��4������-y���?T3��X3�dZn�p��B���]��P}l�kV:�D�# Gu���R���?"�b��w�u�n�X��G���s�p�v����Q,�� c�k���.,�*��A��p ��ZbB���r�r����K�c���h���)oegj\�*�)��}l�O ~�Ǚ�f�Q�������e���s�mx����0�ab�S`&����d��h���x'��"=�R�7R����� ���u���g�pc�=�B����/2>%r+;�����$�msB�js@��$�/N,j�S^�[�	���d��/�ih��Dnj�q�~���B���q����I��@���=��w�j4���"M�)��|LQ:J�J���T*SPSx�D�d�@ilS�G�#�n�1�3�:��V�٢�?��#�F��� vD�qxJ4��N�ި��X:;uf�3��ӌ)�~"���ԝNy�_��[�.a����ڰ]�A��1��}��}"ǎ�&����j�O�Ԍ��'�fsɊ�W��nOV8 �~�9 [����K��íbo)k���������&Ѳ�kO����o~��q�q�y���f�C{=��7�(d��d�%�Ah-����;����u~�L+r�l?�6�|�[�W#�z�駨j ʀcMe��R�5G z	�����V���Ľ�&�^��Y���;������-(���E�<-�����N/b����<�Iǳ�ڟ28�,�BƀQ�d@-w7��)��<l��ZS��_m�Iw��Jh�膶 b�n�>����S^_O3���6
YW FO���_R��s�M�6ml�lL�}@8�A�M�so�6M�����'�|�)��w��<�^�k�pqgm�I���/��X�H3�B������"�����	�S��߽ޮߍO�!�M�H���O
�<�W��|�r�Z�s���4#y��i��	u��q����+Y�'2:2<��4b�izD�h���Hy�v�b)D�=r8���b��"�	�����#��*͈�56�Jr6#���4[FK?�V�Л��3���q<���/�w���}��e]^U�?q����#Ӏ�Y%49̴�m7�nS'*�.��k��B������g$��J��t�r�_��G�;�G���(����%�Ϯ���b4=`v��@"Vܑ���K{�ha�����N�t�X��iIu#(��G��W�/�k�
<��8�l�˗@�Qke3�+Q#�	��S;Q^����D�*p��>� /P��ۈV���_s%���9[�P�eo$��t�۔�}?b�w�q�rD�B_Ú�n&����Nƙi�厩�+��=�=�]_gW�y
��5�w��e��ۣ��������F�`����3�o��]Us�2~���B�o�f��%�P#w)k��֬��{�E�vP�쯯�3�Ι
7�ǘ������7�����B@7	X�����&��I��{He��A��J�մ�v�r��(9WAY3�f��-m�E¤ځ�X�������n���r[$���H������2�:�B���?�9�d�}�~_a�\��q�Ә�ક�#qt�h�J�[���t���Ě+�4N��*�������#.��VԔk-V�,r�����Vh<�ճ��2ĭ��^��������U8��.͵�6z�]#Xz���RΆ�\�aǍ�Ě��ܚ�Q䡃�Kd�}��A��y��,��@a����Q�����n;�RJ����M�'�/*��a�خ
�#1���}ɪi)e_"2���Iy;y%��������A�{i
�wN[5W��A 셳W�2�_��=������A���޸|[[/s�t䁥U&t���8�l*�SzR�(���ۏ���xQ�ڿ8͗Wy���8%�Y�"��打�k�X���^1#yB|� ���H���*�r�EJ5��;~���3n
b>���=#3LK���/a��?u��_�7s|ɫ��f�	���!�8�m޴?�	&B���a�������\la��y��AWy�6Az͒:l14i�q*�;��X��� }IKD�S,l��$Nt�x�S�l�٘o��F�����\|d����������Q_T�� MD�����[���&-�o���	�6msZ�\TsSn�y�2���8G�&7�0+�����!��r6�wF�	B(m�+�-{J���s�����8jI<����a�e.�o|V��S��I=x#�� N����� �vy�o�_+!�l9��;G�-��	H0�.��^\d� N�����!�����N^8>:���� ��O�<��R�O8V�YL�2 �#�����ЦS9SM��,��$_��\/��X_p1E�'�3x�|O7����C/�O�$��:3*��B�D�J��#3%����<����9_G��x�t~�9kb��F,+�����V��(�]�#�hW	`�F�&�[�� 1z�|���?U���v��r8�B�jD4�w��j<�Opެ�`�I�v����M���v��$�4��2o������}�Б�;"�`x \��ل�r�A��3��.}����PS�G�d��jE7N�V�;ߢ�/\-�c�0!��T�/��eb�F��r�2�Y�|������ks��8�=T�L��&���t��^�n�Q}(Jh�� w���U�Ϸ��vs~��������P�O̚4�:�}"X� �����C�a�:	�3^�	���k�N���b�m��QYM��w�)�0�������0b&��Le"$��I>|�Q�f�`���dpÊ	qb���%F��l��?�Wk �R&�w�,�~�_�ݱ
�ޅ:��O��!��|��ԑ����+��W�T�5���Y���2��k��6%8G�S�[?���K���[֭n����ݾ��ї�����*/2T�l>ufOJu蘏�;����7a�Y�ݮ� q<՟�f�Q)׏��	={�����U[�T��S5��%Uխ|�qgx�D2���gSlo�v��ƺ�^oD2��˩�����{��Xv���B�E�u6`Q6p����*����_ۮ�HmU�-d2oQÌaf����
���.]o!��|JK$��vF��;{��i�q%����y��<s�����I��
m����sky��!�8�|`����(cB�Ŷ�-�)}�*������>K��Z���]�3�+9��4X�2��� ��
�������t_M(&[>\�0��{������G���n,O�g!�NG���3Wu7tky�>�'�i@���%�)��p�GӤ����M�I�q��*�ϑm����/f#��h�?�+�PJ묤 ��+ɻ�����=:.���?O[&7a�R���,�ÛV��ıv����C2��q�K����sd���;�jD�U�ޕ�0"�_O���D����+�=��ͯV���h5I��yh3͒[���;���. ���V��Q)+�Ѩ��������X7Q���\�Fe�ML�F��!�TſIʜ�w���PH��}* ��B���U�.���W�0�,�0�k;ѿ�F�g�.��.f�6�c���ر��$Is�)�����
���M=�H�Yj2��i�6��z�4)��H5��0��.KZ��`�	��+W�^˒'�� �M'A/�Ѵҝd����2r���.�I�8H�SME��4O[T0�D����h7�W��.8tFU8k���(�����9ީ%ol�����/o�h5���p����6�|=�d��D�JN�����jrm�:n���z��q�I䊂� ��kpa�ޒ��Ґo�kTа��$<S$}�I���)��C_d���1F������NU,㺗}������Ԧ:�n=0�~�L�� ʡ�@�P����'�_����V��I�>e;x�Xl��JN�q�dW��։�Q��s������ &
-|�d�^���:-E���>e�
A�1�ef�nR��У�Ā��^��C'^��=�ֹ�Ak-��ӕ��ޛ�m{��f�qG�[|��(�Z�ї����b"y�v��F�.V���@^t�Ĕ����r?H	~�A�w��s��Θk�j\�4^�oL������<0����޼.jV��p�v=A�/G�㝪��nb�m����𐗬��D��8���a]>���>�|�����+V����aI�ȏ�+��ڕ���Qmz;��k�)+X���	�~�18�f"��:�����M1{��\�L���0Czꌀ��Hw�y��N����v��;������1I����b���GX�_�g�`��i�t�j��V]��C��ԏ e��({n2՟1(���B8����x�qL�n�O�*쮀�O���N�y�}x	�ʌ��E.�VA�|Z�����8E��)�B>����A���Ŭ:q`��a�S�`�^�����mt`��v���ƚR�+�����l��:�\�̪��
r��Qy.Ƨ�?����p"����@�D�VA���kt`�����[�ˠ ��jp��#���O�/�1���B/�~֧�_m:L���O@�����,PNu�V3Bʩ_Jk�.^5D��hwi�L�)�Q��=?Sv���,��n��/=3���ܮ/�|l,Ԙ���(�COW�e1���0�CX����!)(��۹C��-TqtY�!�m�\F�u�\���f�`���l΃N:ψ�)iH�p�6��,�d��S��Fn$4b3�&z���u���[�v���!��؆p��TN�8�sFW�|R�b���Hl]X޴i���	����VSݹ����Xا� ��j�qaI9����Z�
9�gȠ���S���y�h�,=�R���7�QQ�C�j?�RK� ��[] �K��RS�\iz��C��H���-Hz�F8��D��]`�L���n�?�-�ܾ�Y��x�+�k�v���N�Yŗ�(�"�1�k;Ƿ�@�{���z͂?OÿxQ��}^�%cﶣ���?{�Haf��c��v�XB
�ƋOC���4�Kw�;�����ˍm?S���#~��d��葒�|ϋZ�0@ie '̀�?	�=I�h���ي����IF�A�ϊ*�6�����i�d�b@���THZ��C����O�S��c*�~]*9:�h�-N�Q,�L�j%1 �3jN�h�&L7��| x՘�f@yD[��*߫v|q���q��	@�L�s�(��X���G?&�ꖰ���i�-�V�}��7�_1�CaV[aՁ�0̋�7 �"K��e<+�� ,�M�`2��~��m��$3��V�������c��Y��ݥ�B�mA_Ey����U��C�!�@Tt�`���ϼ�J4ñ��A�˃������?��9g��+���z(I$ec�O�Ѽ�]X�� ͪ� �D��K�.���wS��u	t��C-e�$�M��p߳����l����+>��樥��aG	"��؟�����2�A�oX�	��D>�>Xf_����T �j��#n;ċ��e��G6۷�w����e�	�3��g$�	F�6�jL�' �|Wl(yڑa�S���zcT�P\���k�y�aw�H&�����H��J�s�_�,�鄎�"~�v�d�K{���3�+m�,��9�Mr�
rs�X�L��<I�+�D��LU�y�)٢*���y�V��[]����9@Am2~�%��Az���l��P�>W"�ZYs���cƽ6�~�^5%d�*�KƆS^JV�C�~�Y@�<Лܑ���׍Q8��oUC�<��_��;�xit���r�`;�Q�W�vğz
׮:P�j��Uե1��-:�2�����Sݫ��qK�� �4`.�s��l���ķ^D��������/�!F��lLc��Q�o-H�r��8���	yt��ﰩ�o �ITLz}�E��S�1ɒ:�I�E�(Oƶ�� ������9C�j���&�8��%��gO��".��w���jP�{�$��_vZ�9\�@�9-��jF���8u�x��m�g��7!�%G������2nŉ:e%Z#��q����N�!OL,{?j�����VI�:�!���4ϛ@7�{L|��%F_Ev5�6ʐ��YtE��S{d����lr��H�)��2���1b�<�	��g#�N�J,`�c��	/��׮�Qc}��w<��'W���jh�-�̸��1������>+�}���j�N|?k`�:dT�$4'e��2�u\��<6�k�2�v/N�ΰ\�1���
"G��ǭ7S�!
�F+kJ1}Ė�|�5�#�x�4�+�ʭ7��1|A��/��B-nrV.�G����
�	4�\ķt�]R��/���o��>�z��P�)B���؛��_�*Mǭ��w���S�6�Pq ��8��ע���>��* ��o���l�Z���j��5ۑ(v+�L���Y	AǪm�!�t�DWYt�Ozwi�(P.'�YN�2t�hR�⊵L_�Ɔx�+dʕs��di���aЄCgPD�t�0���_'��.l�#�y��G���U��>�\H
�G�:����m5F����4����q������V�� �R����>!�c^f�B6צ�3���	�r{�X�2ɞX�ąEP�G�{Us��6n�ϖ��E��E�
�%�X�������^�;)ŸQjg�������H�("+t��;��-���4%�&H�s���&j���!�$�G�큽E��B�$'>R����n�U�A��ĩ����n Ɗ�Y�Y��K��j�N�����3_�#����o#�������w;M�c	e�V�&��*��Pw��9O���	�=j��I��Tt�{�u�����J�|�v2�c�u��5�l�@Pl����B9��f���}ePt<z/*����7��(���L��(�x-	�4�E���¼�����L�Íhن�o�B䍠���>����&zܣ����UJ�s��V1С�X�j�o�^w��C�*���x���`;����
w6���� �ppc;�.|@�!���W�/[���n.W1fP� �(��fVԾg
)|ZP0�����U�{�
�Yyadz~����D���q�z�("���*�v%���	P�n��;�M���"��.�[�7��H 7E�FB(gYC$p&"5�A������k���ы������N?y6�:�*�h^��)P��A�@��j�양;��_"���CC��ڪ�wBa��tk�;4�V�\������R���B_̕���2F��+:��֪��Kv�SY�c- �� Q;G�l�-���L��`����9x&��A��%�!gmi�� ��Y��g��qo=��X��!�ʘs��&�F�~�G��x�w JP�Ld��3f�w�׏�C��O,�_r�Z��D�E��tRp��X(�Ԙ�؎�A��y�Bݳ\'@2@��D��6�旜�N����8���Ğ����.�@��`�Ljsl# E��Pem�g����jV-%P*	���S.��{��42��qf6�W���?���[S��s*JȆJI��3}�,g��ҋ��k"���~i��S[��!D�"��@X��$������A�y��P�MiJJ}�߭�ZHWu��J�`=��!�.� �Y	Z����΋Le�#@�hn��P��n�՛�f���A�N�c	~]��N�r��3��ny�q��&���y�*�T�	��@Ym�y���W�n6Tˢl�ʨRF����Ġ}�0����I"����/��+O�Ϣ��ٙ\yXD#�����а�,���$�����J�O�}5fHE�ki���M�������To!����ȵ|]�N��4+����M��.�"sD�g�7�7�P��A�)��4xp��C ����)�:5��|�'/��8�ˮ��'��$/hW�u&�q�
�\J���,t�!>]v%�����A�M'����_�\�'/'�m�<�����۸l���d���ppb�%�B�g�+��%Қ��G�ѢSV�-�;���T��U�?�j{dye ���я
�TX��=�uqo�K_A)��d �v#�B��A<�:|p�,��B����{!�v�X,��M�#p%ɄFC����q@G�׬�uYR��9&��yzl���ݍ�j�-�is�#)�<b*�kkD�}��;֎����> Rc8	2W�=�u�!gʑU9�\��}�OFJ2l���>�����B�_M��O�����F|	�)'����u�٪~����|���A�6rʸD|��pQ�A�'��2�؋�Q�F	`Ck�z���Q�I��Ѡ�ߦ���I�s]V�vId�X�G�R@>�����_�y7mU���;������[as�>2%���N5H�>\�M���#z�p�M�u0=����y��A��o�3n���>L�Ѫr�:�3����Ƙ�z`(\ɫ�+�rH�j+}�?�A`u�����I�e!.��>�N��;��n���]�֕lw�	�}�v�=�h���=��R��2�ı��7dվz���R(�0L<�Y��`^�c�Z�*�	�V	-3됦���}ݗ�#�9I�"�$��9HWq�QY����Z� m����x�(� �3��#�
e!�T�X�\���Q�.� �n�K��Q�MMޖ����R� /�_�<��Np�ª�� N�E��0CbsE�TF�Ht�?�Ń}�A���om[3EM$����L�-t_��mJ�x�^-�a
���:��_4���%�Cކ��fm�F�g� ��PQ�{�/�x��w��Z�]2�"d���JZ�����6��j���0ܩx��iM$�g9p�~��!��ò��$P�N��IJ�fD��5�`lg@� ��Mc�wse�#��,��[;���-�ڒ�`���iY=
��=ؒ�a)hE�����t�@4cͭ�T�dt>�?�@����&��kr�5N�^�9-���ʶ�I�O�j��#+�R�|?��a�@ʳ�k�,�(����+:&JU�1Ŋު��6�+~�O@����6<��A��n��*ۣ�s�a�I�4��������"��K�'�X�K�T��O�R�!p�H^��G�^������)�?$�)
O5�k�&f<M�0c���7L�Z_�n�6_2�u�e��W���$�9�݂K��*���A�K�Wu�[9��LQ���w.K�1-wY���t������b�T?���s��1S	o���ŗ�~� ��d�Ʒ��L�+��n)��0�D{������z�BBl�w4oG������+���B��zY���Ѭ~��~'0�6Ghi���	������WI��=�8�	�*Z@S�M��V�~���3�'��)N^X���锍��h��-����Z�#�-��j*p]_�~�A�������x!��ą��=P=[�����硝6�K~X��J(�z��U*���;�<��|�A����M�k��o�A��8o��]!X���jOk�"�?�6��X;�T�i൶#JXT����OWN���X'W�@���2J$�_c�7���tx�=nl�<�Q"d��b�)��J<�fcgvF��rr���'�'�����
��;�G�Hf�ܮC982�/�Ǝۦi@-"$o��B����%����-P+����Z~�1�����k���c�T�=�R�#?��w�J�_���FϨ��eh��#�P>��u�X�U�5l�X�c�yZW@�H��U`Gbo�N���*>d�@����J�&���'�8�6�7	_3'�y=�?��v/~�]�1��1	���v�N��������z�P 6��OC�������q�&,~#��2�%�x�����q�f1���o������rwK�ߌ�aqi�e߭|���x���:w�.��Z˷�w�5�H1���kX�Zu��*d{�����z\x�Dk�,��큖��/T�%����Ⱥ��b�I[�J�0)�9���K� �cd1��Ak����Z#���ȅ��e�{���9��.���Q9R������(\8n��93�um�=��W[�C>��:��*+4v���3s_�N�k����ƣ~��a����PCN�������bR0�U���Lb"��)���o�&u��7�B��8�����\m�8F��kc�>g������..�'����l�#Ȑ���1C0i?��cd�K>���T �H�#��AqƝT�pZ�"@)����jW�4U9Z*n���pQM�Q�Yk�������S���y���#�&��!�Pw�Qe���H���-"�-z
X�X.qWrJ�PL�G�ܹ����@��(6ʮ&SĈ��ݽ���@t�����q�{��ݤ�K�Z�^tkU�uQ7���v&:�e���s':�t\��VI��� s�<��-߀Ň]��-ЍU�b`u4Sڢo�V��J����+���1qȅ�(r��9E�Շ8�~�"���H�ŋ��8AGzD
�`�3�$�6�1ilP|J���k��Nf��������݀����X������qw�{����躠�����U�j�z�*�@���?ߠ�Fj����1�,g����Y�eP�!	��9�~��ۍ=�Z��8��P�.pU.M�į�!\��+Srՙ:�3�W*����&�
H�"�a�=~��Lp�Z�Q�
�Zm�{��;<�h���#�j�Se�+՝]H~mT�Ip�Z�i��W0�����|���y��T�Xm^�&1.ڞ�6)X�q,�
4=�1Y�SY��-F@=�I�!��j����	Ub�N���;�p8;o�n��QįϾ��/�������裡_�Է�Z�ν�ҋ������Z҈�;���t����q
¥O��A�N�=ӹ����52��^�X��<,�,
����"3a��e���W��e4ɬ/Y���v#Y�%v۷��W�pt[���-�p�Bi0�j�k(1Kg�aş&��t�9�u��q3��D1�`e�%�XE��pv�w"�u�Hh!t��k��f�0v�>��M�H):�V�;R��GJ++��Ǣ���Ǧ�y�k�J�֕<RQ��R^ߟ�܆��IL}{����:#�C��d*�������:vR��եC��li	ޫ'������-_G=h��u�o�b2�W��.9�u�̽�8IT�:�g[��Z�.����`�(/N��[~�����w�3t�+*�ԟ�t�'>WOV�#`Wp�cP]�٘G�IWjΒ�g���801G�ڢ=�
�7)����[ڧ���O<+ӡo�nMxO���rB}!��m�����Cm�u��9��k�f|�.�Φ�Ft
�c�c�|���rF R�Ղ�%5����w�Ђ{�,�[vZm�`��y]��͗\������%��ߔ�3ZO��V�EDa�@=����:1[�j1R>
��̰�e�uZrAk�6��8� ���Y�G~��(����ę?�~�Sc���	�e���,v{,BUiE�����-vz��}��r����o�e2>��O_�1�)MfB�����_�u�Z�)ݙ	�J��LK6�f�3��5b�\x��D_b`�s$�Gz�l��o�~�C��)$�H�'�d�b~��x���](�$*N����%��2���2�*�
D���`r�9�}]L��z�d� ^�]�
GH]�6A�{��d��@g�b`s����)��r�*} ���-�}��v�{a����=g�̜� �C��5��&t�1z'�ۯR��a���,\�������sf�o�^F�Ejw��kx�3vL�e'A�z(��0����/*K}>﮷Q�����]���\�n������S=C�i��ю��G�!��jEǟ2�n3ğ�Ս�>Т�ӊ�%���#іN/:���u�T�Ǽ&("���/�O�QW͒A���I*�Amİ��ɒZ�P2"�4`�ڡ�B=�V`���)���#V�P�9�������ʨ&����y"�)a��'�l\r���3�y]#����n�KR&U��W֦(3{���j�j�9�j��
bk�`�Fl����s�0�oON�	�j幟 #�jžk]U��Ά*���R;�T�Y���*��衩����#�-�\֍���J2{u�E��i()�#M�n�9�a<�WS�u_^��`-e�����"��K0Ϛ$�'���s�Lك�kB" .U�)]�����e�F���͈�?�>U)2���3ڽx�V�#�h��S�j��F��Q;8�<�N�m}��,�+�N�#$��m���v�Se��}��B=v�zQ3'��m����]�L+�`��yX�	�7ՠ������؋�R���Ь_{�B��P��g�Շ�U��<{uѻ����$�JWx�ȏ6U���e`{�2��F`.��,qQ��֔�� ��|_���V[�SB�޺ ���&���K���a�n[&���:'|���"��;���B�Y�/Oi�4��Y�Ƕ�:�Uy�]����
�B:��^7���:���
$bG5�s��,x{��J1���%W�����y煮Z1�?)U"7O�n��v2tlJ�U�YIQ���\l�q����[��0]J�Uǳ<b�m�7i�l����%�����c�Y��c?j0��& \][DPZ���#C��d��jħh��*�N"@�ų!�#���H�2�:tflK	N�r�K�T��"�%�N�k}pD�%�N���(�
\�xZ�>�2EÀ|������&A�z45��#2�͠,c�����ùS��l���<������%��.j��cãs��3W:5�v'^G��l:Nq�'y ]��3��LZ���4���=�ǐ���LV��6z]�(�&���(����7�i�
s�D�)h�����&�nAD�I)�ra�ɌӚ9VdG����ΰ�@��ԯjcZ!��.n�1Uݿ:��J0���Q�wp�N�"��s>T���
�qY�9���2�}�y�m�B��^�|B�Ճ���9w�@������r��C�` c~ �@�
�m���7�	7�*���\a�*[�~�?kd&�WR�o�mv����YK
��LO9� N�6pB�fwy�@�_�����{�Qp�`Ӥ髋]����Ade`�
Hk��5��	���l-���4���-�T�%��'��Q�쎸�n�V�|-T��<B�;�����mf�B��{t�5M��>e�*4�W+��*�(�q��y�ʕŸ�jkbzK�m���b��G���|x���3m����Q9��j���%u��2�� ���TۻN���Y��h�$���1?;S�p���Lf�?�0lr�R��O��W��:�;�˖��O��g���OJ�|�bOq� 5N(�Qzs9�q�}���k��h�>qT�pX
�ȍ��n�0�����H+�B�ǭ���
�J#�.���Y��Ƨ�%��E#=�1�5$)�:�u߶�Pr�5����u�0�NF�Y��`g���獏��ixT���E�� w'ICzA�f���ĉ]����o�ꬹY�_E4��wء�Ȇ�8	��ۭ���9ɋ'R��o�E�e��� �R٘t�kIe=��5�0��1�-t�<����-ygv+%�̡�C����+���|���l
4x��2��cJf�q[����
�d�v2oT�c��s���9U����T�E�fq�!��x����l"�[O�X��("ڂF!L����,�1�B^�` Xv���@U�kx�����}\�o�~�#�^��E����_�4`�}A�u!!/\o�����,���E�Z�9����eCcg@-Nii
��1��u&H��b\������&q������1��fY}U����.B�"\9d5��߱9�{��ge�`4ը�Gk�J�j�+z'��|W�qS��Q�Kl�l���v�o?��{�Qsd�M��ϥ�����.θ��a�j�����0ɉ��<�I2����cP����S�x������'<�kB͚��G^�X�+�XY.���zꐭ�ӄ����a+X]�K��y�V����c����I�ߏ�DѐL��G2�����R4h��W?Ed7�"z�y�2�@��
K`_+�Bـ
���T0G�G�
>P5A���������B�������I����/#�Nb�-CP�-/
��Rl�wd�k��.-~�����{)Y+������t��M8)�-]P�)�7u����%.,DX�����N
B��_df�E���^t:��"��%�݁�-S`&Ŝ���=��RDU�:?�Y8��8�世\U����ji�۹tꎼE����T��D!��[��i�!�@	�<�'`�b�gc�G��dU�}"�(l�5`	ϐ����*��+C\�ԫ�e�DG'-�4(|�4�[�5B���ѐ�)�}~Պ�fE J�f��
�Jc��xɺ7YM.��/O���Tj B���m�F��='X����>�z�����/9�X���K�ی���x����t΁��#�$^���j?��,��?��؝�r=tW�gȓ3��L���Au�H2�j�^�m����6������R�A��Nyݥ��5�՞�?�#2`)��}�;�3\:���HG���? ���%�vJ��@�֭>h�'4�c�������$#2cf�~ux�3�0�3�����y�xR�&�Z��:��&�/��alQ�1=c���4"��N�q�K�>즀y��%����j�$<s]fG�YA�QN�m��)�zՑ����� ��r�߷T����O{'�d-�_�?�&� &6p�������OB�M�n��/>��{Ӡ��޽x��t� �'Fn�Ħ�>
!C4�c�O<�e>�2�A�A�r�u�e��K8i��U���� ����p�Pv�֡*z,xr�S����� 9o�@���GV����r���|\dC�����fO�?N���I����[ipjb����������,�l�i
sIR|��ޝ��N_cI
�j{䰙<y��`�GW9���������L"����ȴ�%�w?*?=9n���^�Q�,�;O&r�M������]�$(��n�_LL,C�h7��o&#Y	"�������	��A4d��TX1���R�
���n��Ί�������QK�d��L����6��@G���P�+�vl�g?�@��M&���+��8bg]��$ڷfWjZr�U�WS�Z�d���.�C�8�����R�������^ܺg�^�*S
�4<��nL��D�Nt�׋~���d0'���	�N&s��;�E�D��xt�{z!�$ ?8��ߐ����\EJ�\	D�b��<]�����
��j�n����mZE��b#��q^����T8�����r���KTyya'�ZF��jH�ˀM��2��ϲ���%���Y�
�S���,$���
||z�i�BF�I�MTUa�L�?�*s�sG�Z����j"�=��8��O��Q�;��A}*-�$�[�4����D�(9�����o��O�:Ы-��Mf�{��t($��ֵ}���u�τo\Q��þ��K�?����/�i��Ј���5{�)2�r���g�����b�o�XO�|0��v�Ib��։���wBNi ����� �+�9@��V	}��x�,k�F�X����/g���u�T�GC)��_L���^�����7� ���)�<l�죡k*q�7	��^�{�0(�k��}�=��j�n\�]NM����5}�p�������ܒ���v����=4��g�0*Cա�׽f� #VH9��� K�H��302� �D۴"Iب��	�1��2*��� p���.��']�D��ڑ�6���4p�"<����tBMj��{�ʍ��d������}�*����t��Z ʯ��ͩN91 q��;�� d��> J疗vn�3�QHS�nⲐ׻��-_͇��ّ�əK��d���xk��A���aҩQ w� U�E�1����_v�7� 5�����k�U�QөKk�q �I�A��| �j���	��w�vY6X�����Æa��7�tR^���	eN�U�BW��%i�`r1��C�mw�/�3�|޻�ł�S���D	.��.s��U�{F)l[��-�#�6�;,�b#��ʯX�}��"���-!���d�YA�K�6-����H�,���Fah=<f7���:Q+g�:r���,AO\�V"B��~����ۦ��R�X�w=Cus-�*�Ґ��3÷Y[���ʋ6FP?M�_~���n�Al�ﮢ���^.@�5=��NM8BU��S
<�8e�K/砐 �)x�-��k)KnF���:��D�����љ�(T>25�&�#V�EGA{DM �[��vE#5�`�J3�jj�2`���5jJ�P����tk�XnXI�*CsaR�i��ˀ�I���dM6�,�׃�k����aVʁG7����:P��Ӎ���'ڎ����o������FE��$�?��1&��� f5q�d!�l�%�u�A�5�2֒�K�{E3ݥIȋ�8�}x�������{�Da.�o���)��8�Q=��J^�̏Ћ�խQ���/��
����f�3+g����U�e�o(��DvK���}�Ͱ��>����l�F�h6�y[B��.xV�} %����N`�ި� ��7�e�\s�y�������f����A�KcD�][h5�Dܷ����J��3�/�)�6#�NBa�� `(����I�qMN����1Zg���&ܘQ��J⇑):��>�m;)���8Vcxe*�5)=~Tr��i�#��;�,����L`!����Nq���Ǩ�4���m�q8!Ӡw_�SZ<�0&�9x2�E[��~��9;�DJQ��X���@{�O�?M���X]#��ME�g��g�B3����O�Ï+*Bf�=�{�^�(�>KW��q5j9dn�T��~R)�z0�� �� +����b��§�V�����5���,�Cmp��TF�4�_�3L@5�E+���a{�L��E'�����U������um����3��El�]��4�x��Lq�0��?`��1M{���y�r Rk)��K[��	���#��՟T#��"4���{F�Q�>=�i�W�ľs���51�:�Y��b���uW�����&ȷ�^��.�j/$���J������vr���U��O���H�p�Nޏm�k��x���ޥ��-DN56�t)a�k���K���(�ཱུ��r�"╂��#��,��{rb4=��>�;�P�C��	r_74<kr���F���g0�\�h_:�mi����E��Z�����*i?C7=91�Q���/	�y$��H4��df�/3
x^%�zNىJ(�1蔯rK
}d^􌄡o�Wl��M�'�t�	r��@9�^H�W�����.�
@�bݜ�B�2�����Z7��[����ȓodd��"=�5��lT�1��Y��/1.�L�,���٩�[J�BK��;��|K�Ӭ������W9�p��"Q��~����7�ź J�Z&�����wT:T�T����6s&Y �ywx�L�
�b*���[0�p��P;�/�x*�J�j�ށ���G�5�n��3�Ũj�Yjj
�)"+{WV��E�1�7���Z���iw�f�#��8>_����>�"�i�tǢ�!�!k<Txn�Rg)��d��s4��wc�IJ���^u(��η���j)���������Ô*��og*BY���f�˴pB�[��3cc L�^7���۰��K�� LG3�r���٪�X3.h�8x��NR� ��Ɖ�����x9"�9�M�i��0X˟�y���u��^〄� ���2�)�ѻ�3�ZQm���3��:���b��z0��XOW�%�yV�c�0���iAY�릿�:��׆�@���Z%�C��>��pe���S�U$�;2�ms��-U6�����_�?�m�~��Hh����r�l�4~�e'Ì���� �|�<��AX�h-G5�Y.(Xt�x^��C�8"��e9���u��������A�����#R@GQ�9}Q�ܴ�B��q���TD��J��8<��vzu���T&�g2cS`���=�#�>,�Y�˻��O������u͏tL�8��]J�E0���!SH��U3d�����/��X�I�?�y�~J�R#���o�T�NF��"Nu�հ�n�ZH�4���h���;�ڟl�O�72X��;M�a���nwlM��%g�� ��N�U���������s�9��&<l~�ctÅ��ji���Ä'��WB���ċ�L��q_�T�m�bkr���^�n��H�Ac��rI�t�s��ĺ��Ģ��u;��|�c4}�P���Wh"ph��OR��j��=�jv��e�g�X=0x���a�z�M��V���z]�\9>�޵ :�J�{gF:l�Ir�1Е;���ޭ�뎯b��~�gEh�(�Ϥ��$�{7�(V5x�����'8;�&{|��K����A[˃�)Z��r���PD�a�||=��gNv����83!��������'�HN%���&��P���"�R���;�۲�1���w�u�����6���Ր��lb���a�WHL��
�긽-&�'~���U���Xk�-�6���m��0'*�� B��	�2G��3�5����������&n;���|jT�eۈ;~�h�s�Z -���%�����^}�A$���bAGҷ��x\�8ֽ����'x!�[f�􏰮H��Y���5�Y��I���SK�~B�Lv��#��U��6�u�� �9}G�|�Yw���D�Ule+�KZ�ؽ��IxL�[�wF�&��+̚�D�M2�l�;��w����7r�	��o�h��h��̕����ַ��P��cJR�� }���»�8�y1��''3���O8�f8���<),>�AL��a���|/���� й��v`�^(�A[���@r�:`P&�d�J��D{�f2-�*��.y���@M#6��C��ί�vF����1Y�*%%w�������'�����5�J�\}�
WT��,y�n�p�|WZ{�
�;u���qp� �܎��W[�BtǦ�<���(_F7�����4�h��«?}�eɞ&�n��=h������єC T��EJ/��y�kO̀���*���¥��	�c������:����PT喘���q:�!�'��·@h�J��e��n�ԆRqŭB���,����.A:�%�,�@ht�f��eQ�������)u���u!^s��E�N_���s��sP����dE���u�=���X����JAO��A
����BŠ��+j�k�A%�ba}U
)��FM\�n�j����&fB�|=F���D��b��?�yz�)�`O���	f��ī��]r��0G�!��}Di1��e��@����6�D�B�V� �$M�R����gU5����qF�t�� ���:�9vl���F��_tK�%�{��:�؀-�3��njL�*Xh��Ld?]�עB����L$��B���ԗ�`]��
�Ǎ�\C���ܼ��/��5e�����Y�z��¼K�b�7����c�(��ݍpj�M�co���2[����r�_t���s7�q�՜cw�Ȟ�=S?����ܾC���aɮ+)�-Gŭ��XC�ul����6K��(��Q�s�v�F�K����2��2k���}��z�
=�
)��̘�Q�b�������}��
$��\�3!�C��~�7��������ڙ��<��~!O_`5��le����<("r�3G���Qq=qIf� A�����������Gk�\�U'Z@���{��49e(��A�/��zF���WQ8�N�c����\�ݟ?yP�4�76�)����`e�����Be)0��\��2-�;�<�G���>�X�X'��~^l�T�:��}�Yq~��|pȅ.�V��L_TQ�P,�Y-���&U�dq�Bi�A����66B)[��`����c���bY+m����sT�ː#c���gK�`q��o[���!�\�XE��e1��S0�*�9C#��M����P	���x��c��h��p���`�_��æ7{���cD�ic��c#$��iz���u��g��8��ᨎr�TVD;\$<6��� O����=�0U�q,�x��d�V良X��/&��\�AR�#��&�C�iJn��8R�Ҝ%e�F�5�S����Dz=�=�E{�ZY�y>�s���]Yr�����^(��Pu�R'�2�i����?�:����Z�'��r;�l��߰�;�y��=gצ|�Mo�]�� >�#g7FE�`�ME���6=��U��E���!���[��?���ؙ��OV�3r�F�k�X�d���%)³2e,���^����b�l1s���b��y�<c��Č����X^�9�D:4�AT֜H��ga�C]�j'�n^K,�a�M�Ͱ	����6۾���Tb%7����=
�Ž�|h�^�<d���\�ѿ�QU[�Ey0|�7���y���\K�:����j:�mq�&r܈�Q+�B���HsIYtX�����ho��H+nj��{���A����t/���u�;-`ihs�ퟫC�=CcY'��Ս�J1�}��&��\�"&>�ܠ�ЕF�4+�U���_n:�7Oi(?�����cQ�B��v�Y�Y�/�@�@���=�e!�b���EK�Z���%�x�6��KM��Ş(� �P�R�PZ<�A�� �3�.�`���qo?�Ҧ�F�Pm�"��b�)���Y@�gC�3��*�z|͆Q��w,���Q�%�%��s@��n�r�cGe*�� �H�V;vC����`�Ya��1��x@���)�4�ܶ�B_���~댹㾷Y(#�ܮ�̶��>Y�+�YJ�:��� �ĒP}�<#E�ř0%��ƙ�}Ȯ�U��v
U����{��()����m��j֙�T��]P����L���+[~_$Ok��0u�p]�R����;�3�k�����"TpL04�z���$S���lpwD��}]��'�$U�O����X�Y<(#}����J��G�G���A5D&��K^��:oK��e�
�v�l}��m$��``-vy�V�[�WT���Ll�b�>��h�}�/�m���cxADh��
�k�fI��+�X֑_�Nn�O�[�@����%_`���4tsֶcj�ς `�MtyV������we��4��J_%[�k����K���MM����s�a��cx��2��~�츁���Al�'(s�Q��n�/��u	���&�g���s5�
9��)��v�d!���k~ӱ��U��}m��\�JOe����hz��^���dYJ�<�r�lԑ���A����N�0��G����l�La8lD���q��Y����|6eGޥ���b�z���!�I�Z�sڬ�m�*���
!-	�F}!���$�c�=�s��6�цz�X%�'q
�'SJE� ]�U�Rc�r�#�/b�X�L�	����EhX�Y�K�I9ZJy^�U�\����0K��}�������#Y=�@ ���5�:U�6Xs�)�F{�@��lsI��ȓ4���#��h
Uyo�����GPۀI�N�>���Z�:��E@OA�@7J�Lt��0s#Sǯ�δ�b���|�[����<��E'��꿋s�����7RbAv��R�=s� fc�\fW�m§v~{<���ߕ�@_^��>Y=J;͟��UD�t�M�$�5U�7�\x�6ux���J��a�ͩn�Y(�"_\/.�W��91�����
��|���.�M�D�!#���d_�a+��5qu�+�[5�]���9@�lqƋ��}N�B�T�m�A��)HqU|_EN�4�cS������!}W��R=�Ե#�/I'���C���v�A/��%�8�-W��Z�@����A�=�=2�O�}�K��kO�	96ڔ�M�L����\�� �ଃ�0�[_�.+s����bb����''?�z�I��q$��$�g��G��`�b���R_;2��W	6s���|�Ś��͘��Pd`L����i���5�2�d�i�NS�B����ge_�����F��u�ّn6Ɬދ��ޏ�τ[HxP2�<�M~G��y�
qʝ�N|�\�	
�k��}XM��$�}o� ��� d�+aZ�x}.���H�y|��;4h�����A1&�ę�~t6�k�"шO�*g��GѠ<�<��$8lX�_Q���Y��"mfĬ����u��m>D��4���Y
^K~��5+��(�X�br��d&�?��;�6Jj�\���1X"�!�oP�8|��ypzX߆嫩�����$`�����Z��{�Za�K>�_�\)�i���x4�o3@�b��ȝ4r[�YM�vKp��pc���n �Bֵ��~�� 5�+=`M_c.�S E$���f�4�3c{ 0G���c�Ã0��d�����݆�'� TYf4ePX[ͯ�0 ]���J���SE۞n|���*��7϶����n��n��H�Pe0%ᱪL�g�Y�3���bQ�q�ӿSU;��y�U��ʢ9c~�js�|���]���\��=�>�ҳ��|9/v�@|��`��9�K|6�'���sv�;�16�d�{?��'�;
�����(�+�]!sG���rr�ː��s��c���<n�H��N_,{k#�N���)G�
����k�vRT���<6ѧfIgj��;�t�6`��^"'I��4R/����&��4ϴ�h�R�!����EcD��G��Y���;�}�4m�_p��V������h���8�tegC3j&E�8L��J�|�cvA�̍u�rr���2Q��qG���@�w/[Lb�2F�3[�?�����B�}/���+W�}l�?�3��-���;�
D��>��\B��j҅~�۰��7z�[�%�:��|�f�2n���"����
��n��)�\4Y��&=���8v#X#uC��Z|���� w.]�(�3�����@���v�z�.�#�v�LZ�;��.��j�@s��v��X��L^]�Y/�s�����g�,�pT���h�w�4������!�)��a�k,��5�����X���p���(�����W�/�3'��얇o�.D�n�S�k�a��޹w��@aF�����v���E֤O�I�ڄ���X��U�����6���cw3���h����0̕���}��	��f]N`��B��9m�͍ʟ�u�&����CD�����Nڅ�5��L	��e�ONp{G��%H��i A�q4�.��������V�WVEk&R堛�������D�簑��?��w9���[���c�D�΀V�˔�,�����YZ{�� �~�Й�m����@�����n�e�	׬pNW̮�/�w7W��"uj��W1�����z=�d��j��3�(ꎜ�b�I姃��پ��>�Eg+J�{/�G�d�4�StQCF@�����I�Ѻ�E6I+ûk��~���!��`=O0�&��V2���ϲ'�g�.�9黖��{NR=���PL��@�m^/$x�1��������F���8<5��W���] ��4=�6zd�:�0H��C���S��9�c��i�_��P���:����wUs�2�+��A�*�lB�曧Q�ӒkQ�n�L�v�����.����?�	evV���� ӓ�"����*�J�uӡ$�s����s�6�U&�`����;�_�k͍ï`�ҡZ�Wt�ma���9p�W�M�Q&^V�����d�rʶ�Τ���uS{�? ��+���0��9!����#��<f�Ϣmg	YE]�1W拌���D
�)���$%�v{��_�~�����z_�~�$ʍ/��t�^��	�o�j[�W-2��w���C�o������Xoh�i�1w�䊼�KWkn0;��k�ߊ��.� ����s���@��#�N�.��¢���	ų�'^�u�
7ێ}��u��p��D)ؑt��P����	���6Yo&����a�E��S�VtcA���s��22�ۄ�K�EG�ا�u��g!�5�[��yǊvd;7��,��cmI|he8n>����Y)$l��Nޯ4�M"�rSW������Gc��3�)���ZЩs���k�� �Sy�8�A�����)0��T�!i�d^tr>D�~5�4�8/e|oW�p����%�r�7\�\w�H
c��3���~%�wR���-І����.��ǰO�G^R��OPj�4��D�/|�N�����@���W <eW���K����A2i���e��L���x�j��F�Ӯ�b���E���ʠRSYIhB���s.��Ȋu�&��.���-:�C5�u�<(��d_ޯ�?�qA��fDO}�u���Eı��Y��D�/ �9��>���^�7k�4�ߜ��wS6�"{�x={㌟��^d�0�)�@��Z�����%�-�j��J3��;ƕ�o,�M�4k٧�9>�+��!7J�x,:4��u*UW����x>(=P�>S�7M2x�3j�_#m���<�C�c��w��i����s#��З��Nc��>Di�kױhe�ju�HQB��^��ꚸ�����+�� ���iFr��'"W����69�X}�LIzW�nbs�i�������co(?�[W�	��_Pb�ePi�xf���2I¦�ݵx T$!GQ������2���x�p�/��ȟ�i=�"f��A�����J{��}4,��T�R�F,�n���]�$�nu��x����}A�C� ���_�g�S����\Y3�A�X��m��TR��] ��H�+]`\@����78#��*��5Ig�Y^�3�߷r"��S�N��^��r���o��u �zO+FI~�2k����:���X���w�7���VȭϠ��}�sa��X��F�/�m�� �֑��\[�nVҤ]-t�RɈ�^�E80�ⴿ�(`h>`Yt.��67%����Y =�e�?Z?@p�;�S;��K�^�PVW��
���-&���0D�k$�&m_b��T��X�)�����&�x����Yu�eO������pL�.�@|�����7U�}�,dpC�G�ߎ�]�V9$D�&���9 V�[ɘ@H�����>2�����*��9օ�{�ui�p�w���e���\��h��e����e��l�!�<uE��El2����_�*�����>���
���9n]�ܐ���دL?��kq4%�FK|;�(<6`wHk�u��U]q��C��|t����)�U��3$�I������:��.|~%.��?؂�JR�⢡��W�%M�Y���ǓG��1���+Ctfa��Jx��%ͧkejIJ����9��xu�5����í0Q��u&c8U���ն�L��c�(��Rj�KQ�����#B�lY)��]���l���w�sR�i��*%�92��"a���0���_o�~�)%0wʹ�%O>�x\��� �^c�:l�Λ�V$��XN9Bj�<M��K�KZ��t�}�ѥ|�����f�U���E�ƚ�o�T���T՞�\z�`c��}�D�����Ú;[�@��Z� 	q���Y���b���&E���<B��m��|��=wc�w�\�;���
�T�ǒ��.���⋔�ѷ���qZ2������o�x��h'	:]���k��c:�xY����q��ٺ���"�Qn{���?>T��H*�Һ휇ꃖ�����!�U����dU�����~��4W��dW��ן R9����f�C(O�P6$t׸��Ϗ��^��t�E�!�g8�m]SL����{�M�H����lN�?q���GD�~��-��Cb����c�y�!6p�f��0}��5�d�xT�+�x� Z`=R$�R=m�K�Tr��wmYc"	c�������i$F*$�Q2/G�k�D1�b�j}�)| !�)�'�f�s�|�_���Ku��5@8�����P$K����|GeKF/ꎦ5�$R�nVmt�Fx(��`��p�tZZ�����݅���|<!��jx+X���앰�}~���Iq�t=�^�A�|т��W*��!�^<`��c|����c,���D�wܵx�'��6}q��ى/4���rݟq�_�hy/�݋Gė2F�kV�	8�/'a��3je��P����E�ӌfW�H��<�C�m����h�f�~�����ǖ	��	������N(_4�W̼�$y�T\�/Vhس�5,�ǆ�a�HF���N����:m�����rJ]�U7���s��~f}��ԥ����S�$a˫'K��{���T���˺*�j	ל)0웓5�Z��íA���v��QA����y�}��$��y����':Y��(�Պw�^���I0W���n�����}E��<���pT����a�{�,knS%(��=Em�;�0`u�;���i"�U�b�sHТ[��'��Q�9Wn�P���Fng��&����jAt�'�$[jb�$�w�eV0?oz-��-�Y��!uO��Բ)��ݿ���=TTƊ��β�4N��w?f�B�5���Y�<{�_y6�fÔ���o�G)�(�(Bi)� ���	|��_y��h�L�rI�.��i��-<=nn�F��|K��� ��J�"�wo��^M�z��j�Y���6���ߕ��W1�,NL��T��� ��&�
vT�ȧ6�y�Xt��j�7HkJ�_C|
��}��H�> M��ؑ ��e���-|��9�vbSL��84Hn�X�Z��}��C����������(�n���0@���DZzv��hW�:��mǛ0	�fR���N����2��qN�u�t7�s#����K�E�O���t'���X
�����>.�{�@�u�~� ˮ���d��)k%�!^A~��:�n�`��yj{��D%�BEQO���W�����9��Mـ��/|�z� �/������Q��%��>+)C�@C�6;���kd�E��GgP��i�6��@�1�Ze[,}�����/ZO5F���)/���ӫU=4����:$�� ���88M��*Q�K�b�j~�;�+�(�v^C:�[*����	����vN�h��:�6)���c.�U�|&i���^��!*��IWY{�3��38m��Z�vf��K��J5�գ�\<�v�rd�@�%�����c�|<2�����6W�[f� 
{�*40G�#�F��;�.iJL	���ubz�疮?����l���Qu�EY\rZ��?��v�p���5XtU��(�s�V�x�u�i���FV���-��sl��U���A� �M��vt~	��&��2���}m�|[ �ዤmG�s�4(X/K��P�T��÷yo��#|��ִ[��{P���SlL�am��5-�K5�T1S��}VG�<��BL��������ʍ��5�%�?7��r�,��ݾ+��w�<�Ċ�q����� �O��uw��x�i��}ٝ{R�Q�<:����ט���9w�!��-Ǎ��U�Yt�a[V�A/��Jt5R�� %r-Y�gp&Cg�� ɝ�f��X�V��g�h�6{�R�}�o^@h��л\����t����)}��+M�s�1�c[��s%���v�g$��ρ�.j>����_$y�b��	_���8��՞\����W$<�}����Ѧ׹K�2��q�h� �Ώl��"�24p|���8�q��cC����OR3����J2�ux>#'OYta!J��j���z��og����,��GA`�\E�?��Ů��׊�LW�&�ɪ�"��j��@��"���X�k��n;��������N�"v���tUNa�	���r,��W��8�^�u�;�)j�uR���K�\��#��٬ h
������X�Q�m�9�`05�]����|�J���L�!�����l�7,�Z����պ��sl���X��W�\���+�y��q�������\o��U.-�-M�Yv[;�S�WHEЬ'K��2��HS�*R�<1�PZ�E4b�N��K1joC�8s�p�f\Ҍρ�6oВ����9��s*��kx��Э��6Qu��?W� q7GYTG�l���/�zV���#D0��Ԓ�-�k�h�9N�8���b�ڪ<\Kݟ8��?�z��&��G�=�H�=9��x�+փ�һ�ǥq�,jO^/�[�^kP:�^E�Z��e�'�	O��y^�����Z�w:L(����}�?�����cM�I��q�h��J�o�\L��P��`	n��BK;����߀y>%���(^"��[���H�
��|��2�W׈��oˁ�D�f `��M�����ÖR7��u�2B�x%��& �%��ܔ8�H�q~,�!8؝�4����zխ���be����ɸ�{@N��b�w��*��f���S��_��x;^�y�j�<�.Ç�����f~�)���W�k̛��Y��|�������040����ͫU�^��5J�J��Y�qPN�u�ex�/��M`����?ۖAf��F��ς��w�Ę���NMX~� f��8G!��B�y�@y����C��yR�1�� �w\u�I���� %�����0v����+��޾�RM��៧�E�{~�L}c�^�����B �%m�p'@
��&2ޞuʭ�5Ea]�ew}*��eh�٭0�~3��;��p�#j�=L�+�G��	���T��Z�;�K��(�p`K�*���\-�����;Ȫg�x�ݙcr���.�^�Ͱb�r��%�Z�,/�o*"��[j�D��#鼶�A?��Y:#�����P�B�o
��K�7,$#��UGB�׿@a��P���iETƭd�G���s�%US5z{^g�%�F��,#�_]2�y�E��''Mx����?;���b���d��8wĩ��.q��."��|���-�����4�MC���lA.�kK�q��w�阕]ɐ��҄)�6i��ޅa���^�"�Է�]e���: p�R�������ˋu?"OvN�vSN�5FI�lt�<�(>�������ps�Q]���R�:�Rǃ��x�_��FH�q�w��b_�V�րj$������n0�	rYǼ�7��T9R��+�N�:߽� 7	�����Mze'��6����Y^�pt�-�
�v���ǿ�>ۣ�	�e��!7�ف�F}N�����g	Jg�����e*��c&��������M�7z=SR���/�!�s��}h����5�l��d�g����q��Π�=�	�"ξ���X���+�+�3X{x�w?2�	�+=,1�=!�R�x��0��z�f�x8�Z�Cz�eLNwb��&\֛0�9��O�׫m��\�3�q�I��8k)=H-��h<�f�4r������vr���Zg�W<�r�O�*g���pq�l׫/V�oR7,��ƧikZk�	~&����	�	�.��qR�h���������ص���>V�*}s���̙Ht��&Q�ѝ��T���mMe����
�n�~�}ş�^GMF�~�G�W�(��v�eP�j�i�T'u��P���^J�����
=��D� �n䫢���p1�$~���P�=�R}Q`A֤1(t�FK�ɰ���(���"ц��՘j�	��R��&J�p�#�ۙ��ʇ��b��VHb5�Z>�(�2r9jd�=�8K��XI��b��+Ω�o���qY*��[��ܲ���Rvҝ�}Z=3ˉ�N��'�IOПo���i
���ٹ�]�Br��5�A,	M�:�>���+y�Q�S�
Q)��U<�&�����
ْ�O� 멺O�V~��g���Y8@�!��X��BŌ^y����q7���,�� Ι����u$g��S{JQ "����3���H��2e���V X���Fk'w(�Xcv��YF�{3�q�둌��E��U�xa;�
�:w�MD�7�6��Yw6�W���H9��bnN�	��������e��@@5pd�����d�z�r,����	}a�bi[M/�ܸ����h ��|���I`O��_�ʵV�+���v�@���i����	6�Lp��f���F1$�j��ީ�y^>=�Ǒ�}�Po�"�A�X����a%O��R 2 4�.��k����"�0q��^�(�칷?��1�NN)8�F�a�,�P,Dc;���u,�챮��8_%��ַ��<��;�o�uD9��� d�s8��1�3C�k�k�R|f���H�7�6-�i��L�-^<O�R�`�}.w%h��${���k�+8��
��`��Z����
V �7��<@�
d��L�7@����Ј�ϟA�6:���^(
A���璚�f^�:���[�%Q���E�	�4�?�A�����U���$լK
9���3��7ɥб���ǥ���)ժ��^@����,n��9�: �Tv^S���������@����B~�Oqϲ]`3?/�����=@(�Jh���dDτ��|Y5ȣ���K���������I��మ��{��>t�H	���z�q�9�1[4Н�n3:��c-Tp���G#/60&i�Q�`Q���6�b\����|:ѣ��{�1�B���-!x�[6s�r��'65p�=O�X*7�;�2�]�b^��,�X�+��4GZ�\����KәZ�\w�m�=��|/�����4���{X\�f���2��%Ϯ��m3��� ��@Q����$?�Vp�9u����V���'��:bGܕ!�\�@�f�ޟ�]��F���AJh�X0���Q�@^���[K
�7��/�$cO��y� `?'	�B��ٛ��ſ���B09����D����4�
15�YX���6tWHD�}�L��bԜ�ų��VS� �[�|N�����8��(Tڵ��<%�ͪ�Z��{8����	g��Vi̐���d��P5ͪ�mՏwb芴��=��ȷ͜g쭨�H�6����q&o�ɧT�˻�X�G��+f>���J9��u(���O��0��y��C�0���r����V�Iѳ���3[^�����vq�mh�Ƹ�8���:rZT'{a����C��k�Ttz1 �����+N��A5�RݔȱP�o���u�녋�b��e�#�v�E3ч-�0�<�z(�.��7��uV;�:���TLg��icڒI�������=h�kQ�o���������0W��4�l��B���H��7��՝�+�w�����@T��<�Ϩá� c���_�`��JK�3Q�Ǽlb�؅Ӯ���qi�K�!Z���rw��e�u��D��<��oͨ��a~��$u�^E�\��Q�UU�D��(F/�����n��h�,_���Fi�E�ݶ�۾��>��~�zZUW���2�� L_^3�9&��J�3�쉦6 HL#��ZG!<@���?���"1*Uנ3{�}�{�Ō6N,YL��G�A��4�J$Y�j[ W�~��U ���&�����Q�� %?��F�K�K��2c�F��eFb�������CSXV:��(���5#4iJ������<i�UA��i��r��Z�k(,v���-6@QU��&�8?x�0��H�iPpXR�T�[?�To�
�P�Y�%���.�:�c
I��Oۙ��DJ����#!��!��솁�GP�U���6FCDbQ �:�����J?7��-Oe��/�f��v����Cy1�	K�������'�v~|7�p�+Ѩ���,Qx�d|d_���n<�HH��
�TϤ�i�H�����Wn�� �r�/��]��G\�򉸥�ٷ���;A�9�,�:�E�|Gj�6�8o���Q��}�c�7^z5~���!��z��^F�"?��y'��b5��/ڨ&Ǒ�৛��G��&��ɦp�A��[x]U1b^���r���<C'�2v=h�K'T?D@{���4�Ӟ��j�����u#�BG@�bDZ��Ø>o��@�@r��!?Fr�"0��q�K���6��ͮE�M�zO�}�BS�1B��n(E��<�L�u��QL���v��w������&��������+u�i�(N;�):���܏���0]�=A��S����+îs��X�s��)b9��U��cƼ���9�R#2�@pD�=�<��+���>�Oۀ���r�ej?��&T˓��p��8�EVC�#�f��AH76���n_)�p��|BW�ʘؖ�>G
�vșG��5��'#
�hD��PA	�U�ը\�J���OS��Xߦ)��.܍B�2 �}�<��>�W�׭�	k	ʳC�/�¾:���f����O��3�._�q��&cJ7��ʵ��9�v'�J�b�B����)��``��N{�j�'�<����ˆj�X3sUQg7K�A^wsa,&�@��?O�M�E��=�����Zl�K�}����v1�Y:�$M������B��A��vV��Æ��OwP�NO�4|��9�g�,��:xY�;c/��AM���SGet��u��=�1QJ�=D`�/��)g
;Ä���� 	�w����!����z����-���
�2*L��/��Xѿ;�&�)�bb��pZA��l�T�(-�����䓲��J���z7}��tZz�+yA��ɕaߨе�H"�fO��r�t��Æ������������/9�.`v���ޢ.f���+X�r[�6�~ ��l�����Ryo����l}Cn��ϓIWPɪ�5�S���������5� �2��>3����Nr+M��u��]�c>Z8�"��5��ۢ�!1�^҆�_�^
ж�b��N� �$܅g��,���Ҥd}�u�B@�^�'@$x��~���|�}=V=RԘ���Y	]��x����u�I�2U���o��K��;�T���
����������9WXP�5l��`(����#g�i7��V"ݓ�$�\顄�e�(E~�n����WĦ���� �+?1���@�\���?3�!�H#��"^���G'�ԋ!�7'2��^z�z�BZ�r�����wwu���3�ȋ�v{j��h5(Pw�}&�6�;��L��U,f��;�!�p�W9�	Y��U�k�:izR&r�d��m�Uo@��]�6���<��=kn�Y &2$J#����p��ͨ>x)��¡k��q��Dj��8{ָ�\!�Bh�$ѣ� n�c�NZ�9�ɵ6�i�\G��88�}	W�7�vC�HB���BRDNĔ-A2Dx�N3�o9d�#I�@� $�hN�oefH�ё��ա/D��.g�Sw�k���c����]�˕���5�6m��䏹�'9��7��
���2�Au���r:�SX`y��?�ܧ��g��/���o���Ѽ��IʯYB���w�X=+4ʱ���j���P�GR@[� �k8n����Vs�Q�Nu�?/S�éX��c&X$��wv2�e��SKC�8�	:��\�t�IC��7$1���P�h���}O�w:H�kQ~�*?$_>�&0ߺi,P����d�d'�^l�Φ�4&�������Hyk��2������#ȸH�!�Ɯ�vO/�5��CF�3@��U��}@�m�@�J�>a �}���E�����	#�8{=�mw�a��A)?��1�!�.���U��(�U�������:�߆l��������N-�_A>#�0b��	� �"f�6�iX�F˲Ik]HT>)��#������c��#�zZ�)m��aył?�xg5��v�����oM34���cOx�p���;�I��Уi��
3g|�)�{^z͙Y�z!��=2X��I�m����������`�E�&�~��`�i�o�I���\Ɋd�-�fԯl<��;A+R0`����<�/(YD��Ģ��&!b-XKF�)Z�a�r+Dj� .�d� ��az����Ҍ!���B�X�WU:ڞ�`F��8�<�z�Ug�|f0gF���Kq��-5mn�s�kp	Z⤛�����3*8�h�Hfk#܇ah��FӍ�a�P>��1��ZOs{g��𒎹 ��l�jҨ�����v�Ǔ"��7�w�t�.��n6�Nk����)����O�:	����t�ڵހ�W���5�mu-�0.�	-?F���?���E�� 
Vts`���R^�l��<�n�Q��(���&������o�j����j�Ӵ������������C��|��pӘC�hM0O1"i�=s<[x������ܭ��2��j�l�����Y����HZ������_nM���F��w~�vM:w(������.E�X��:�F7���#DS��b��k��7�-�BhȠ\��=o�\�Б_r�y�}�fz�Y,�uWw�Ӂ����٧f��6��/x=@�tM�/��� ����v��y��?P�I�db���B@�2;v�C�)&���0��X�,�e�w�F!����f�X@G����g��l�4�I��#��-�9�������뼰�G�(&�����!�^V(��9�c��f��l�'\-}k�-+�W��w��Y�����Σ%��
����1J#�s>P:�~d�Ԕ�'�N��ާ�뒄�!�X��9�d�EHd��\"v�	ˎ92�va��{�=3�<��u�U�P0@�5��p�Y�N�T�]P.P�_=�,5j���M�p�	�H+�$���'��]���/J&=(�q��8j����h0McUbi��wu֍�Y����/6��b���҄nz��<���ȉ��Y<'b���/�o�J�<C⏺
�H"J�8�ȝ|CWU�E8��h�����������:I0o���9f�������i�Q��V����n4���!��S�)@��>M6xW#��Z&\�I3�u��Y��f��X;�:˒(�G��^K0- �^h�n����
��S0�m{	^�ũ��%ș�&G��k5?:���m��)���`�Qrw��*��B	U��h>�w��{<.qo�y.N�2N��;��r/!U@��/�ۦ��t�(3W+���{��6����t��K���VD@\wN��ӎ|�]hC���
x�;p8)D��3�霪nV�(��tÜT���zT���Q6�p��Y4m�"���2�D�"
8�Fo4�-�D�ҁ�B�1(C��q)'C1��7�@j<-��
�>�6ߥ�S)�E�i.)�|�sح)��
�9���w�߸�.8{��V��+b=���������q}�[�C�g=(���k�m��~���c�a%��'�X�e�<���z����ō}�Q5hM����9;�W�f
��g�ϐU/�l?�Pu�J	�c'��Ip����̔������y�*������	j��ǐv�/�L��0��%Kv�����M�'\���
��^[��q\�݈��<i������Zٛ�P��ÑD�Z��\J)�|�[���\�XM�k\l����G1�ĞK
�u��W`��
�~`����# �n��Z=Pa�o2�Ӳ8ZFS�^𼿂�L�?�P�`�Qwn�_��g�[��a^'��1�[�7tث(R,(q�!�D ��1��G����|�@ELT��!�����"~h�=.3�R���vg,��h���۩u`u��K�S�������C��	�����3���^�]I:�)�oW%5�ru"�DBFL:���l�&rd�r�v�K�jaگ�Ia]1���@�+�#g�|Яݚ,����L�Y�
�9%O�:��[Z��4�VG�ކ��Q��0�->��G=��H��#����ߑ���.��߀�pmO�?����Pl�E����OU0���M�4m�{Bt����>�R #ػ���IwܦW���w��+���S��t��'�0a����QrS>�s�\ob!��H��Hlj��E�k� %����1G�R�vd#�ū��\���aZrj��m����M�e�t,�/�:��ݞI�y���;��i�2ذD����u.w���m����2�@WY C�f�d�������O(��*G�?
zB��f���U���h����?F��lw2-��w�n�{��
�Dڇ�,q�I+�|�p�z!�)����47��Oe��Dqm?A�bE���3A�^��;�Se醓*r]9�3��m֯��>�W����٧�A�D���&+�!�����j<����D>Mw"��^���I�h{�0�Y��;3JƢ1�"4�{�l�P�Q>�$3Ib��A�z�A������U�o��	l�)�����Vļ�y硅��"�d���t{������������9��D�)J��f��P!~)������..��)��d|~4�Z���`k���\f\R����ҡ�jy�`��0�W�{�/��l����vj�e���1RӸe��A�Ŭ���ɍ8V�GR�C�"7@�A�P&�X��ҋ�u��$���C2�G0c�A֘��JgҺ�@�\���{�6!�ⴛ/K�?V��d���V"7�rW��U!�)�*#�C�g���ϝ�{@���?'�� _���Kdo;z&s�i�=�b��ʗu��A�jK��N\^��Z�1+��:����Jv78��q3xb��Ѡ���)=^V6�Z�j�M mץP�sH��v_�d���`��Ԁ�[�|m�%ssq؈�,{�8���Y����M���i�k�fc8E[UCq8<�P���8��#�a-�VU���w��}��~2�z�r.�P�u�
��.���Uo���1H:H�G����A��}ef1u��n���y�j�1�c�!n7�h^m�*����@���4�RI����ފ��VA�eT��K�\s���b+@VD�%dEI<fR���W�X��*W�����$�ި=����[��A?��
�~6R�+*�D.J����x�tx�������x&�2yoA��U^�Qlz.2o�n���r�^NУ=vr��^k5FJf	�ݼ/G���|o>��!AWQp�ׁ~����g��2���yw�*R�J*Ө>�u�>�����M&�A�>u
}�-v|2� P.v,��'�̄`���4��ݏ�
��C�2�Y�,��)�'���v��r9#���!�i-����zّ�xr��9���b3)Y^��?Cp�KE��/�'.&�|1��̽`�9�j����)CM?`, 7|3Ll�V���18%e�#�=�c�����P�7�B��Ej�� �oA�;������%�M�O��% |d1:q1�T��1��y�˃�����^�l��1C����+���ļ��Ig�z��8�F�]l+�L0���	�W�Ws���eT��c�󑞕���5��dh��?䑮x��q��w�}��g�x_�=S��$�V���F��3��B���rF�߭�%�OrT��TLu���Y�"t���C|;4:��o����G����L���ek�<J<OG�n�7���!3^FQ�es��W�o<���)5S��s?z:ͪh�y��m�Q�f��a��')�׍�PHt�dU7svN��+_����ނT�����QGK2��9(8�����5����	�r�I����_��ui��<��?o �1�^%��@�'4���"	N�����J`*����3v��*̏�-�'<e�u�t#o1�F�auD�F�j���fO=�s�G���wb�8ʊ$�ň���}�T1l�(TŘ/�L�&CTo�)�EP)��{���my^➩c��ҷ���}./�И�篢�&�E��<	U�����ipz�z��#+`{����}&U�6a�<�hi�6��&T7>\��l���=�Y�.����Y��S�{B8�gowo!SflP��A.We��c6��|Pz��;JW�x�mH�.�`t��ݜ�+Vo
�ś��oT<V��L�HlƍK7���hA�����[��9}x���ds�P�^�f �Q��B�8�(h�C�8�����qM�$����>	�2>�G\����r����w���8��q&���Em/cw�`���~��Ƴ��e {�?���O�d�\����}��u�f�#�PW��
�β+	qu����7�� a���o1D���%�x�mM�������9�:*Xg[!���dE���=�,�*�+��@�������Mp\xO:�̬z�Vv�a�-���3�r�2Jޠ���d����0�L�1NI�]�4@"�JH+���Dm�ʊ����K���z���1hkՈ��jyՕ��4��5�y\���D=�;���AM�2��:��u����z��F����bB��!��tӿZd4��d���pP��d�LD���2���Oy��e�nb��s]����_��3:��}kU�7�5M��ϥ|b��+O��]0^�֔OE�1�����i���5 �gƎ��$}	��E1��� �C�fs�h���]�OUm��=S���q�%+�IE�%X`Ln]q/.)0�fl`lg)��AU�W�T`o���;�зg˔#��x� �[b>�ݒ�f<*"�;ȼZ��1D98L^[fht�#T�eg�յh�,:!Aj��A�L���3{�4���,Q}�F*D�������yA�bp���=h��ҥ}y!���3W��	��&ă�݇j��ݷtM���3K\��D�r��{1m���g?\���DӠ��;4��6p�\bJ�	N{j)E��0�,��0�b��||��]t��g��|\�m�����Z�`�S��M���m�W���Nx-�Vv��Q�=R��mh��Q�zJ�oNaU^!?��ՓQ4��#����L����2#BC�U6ǉH&=*9�?]��f���B�^Nh�d�P4�V�m��zKBk |=(���}{��X�6����\E�v֏�۹�k%q�SERT"!�S��Q���U���� �X<����9ɥ]��^(��䛿$_�u�au��J�1\�J���"t��a+[knW8ώ�Ά;W$�\�Օ���'���ߣ��t�z�M!�qCX�8~��������x���d�JE��@8�o�ZM��l���y�g�l�`	���D�ID!m!�v[vAC�ft��F�S��� �$���7��2����5
�>[{�5hk�H,�c�m��0&O�k�����umU��?�U����>�l&����:t��P2}�a[�r�&��#[u�6�k�i9�ƈ�Q{��阧*^��'`MTR�w�'�]B��I��8�8�Lm �����,�8���(h�]|�0@'�!�9�ƥ(��襸'Wf *�v�>�+LV=�6a{�u0$?��yo���8-�r&���9��KQo%����<�$�HLo-�@Q��A.(2M��a�o)�� �E@�\:�!�>�I��5�}�8����u�+�iO�$�)�:s�m�f���W�p�������0r���]�nu�-�e����	����ù�[����-���_m���_5Í�ǵW(q�lk���/��o�VWp�tPl{�3�+�"p��寴��
-;�Z��$i�6$Y�>r.�hB���A��A �������?��d���|�`+��I�Щ�>K�HZTV��:��Q��� *ʁ�r+T~�.T%���=٫�∠���g��-�nR�	+[�#=� ��"摖֮U�����DL��8�U�P��vU����ĕ8�}����d��bDR�l0ϻ�nW��F6�R8NP�j�#s�Y�=����W� �E�}�����*Y&�M%B4Z���`m'�5U��m�@DP*Mp'���
������O|�X�7��,*q���k��|��ȧ]B���t�����vZ�$v��������%�"���Ё����i�P��I����v��O�'�L.��53��$�to*!�ꎸ�v��u����z�5�0�,G��fz*�5���~�:�籒L{Gv���+YN�.�����ۃ4Aۍ
��6�T��؉@9D$\���Z%��r��?�Avp�)�Q�o���~�SeS�XF��6�7ֺ�����5Y�v�F��S�򗩭��R~��	^���U�(��SK��(ᙘh0?7R��
�)9p+�:��B����_>�޵!K���n-��A�!�V��KD�yT��#P�*��E��3�B��Ж����?-H�v��Nt�A cu~g�hN=��r�n�'R��L� q@R ~���hwRP�n��\u1��ˮ4oӓ��3�cH枞�L��{Pf	���J�IN��R7�q�����Kv��:�\�#�G�4t�c�K��S~}'�K%�C�Ȫ�k�UKɱ�J�Ia)s������YiF;��g��ݳs��ߛ�C9E���Bo!�S�!�t'se��	��"´��#{��E��J�L뼎ϱD��CO�֋W�G��+�s[&��;t�9����D�j���+�u�Y�	#U�3�,&0�Cu��|Ʋ�'�r��M��I.|1M�W����`�u��Y\�:ke%�ѡm�g�f=o�zʯ�M���2l�V]
s��ww$�0$&{kC>����1;S����V x���U�Z��
�t���eB�������n�&���u+4��*ܿ<sp��7��SX�ml`�� �͛��}~j�(z~d�I�L\��P� &�@g����B٪cýƻ�� j��ar?�����dy}�����ߝ47�j.6���m��84Dm��1]�z(.x��A��0�2 �g. �x��n�==���q���o�]�q��lWt'�+�b�����i}�z()z����̙ip%S�Uh�TQ�̓-ʖ���"A܈��d�O�pN�X��}Yr���`��*�YG0�zuǫ�����at�Yl;9�Co�5_��~m!�a&5������IxŲ�*�)|�bլ.I��6��G��|U`Y�-	�av�gbt���n�~�0?-�k�ŚI��!j��6*��C�6��ʺ;��K���=>0M�G�.��3�C����Qx�4�-��̪7�$+e'�q����q,����@��Ң��s������usV踇�W�c@[��L@��긍?N�.�~=zh/HJ�9/��>�5V����/_�~,� s�O����"wx�ϥk�o��.ŗ�&k����
��};?JR�)k�8��hɀ38�ڑ,����9�ToZ��y$}������9��Q݇�P������*PF�J�KC0�qZl�'���D8`{�3�C�NR���l���n{5����\�o�Hyt���ǵ���p"��v?�$c�_��0����*�m-���W�f�_�RaL�-/wkY	����F����[�*����5��1Ƣ�l"ΥZ���r:j����=����ߗV[g/���n%̇{w���,�ϣS&uGŸ��+��n��H{�� M��~��g�>+�^!�L=�4�X�@�� ����Aizx�4����`�g4�V����JM��η�E���U��r��ֽ;hZih���h��L�q��U�e�u	�%?��T�dc�*����Ӎ�D�siJ����V\|��b9���	q���/�ß��&hX�/�'DP� ���������k;. ����Ic۴pY���Q�>���;w��>\|���2���-�ff5��������W��mU!7�B�����jc��d���k9�;��=-�x�������f���o`��M[���Z����"���l~�逽Չ j��В>�G�IN]��{x�C �I�Wn\�`��o96�F���a�����Ɔ��~����0�>��LRRo��	�|&BB�޺� �<A�`\z���&�sZ��&`��o`I�b%�|�
4��fL�Z{���v�g���M
�ꜵJ�*l�w ��e���-�*���XN��k?9�*f��nj� |�]~!+0K�=��������TX�C�q*2���ǽ�~vح�ЖnH�3����
\��ı�rRa��բ�X	���sq��J�ʄA�U#E��.����g�9�;�2���5�f�$i�^/��B|���u�`\�{�D�oF�l`�j��z�_msu��!�7�8 �
�K0����������n�.�w��h�S���c��1-d�=���&V)�-�u[k�1`�:�tĸ��n�5S���T���d��D%�V�cY��	D���9���f�h��Ü�!WI��.�P������Iw�e���w�+������TQ����q����;|�w����%T#�J�x����}�0�V��gO�3��S@iMgS������`S��f����
��R:<e8� ��1�~�Z��n�5լ%^�������R�EO��G�TF���
��"�-Yt�<�}���?����]��:��C
�&��!dh���s}!Dw�e��{t*/�jT8�,g1M�Do�R��!h������O�8|?\8q0!���G	�����`�Ȅ�(&����K9���%6;g5[�^�Ck\b�$H�	�7l�aSc������x[�BP8(d�)YA���nv��q��ҏ�F���W9q�s3�d�Фa�F8,`oG�_��d�k���*Q�u�"oH47E�|7���ˍlYH���T�@�t\o�����l(�R��a5E$���A�!@�c�T3F΋[ֱ}�2�x,D<�-�-5m$������D�.,�٨#��u��IU!��Y�>��̱U��R���F�j��}��7˝Q@��87�t=��%�hW쑨)��E��� �٢&!L�J�Ř^&������B����� 4��]]���C�����'���aX!�F�q� )X��>���݈.�-L�K*JT5���;%^�<���>|5��&�y������?���"{{Y�ڧ*�&��J�kY�����c-X<�
��|�e_BS��ڑd硜�dNy�kv������8���w�*|�9F�M����{�\��i�,M��؏�]����s����O��^�?��s0+��h��4����k��!���쀟'ŧ8;�^�ϸW7�'/ *� 6s��w���]fߦ�s�@�)��;����XQ#�͂i���+bȧD�����q�$�E����<Ȑ`x���4��DJ;vxE{���i֕.�x���bW����'��=�i��]��~~�,Q7�i��%�5d�7���_�{;$[���o7��7��Cx�&�8Α���J7��L�
$����N�m&
�RûEw߃�ݳh���c�V@'��z em���VL�x�ta�0���~-5(1=�q?�
u������J$�� } �Բ�����'q͓�=`��U,�r�}�_.�u��=�նK]0^�k����v,�kY���"Y{Q�,L��Vw%��VcHI1n���@����n*I?�\����/��>�2��륅�4��<�82�<���!�Q5�7�C{a�
#e$�uY&wu��`�2�����'�_�)H�e}�J���gx*oi_�m�w*�7�˸X��y�maa��&1����	���!�ڶ�.�!�n� �\��D�oMK�ۗ�$;U
�/3w�ǧd2��ƃP�e�O���a~�֑WOD5�l,`�����<��<F�HU��Y`?J�0I��Q��� ���S�׼�#��r�ߕ�<-���_��$u�!Pޖ�pp׿U�,��џxcHT_�� >aQ.�9�D�I�j��>o�.Y5NĤ~��@�/���7�+�^MI����O#y
����mjӨ��'Y��\�IdL��3�$3��.ͼH Ӫ�O�͢w�CN�q�Y\fpH^W]�`�s�.؈�Q�~�zv��V��K)z)���wj�x1�J*���CO�t�>��(>�d^��C�YM�/B�֎k�c�H��	��:+�_Y"�2�-�R'�s#l���}ŷ�F�l/n~&"$�=�F�� [��+���bi��{V簖3y��&XV���J�J1�_K��� �?T!�t���I�*���md�
4?r�S��Kta*;���Cy~�1:�T}�M���/��"K=��a�O��z���X�u%{�\�o���S�b��J��t��]H)�ƞ�ȄsF}�B��v�+��LK@�c��ߤ��+݊�r��BqdJ((D�����x���̊Yv>H%�k4268�55���\�J|��i4�����P@b��(��Q��,�7L��@j���q����/���(�t7�ِȰF�y����qh\�;߮r��a��2��v�L�ם�ah�c; ��8]Մ���ᚷ��ϣCug�ά�h!T���&�����B�!�	D�q�*�-վ��r����I��b��r@�hԾ����4ր�8JWfJv5'��eW��^��b|��*�ٔ�|˴�
r�b�)�e�vly�e og��.��τ_�3�O�í1F�9���΋�5�Ꞑ%�1����^��֎s�H(�F�裩 �&���"�S��+���l�H}w��}�J8��;�.����E.1,AG��w�=�����n�&Y���Z���O3u�IC�.~"S�G�ګ���S&1rѿl�A��P|o�7U=�*q/{|',�?�1��B����R��e��6�, w<>@:h�YD?D��W�����p4>��D6V�.g��J������j�R�>�[��z�J:s�l�Jb㋘>X�,$�ڤ]���kpޕj����U�6�_��2��j��/H��\�Շ�1�C
kH7P��FIZ<�~���Cp�Qn_o?��s*i{I>e5���7��t���7 ��n|l�p�qY'���Z����:95���q������αw�Վ~��e��	��3��l}��o�Oр�nS̳w7���^�f�2�èM�Q�D
�MP�����J3�7��e��K���K1�<Eb=J˗?Md��P�h�foV�-����%�؞d��n39�j�k�`�O���^�;@�A�]p�)ȔO���}��t\-Mn�VT*�-{KN��' W�%w�ߗ
�{#f�O��6[�k���h< EG
�������{��ع�5�"rI�FP�HkRr[ʢ��8<�3G�V�[L��~��ND�sD���E�I�^�աۼ���%+|c��:o̮8`�Ը�=k[��oZ��֚%,���Zov�v���t/�q3梤{D\�n\L�h����Wt:v�x�$���;��Y;!P�P�J�
k���Mo�L�iE��9r�)jw�b��jMW����Ж�Y�j��rP/�]D}�֘��k����⡓��|������L��A,.v[���,�nz� �h`J��`ifQVȨ�؜�롮d�t>72�4͸��I���4��U���3W%��G�D'���l��������9r�}	�u6L�I��V�/�^؎ C���?�v�x=�̂S����T62���΂���l�l��A��טaO���4���X
�|I��Z�Z��-c�WT}|�(ĭPH�=޻�z����:���>1I4.k�L�{�6َ���8������ �G�v�c�@�lg���4���z�(��e�Z�'�9�e��J��J�^���=HΨ=��x1\.7���X�68���J���4��ȩ���N��;NGܠ��w��P�V� �t��cgj��SJh�ñ�����W��>�/n�0�"����i@e}Ŧ�җ����7g���Jpp]0&�a~�&ԡ%�I ���?1��H��ǁ1��ǻ��H^{4�@��2r��P&�����+���`��M�(|�^���F���7����A��c������E_tlz,׶�8��B�~%��7N��_��l߆�uͫhY���r��6ԥ��"�̅`/�!�i���aU�yӭޛ�	I̗��D=(�uL{�>'m�3��/rF�e��8����B$?ZJ�@�?���KȒ9���RK +M���wX�1h�F�������V��n�IY��\"���6v�B�kټJ��U2��
8\�#�~ģbv	~�X��x�M@��[����I�_b΅�D��IR6ݴ���h]�`$�H�v?s�Hi�U��6|pIo���{��x�Dgw���1yɟ�|9��aF
���cZMA)7��Y��@"<7�J������K�5�0� R�J�mv�Dm�BX�0���s�ٜ��4V�`�eP ��i���R̭G��ںW��p��8@��u�RyfT���/W��� tX ��Ѫwx���E�14A��X�lJ68�P��
������[��˖53�ׯFn�Pe\����Q��+5BX~]�zףEj9s�õ��j��kN�re�J�@nl������6��S<ܐV��jWE�QP�
Er6>��}�FX?y���⁸þ}Kt���f^;:?�5����~p̋���?Bd�E�f/�0<�z�s��v�ʶ��O��yM�P��L�hE��~�[jȀ��ɸ�m�W/�}��ge� ���Fǽ:}̅i�)�:?�L�J)=�f����bϷ$ /$�X-�j�ׇ�f��on�TBX'�R�U ����:���J��s��&X��仰5WME��P�>��v�WBT�v�V���~կ�"��Rbf���|��@�
��A�����/0<���<�$ux)���i�T�z�r^�R�cG����?�.ᒲ��j��:��G�Yšnj�W8���}7
{��e��7�و�S�K�+'ehiё��BÍ�����<��@m�ii�[���wSm��y��aqp���n��$g�t�������dz�\����Ռ���\�=�ɀP-��*:
)U�0|�o�E��ZH ��l�ސ�x��|2�h��ӄ���D-��e��Vܥh`g��hgB���8�賓�£�����Xz��۽~���T��>�!�Hz��չ�ƀ.z�/�}�w����!<�s k����r~q��FMag�?\)�D�P�H�i�牮4r>�3����S>�K��
/@��"�v»���S���8���͵��9���!�2<WJ��tv���D�f+隁Ӆ�|����a���t�X\�x�&w�J�q��&#���8��~"�j�S�N{��B,w���#��8;��22��n��UJ�|��@��ƅ>����4bkn?ޙv*z���0lF�0�o��y^b����o�(��������`f�s� 0�ۣ����O�Do)�,�A�H���M�%��Up�ܑ�����5�vr<|w�B���ɛ[�����Z�Q�6˄f.��� �#���
�'�.�)�W���j�o�H1����J��L��pf$
�v=�$-d�|�a2�;Z ��H�/�Bf�Mc�|���,���kJ�����GX�B'��K�f�x��#�e��*s��_���ᙻń��,�[���0�gY�jGW�'Z���sԑ����	�
�׷*B��M��g&��h�䉅R��t�.m��6c�ܤ�f�|
{+�
�g:�l_3�(x!)���*��!�gr(ܱR���v������a�W�{����D�}�\��P��9U�_|��
¢�AZ96�LA�#V��=d��ϲ�u��,�MBb�P�/T8m>6g���7_�wb�/��p۝d�����R��q��Xr�ʋ*���ʹ�C�5�>c>�lxo�G���j�?�~�~R��üFTnK�@��捁��a�ˬ*����cG1��æ���b�|�M+��Y���o���A�xcH>�R�wr��ó��ɧ���B��d_��Gg��Q���m�mA���W�������!q���)�#Iw��4�~L���m{wU.��<=b����tl#%Bn�ΐ�6�J� �̬d�=
�s%jOS��1���͚��A��L��ح�[xy!�2� λ�#�S]�}[KݘHL�.�
d�k�V8�o�.�R~��9��]{ڣ��D����P ��q�\y�&�P��b|JSBd+�)�@��IZyP��"���k�w�Hf3Z�<J����]�<�q$��TTLĶ~J��$we��y
Aj��	�9h�? ���v��:DԮr����:��6���{�$��'�oZ6�\��l,p��Y�h��)Үgo�_5/l07{LF��#�$���-g����߃����U��ÍJ����#�a�:����u�u�/�T�KI��^�V�#N�J�y��Ev5I��hU��X����Ѩ�t�H?��=Qdܛ���ƒ��\ӓ�I|0h�k�Uum	���}�1�p���f�=��h�<�I�.}��bk���FN,��KC<������6�λ��{���e2e�,�F�R�u[B����pG�k5�6ZY�5w"+�Ov��J!ύ�:z.ޱ��e[d6ڊ˿�E� �����_,Kٮ]Y��(D��T�h�eN��q�)��kϛ��++�Z�d��w���T=툈�.H9]��zn������J�[����C���y�x;"��o*��S���������ɟh��hG[�$m��sh���d��GC�4���G`" �V>�	|͔��ʯ���O���6�W�V�[n�S���!u��"5dJX��еB�Ǜ]A&[7�6�������!!V�!���i�������U#v�e"���?t���o��@��>�W�gl4V����A����n���e����y-$Ԛ܂Ԉ[k�?�[�L�S�q.����@!�_�r�@�����0����M�CGx ��|��W���������ɨ���B(I6�Tk<D%�.hyHTC���D���RBl�{Lb8k��@��h�%��blhp�p�tFzDOZ۬H�!Bk�3�6q�� ��IZ�}b��i������?�7���۳�����.��X2|�E��۴��W��2n�¹,�G(ݷ{Std)_n�� j����9�f�c�o��N�Ż~YƮ��=>��Ť��6k������hzYŋ��o���s�A������W�Ca�\Y�}:3�3	��ŝ���z���� �F+C��뼮wT��X\��=^le�W^�T�!]��+�JePg��MS�׆
 xR������!�����^�n�m���5�s��d��f cvm��Fr�0��Ac���"���b�Q7�U��٪�?ɸt�^�xTb_Z>��Tѧ�%����j���Q���|�U�#UL�ǌ��i�E/+ٝ�:�X1��"�~��\�_�`�����{��׵�ڑ�ľ����h����X�u/~7�B���)u=���sGj��f霟���T���wB�o��K��=gGɋ�Ъ��!C��3���Z�յ�XH��I�K8�>�����~�R�J��xJ�[n4{�/�2ᶋS�4}Ź����^�&�K9�k�_J��+� 1	�/,"�;�),f��Hj�ӃBR���@��C�N�W�6s�t�~�w�$�����9J�-���������Y0di���
]�����lsS�2yyr����a�zA_H��Q�@�6��Z��*O�6��K0y��,�G&v�T�^�Et_x�( ��ՐQ\2�D���y~Q�eI���ϴ2���
���J��w�e��aj����FjsVL`j�rRG���p�V�8�ʹ���W��7�PM����!k9M9S5�-#FE�|�s_����ˈ�˶.�<P3Z5乛�_l�'߷�`�j�˅g���/8�� 7�����9�P��i�3⪫51�z'��n��l#��h�R�c[��\3��}�w��6S �H��+5�
�7Ga]V�o��������=��&�m5���_��
m)�N��D���Zj�5�R�m��\6���!�nIȒV���Τv�o�6���1��,5��%�Eg���{������m��u2�R����;k�	��fR��z��٩��Z��Bk���I�-��7�*Rt����\!�A���Bک������v����y#�`Λ��_1��u��sD�2�h8G\@k�໸���F�~5.���A�Ve,$o��r���t���5䧮�)W�4���/���������i�ε��>�A�����o'��T6�Z��Hd�0:C U�(2~�P��[ ��$!�):���TM���0�l�o�AmZ�O�ׂ����1�Un�,iqA��T���z�� �{�L���!+�A�{ �^,s%�3}č�l���� �\�#�dNdRYܜ��7����<)Uz�����2H�=�xy����T�>�ٚ�f���B[�}��ID1�� z�)���,��JQc[s�w/fn�V�p��\����l:MT��g��Q߸98���.2GR��"E�-�-$]'Ѓ\gNƆ��j���ٙ�H�b�h?RO�M�!�5�-�^!3��29O�4H)�2��&��|��K�{^�S,�����4f�y���~��)elB������I��"6�=W��7C�Y�6hXw�n�����������=�h�6�"<��c��uD��G?8�l3���a�Q9t�f�,����V�E(���\���]	�8Z�����0ڐ��傊,�=�1?���uf.���v��&�xg���f(M���|UH��R�{�h[1{�������"icx��vY���=�ɮ[� 6��% �f�Aoƿ)X�7��Y�!�����Ю�º��]���_5�6| �Y���e3�A��t8(���:$t	��aQ��e���ٹ��r�y��_�s*�QI��Хh#_F����fIO�*��5F�X��j�~�v�u���Y�.cQY�|����j��7�+3&�i�*i�m�LR��0�����G�R3����bf��|��
{�z�����1��E�T���F���tRs`�jǠn�X;(�d��2����.�A����&�Z��BJv��a���PM����Ʌ��Jg����i�1����%����Ol�{��₊>�c'3�^�|�h"�G�7r|O�	:͵r�����g O��\8�1G�z��}�W^�d~��{�c�z���K�˸K;��������.o�P��޷#�X_$ ;\�Ż�'2U��>�R�G+�8�);)b q�_���/~�c w���0�v8�QLLB�N1��8]Z�7F�WV�z�����$t��)�R��@�=y��F���_��c���FC�e�s��5���o�R��	�����nJ�����4�md�(��i�c�ҥkGM��t`���&w��{��}]�Q�!B�!�gk?\p	�R&~�,6�z�V�2hTT���RCP����7R�Fܿ��1�����j�W�
�6i�z��k�IW=H�4��(��jĻ����	p���{	��ڐ�����P�*d�o|rU���8mӪ88����%S��e����m4D��z ��M"*쀶�@-fW;B�%����$�EF�<J�$��A=�{��3*1��S��<2�j�s�d��( ,B:y�JO��X=��	�z8��ڻ�D��^ȖE��{w����(-�T|T�(Oj�߲�	4�!Oql�KH鉉�FǏǔ�u��^f�󒟨����n@e��M�fcB���,��{ޏMԱژ�0B��[��h�q�G��d�"z/5}�2j-�+�9�^��VC�x��n"m��6�ϐd��R/o3z�ZR�4ma��7�~c��f�(J�;_��e���Xs��	�9%��8�rFQ=��p_������w�՘:�KB���ICr���5a�@�'&����#5���+����9�␻��0�zf��"���5U�fV�"�&!?��s����N�G;�3h��Ϛh���o�I�!�ݵX~�$��M|�$�-�8����"�?QJ�k!�m�������76ֲ��_���?W�5a�%�B��'%Ek���
������U �����^�B��(���g�+�~c|�M��X�,79%���5���N�����̂�ӧ�On��"�ڽ�Z�S�ec�[�g��wkRKJ��S`+���S�e_v�t�h���� �+�K��Y��BEbԳA%�ZuQ�t�-"}�#��j	����F�"'��6�����6F
Y�\|�ұ�l��0
�O��B�M�'�B4W|Ă�|"��	Ly�XS�>�I�j}_q:]G�L��f$�Q2���H��#���j
;�7��6#u���Y�ɡWL=���sD>'���Ñ��; �K�J� ����n	���t��J�˵Mt��F;*�������Ȃ���gI�<�����D\�bt��%�V�i�Yi��V��=^2_�\������Zgܯu4���V��y�ݒ��G�t�9�����T�g�H��x��*ݵ\Oq+�0��@��
��<�˼��Q72����A�K�k-��@#���s����0�ű�Y�߶��!	b��҇*?3��M%���f��*�t����~�����8˯3F��(�4�'�&�5�t�{��.~ QSM8�S��AJ��[�JbM�DD�*�[ٵ�+3?���
�*�tp&@+��I|�q�ߛWd#C�y]2@#�eW���%�I�9��p�/��9���-B�J@.E�=�j\;������l��>���f���t%9R����f���$�_ l�b�G���q	�f�¸ŬA���dl֩M��|�y��~�b*�P��>�w���X���h"���xX
��d-N������>�w�d�?�e���W�U\��k�$w�d�����b����j���Jw�xw��E*�\;�ČotXE��I�5�}>|�;���q;�e�\�+�w���c�FY�?������)q�"A�VR*R��q�������l����Y��d0�����ó�i�θ��('���k����'&�cfv"�Ɣ8����J{��P�c��;8$�^���7	��7(�N4$G�[���u��p��/k'pe"�F�Y�����9�g��!?�����?�qٰ�v����&?�n'�����G�q�[�7�p�|�^���Ap�A�@�F�x[��+m/p!�/n����.g7z9�薉ҌJ<�Si	C��R���7qOt2f��i� ,V��<��x�QWJg鐀�����쨧��!��Xp$D���ףZ�~���x;��Z5�J�����P�oR/%>��޿�7)� a�xki#�c>���E�g�6���F)�+��s���QD��:�0�:�N�4K�Y5
��K�ۄa��]��G*�� �%a�`Bj��w���񼳩MQ^�YO�`�-�J���?'P��yw�`�jI�T箎��;�f�r1�D���3���]'�3�ZMo�tTn.y�l��2���5�{�� �-آ�!��1Vȿ��|\����k 6��Z�䀭h���&D�E�":�dsw�o�����C��������H�A]"d0�y�t	�՝���G��;�7�UJ��{�s{@�l~�i���P7X�$Г&��gИ{�v��H$4��[��2�H��X`!{���~��q��|0'����/��@6|����86C
!���F�2M�`i��J��]4�'��{���O���6/��5y�!-�=@�^�A����-;�I����_%kެ�����1n�LA	��&�:-3�����[� �x!ZN˻^J�
�~X�ږ�^,�N��eF�n�/¡]�ʩ�=%����D	��VZkG[9��8`Gx^�ZE�A��9e�!�_x��ҐTE���u{۲��ї2-Y��s�ϑPʃ�\f�nTԱE$�Ϲ  ���m�
��lVHu��B�xpGo+=�Z�
��b8��ɴs�O��\�o�����7Pp-��'r�έ���־����zQ�������8V�h�Ċ8���j0kv{ &�����3 G�_Z ����B����J%OdvD9��CE(�D�π�����x�:��m��`)ސz ��V-��!��b/AFh��;��E��	s�uE�Z��ʏ��ܴ.7|��˖��J��"o���r�M*-_�
x����[��`H�YK�O�맧ʶZUt��N�ú�ey��b)�q�rcI����6 h1� �.�c}�h��h���S(r$��ű�<n ���_��~W��v���Tf&m(��ı��P�KV݈��^��W�*"ռO�X���ו&`��sce|/׬^S�����H���Z��c��c�qڑ�~7J!L6��?�t��|�����S�H#�*U[�7d���͞��7���C����C���&�2Q
P{d V�B~{u\6���i�&����~DD$�5��G!5����;��-l���JѦ��rƧ_w�`�
�p���3>��X9�!�ٚfZϳ�F:�@W���ڦq�AO
��`;cwU��s��޴ "f�x^�fq�o8��^�2NG����
�W�����B�Kubd�xeS�f����&���P*�R��&��b��ҢG��MhJ��9��� �5 /8��zL�8+ܶyf�䂱�PO�]�t�>;=)s.��lGEm6b�QӶ�g�U+��u��}���Q�o��Qh)��X;\���� �����Z�h��������e��i'q`\�u7�6�Ia���)�t�A��������J���1y�Tc�˚r�^b8^�r�;���Q�s�5�?u��K�.+u��[�2k2Q	�F��	��/���l�V{������ bX�oe��9��Dy�M��$Z��F"di����.��{تj��. hC蠹Tm��O�����W�Ae������x�Ǥ��4B���lP^]H�uM+Y- ��;L��9���Ǐ�P�?��:������6Q�q�	���f�q|$��e:��1���d�F+ceJ��J�4��me���b	�Ug��>�y�p��b���.��_}L#{�F[c�"��o��%�v9��P��a�c����ד��v
���r����Ӆ0���%��guu�J�<�vae�ޭ�건�ʳn�2�A��������U���2睫DC6�����㜋��l4����y����I�����[:��Ff�cY�������O��RU���W�;��N傞���z��c"�a$�Z�]R�l9sP.��!�v��>7��at����5�YƖ�6�'= ��Q��Y�A�`�k��i|g��|��o�t����/3&�v�:g)��&��o�VԄ�8]W�����3��	5W��L�� �:�km�47nJ ���"��b� ��#t@X�k��$m/A���kf1��YP6�
$�WE?wg�)�q9X���){����t����� �nĩ	���&��J�^å���?\<��f����F��'�o7g��y�:��E-���v��βUdɿ*z��Q-� E_�9��JB���h�'��Ru5=)��\�Rr0�\Fn��;ZQ$�䔵P�
���[j�~_�i�����-�%S��z�'!6��%!0}��{�F^Ն"��_L���+U�� �:��p���ߊ%��f�Jj�Dn楕G{r41ڟ�7�+Ѧ�B��a���S����:m-�}X*W�]�����84S��V��>�0��t��E�>�V��$"�	��3+	�UD�>�)��ůٓҹцK#H��$��F��p߈��F�y!�u��1�����2�ZAJ��3���̬E��I��Jr�#^�Ą�sVs��m���vAC�������0� �������q�{�=&���ca
��~E���Ma������O�� �F��"c}�Y�=�J��V�0~�b�����o� &�{Cw����?B��dx_���;��щ�𖺻+/�Ղ�0�j�������:�ϒ���ދa�8)<�G��z	�i�&7�A�9�s�ջ}���u��񖑷�8�*�WȖn���C�ᰉ���yF+�r�&�]M�Y��~�j���Ԕ������.��cŉvqoqQ3��5;�y�7w��"���헡�7RC�/X��u�x�9�NS��\���M9�d��ة~{��lP���>�B�B��~%o�y���2���ǲ[����A~RWT�}�I�*�m+g��0�i���p!Ќ�����.�t��]�i�z�A�twoL�{M؞=���t?$�D�a��{P�'������+w>=\L��L��%x�������]���*;��f�5?��( E���;M� �hB_1�P��&<���I�H��J6Ev�ٹtg��g*q����A�x&x�?:5No0
w�]peP�{}+�Yz��PFԏ���� M�|S������:���qC1�{B�?��$g��m�<>�ps�WD��bj�!��~���_��ǁHǸ7"���Ac��w{��^[�m_s��JǤ�U��3�e�&M�P�[P�v�J~��8-H�eW��_[~�>���L]|e���g����<[x(�60�a�O(�_ AP�wq�Vo��`�V����,V�H� �3��T==\G2���"�ʁ!�.uB����(��9W�{�x%��炱A���k1ʳ9k�O�`��A�S�#�k��es��:��8��6�Q����7>j���`k���[흸���2!*������=y�()[7yp
Yr��[�/��-�H�l�L�����n,3dZPDt1�`�n��I�gX�]�zgQ ��z!m�*�S}I)i%��9�染x2��p8�93�������\Dnc�x�ň���:F��!�`s7/Q��)���P;���mjD�HЄ
LI�<,�(XE�6^�*����$-l���\�K(kә�_|q�{3�#����y�?j��-�럙���%��������BA o�*E"�/2��)���uK��9�;���ťiE]���|�z,���!Ӏ��f�L4���Jqv��=��GU�H�!�oP����k�+ʌ���<�T���x
��J!��pً���4��E$Y����|q�e�*�v�;ov��O^04�x��K�B|9n �Q�p�@�_���̻�O��f��3�m.����A���/N�Z�j�p�D�DX���V�W(M1�D|���._�(vB����w�ECV��t�����{���e�B����m���瘴��hm9iuE��s�smmj�1G,�����hn��a�)e ����J@292*?�8��!��$+�;����Y=�~:xo��C��l�atA1����[��n�&xk���h�.��a�V��N�a·`E�@����(e+D����7���A`r�}����K�yeT�������&����@��Ϝ.Z1� 1�������*Rk�y��qAڰ�Ǽ9��7��P�r`�ŚM�O�򈺞qE�/�{����}���;hܝ�����co9(�b�VcK�R�?2��TBg|�?�P�s�
�*�\���'�6�:
�GY�_ �I�N�2� .wz��xc�p����;�����,/8�U3ɳ�P������"�ch����I᧜~�7���H���l�;W�6B� kce�t��_؋�(�W��.n|��(F��J��.�a��90�)N��#�~t(��D����8F�/F#����&Q�y�S����!S�p�V����ը�<�l�C}��&�����d(������}��F� Y����} ���I����q����䷺M<`��]^�4~SϞWc�qH��
�����ڝ�����M�PD�N�Y��#�x�����~6q{D����i�jH��(��&$K� �� ��Iټn�zR�r�T�[4���۷�v�|Ҋq<�@���/nY�=��^��%�و��p?������w}�Ʀq5f"}�)��F�G��ޮ��H�hd�VG-΂Zs���\���Z�c����˽��G�����&��\�X C �U3�jv|8W�)��X�M�D�"%.��a^��k�u��EbI���{� ?���E�X٣,���:r��{֪tF���@(�h��Z�� V����\�Bz�H5֚����h�F��|r;��)��r���N�2�ģ�����t�@����K�#X�.��k&u_JX�X�S��J�slA��֕�i��.��
�\S�1��-�6�ǀ�ڑT��(�����_U�l��j��Pq9oss���2&W��GG����:&v�d�I8�x<�|��,xtt�j w�Hk����x��$0��w
ҟP�K`I~�xC�Z�4� �3�=�ِhg��`�ҩ h\u������*��`|�|f�M�Ƶ��V]I���Y��"�?P��T9oٞ�
}��D"��e,�ƅa�*���?��Nη�+�d�Qݎ���f�F[G����b�r� ��\���C���icOY�d*ҕ�����7��\1�Tn}^Aen�h2g�'^�D��Ϻ��m6Z܉�+5x�>5�c*�B5�Ҍ}-?9<s�ZfJ��L��ܝ��Z�oz�; Zڑ���w��Ѡ�"x���=`=FR���?������H�D"=��4��.�����#�[�G?�dR��W�'�ę����k �to����ʀ�a��	�}�m�2z���Rd��-�$Y��P�Z���mKɴ������Ϡ,X̯�gϓlFbo��w�g�(�B&��f��($�5���u$�PC����ϣZ�K�nD�~�?�fR0� V�oq���q�3��%���#5cs��F�خ��kD��U�3^�q��'8�+,��Z�`��W)�o��]y���ߞϚT	�zY-&��5���1�����H��)����~�	���S����2�%���c)��z����a��4б(��٣P�_��|��1��D���D�V� ��m(52��'\9���p�9��~�Gy�C���/��DE~�Q�I��~��D�h-Wh�yv����=d�;��y�*Jf~���t .|i�{��\#�R&��A���>ÿO��1bv+����6������'Z�Z�� '�9~�"ԯ團�)����������I�<0H�Ɛ!ֺх1����MTf�/n�EG�]�����>��-!�m���T[Ql����g�X���3
75^��U���?�x�b�2OO6���o�:ިc�딦:�}H��AK� $�%Z>(���B���F���	Q�%�M�1�?f$�G�(DmfǇ��R`�
q�s1�r����������c�1'S��h[�z�w�Q�m<߬��zaj-N�{�{U�;`l�;U��x��{qg|`&m��L�V�2����)��p����7�B�J��oZ
eA�@5w�1T���M���4��]D{'��B�}ʹD�]qC�a=pVl�g��T�|���Qp#\��|��8��m��$7��>�V����74�!I��UN8	8����.FE�}�Μ�#��>!ora��u=&x�`]�k�q���>���3룂7g�n�l]>�a�fr��R*��0Q[{�]���@��-��)7�܃6
g�1��2a���)6��Z��M��:�8�Ӽ	�ݰQ�;�Zl:uLT
K����玒��t|�Bҋ��F-�\Z�������l0�̱^���BV�0��cVT3�ەu�����w�)�'����W�	$�g�9x���h��4��=C��b��rA�;Ԇj��~���>B�H>��es�M�+�dkU��TC-n�;�~����޴��
��Fg��b5��>w���ha�'a)³?͇�,���4��'��N�(*uNQn�*��t�Qr�cT7U�K���U�1��U���r�&�J"����F�7�?�<DP�ŷ�}z1i�*і�3Y�5*Pd�� "}�ܕڑX��.|A�$w�V��"��+?6f,A�'���)N%�^\<�yjf_J�E�_�P��I�ϥ�:��|w���f��%v:�|������RE�*W*�����hEq�g��l�܏#�L��M���WE���}�4����[27c S��`�����?w���ň��pζr�2����V3�n�v 5k6��Yv�6��iܱ����!<w�Bpt�SW�+aAL�@��~?!B
Fl@^(HU�p�0� ��"�+E],�c��p
���RW[�8���S��t�s$u,�Hew�c6D׍�a�Y÷�-��۩��X�ۖ֨o�jO�`��Fi�D��V ��wV�D_oʰ����"g!�%_�%���nv3I�?��߁g�8��Xk�)��3�sAFs���>�r7��P��h>���1^����X�H�	��ܰG�23\����l�¶*SE������L\�s�	���N�	ڄ�;d���R�u�t���;��7
���~�v�����M���$J���F�D+~�<��]F�\��@'?uvEU9���,�mW�@�7G���8ӵ�����^0��|�?�ހ3���vo�#˴8 ����%s
Zj1c(顮��x'ޭ�|7a㡪=vX�ray�-�(�pGr�,���9.���P/��h�Y�4�l�"2��ʚ1��4��ݞ�̸t�(CF���8�}6���ǥlN����?����;�Y%\��������jYD:��h��/�̒�P�^2���z���L:!?�Z��)�I}D�|�,VG�F��S��C��LS�`�q��{:�˿"#�x�D˨�G�]}�m)��V���>C�5s�i2�ن��ōi}p�F�l�g��(���tJѮa�r9!$<st颐a�h>ƫp��eVqo��Cv��Wdm6�L������$�ޭ
���I�y��%�C�d��4B/s�k �<:��(���C/{Z��^f)x9����T��/z&2�q`�vMӄ����;g"����	s��������S.BC�� �ANa��\L��/U-�f�X���Wxχ'�v����Q�tGH�8����N�v���q�*b4�0�[j3�R��@���V����6�UI
��W����v�U8Ӂ@���~Jce��p�oI��\�K��S�k�M�)M~��C��Z3xB��,�A���XuI^+P��\*p�k�	>F
ޅ9V���d�S�>�.�33����m7�����ڡ�u�=v�f����8Y߆x��~�Y���bߟH#��'d���b�מ��sqf�eh,�B������Y�'����T�`:#1���JQ��+4\}��x���'��vU�������!�h�����Gdل����;��j-L��g?�����$�h�&8�����y��:ͪm��ܣ�y�R�:|���s�Ru<�x�sd��vi+����~�<�3K~܎F՛��\!�����ң�}�]��u�x�%� �������0߃v�N�%��E�M�6��Q�y>�	f�0ԏ��� s �(1�DFD�iÅ9�cL�`��A-N��;�z��h�	j-��bt�+,� ���A��:"���_ɼu=�>3�h�/Ք����&��+�Y!S\�T��YV��ߵ$���@1��Ã��@���{�|�p�t���L�ENRPu�R�s���sePVm��ܠ��$J���w�B����(�@�2����<
�ᬓ@"P��'�R��h�o�N7u/ufZ���N���m{�`�)a�N���lB�-����iӅ`�|��ɗ9��He����t�:M��L�LpT�uW������? �5���BٖvA�� ��� ��;s�n�R-��r/�U�pZ��4� 'ê�����T�I4/�	���J�!	Xɍ((�bO&[k�Z���,nB�~��oz����������ɑ��ٔ�?�k�����M��tBH�@�l��%i�.���k�Zd��T��4ɺ~�i�<
�$wNP�!P�6�_�>e��I�l�EKZ�
�׫�����<�ݒ�T٤��C������~��d�8C�����w�#�n�,3_�w^]�M�Ι;Z�����m��;v���(/�w�` ��a��ְ�(�?/�h��-��l� ݤ���^�'���#�&w�s��_Ւ0�`b�?ZQ��TNOkg=�O[�0t�/�����\��i"�f��;���[����zQ��(V|z1�E�-�"�d6����q��rػt�3.�i��XuZ��!
�E�k{�,{M�p��j�A�"إ	��X�0�C�5rGb����B���@_���2�ExG�ѡ�fY�,��R]�(�g
�A�l��_~.�@p_�,���Bu�?=[�ձ.o�L��c�K�N��\�z�g��O	��=FÖ�W�F�!Z>��'O�r"��.l�	��!��K#����ur��O\U��}m���v�jx�k��r\�H���d�=V�P �i|{�wZ)����
���W������<�!$�� ��H�4&�і�XhYM|���'�p�M����+�C�p{U�Ҭ�إ}�(mJ�|"�����\�qXj��ty��;F@$��3��p��?���/�0�O�6~9�czp/�����\�CLG��ڏtUR�(D���)Xt:�);�f��p�f_�8S@|�Ӏ�j�Gw�g�v�-<~�)��^�p���T��dĢ^�_�8�6n��ˁ��AE ���v�	A�(�µ�y�4�`K9��Ft���@����.���^��?�ē8���~̰��L
�7t, �ub?����Q��鳑�� 1��TM�xf�F����F�L4#�;�K
�8�]턢}JN8͵R�`vB�,�*��˖6���5�&*�Y�-�U\<Bk�X5w2R�G�8�"C�Cg�N㝺qY�x�;�\H�Vp�(�� � ]3�.G�sf-fS�.o��_Iߜπ/�|ۋ�-�qh�C�P�8�ԩ��x<"/��`A~������nߘ��Ǯ�����.�3��v�=%9��I�B�8/�Xx�zʛaHN�#��å	z]��� &Z�k�<O)ԟQ,>��u��ǳ��n�Z�w�w���t�g>��IQ�廔�Emff����Nez��+*��v&v:�iY0�n9�/t�Xf�o��7�J�l�����\-�>���uv<	�e�{�� *��.m�6slnr�K��'�c�����8�9aІFV�0n��^���qY��=�|k��$8�nd#s$�Ӡ-踿 ,��<��Kl�� a��%&Y&��� V��N=�7����c��ht^٘�p�:�p����Ą�˘f����R=���3�,�%��DZz��+8Hn"#�g_��#�PY�	�F���jB����j���-�#D������/��0\��"��Z���I����mܫ�6�o���|�/O���8󍽼��?�|9͆XkH��aK���Η�x2E����b��y�|��;��j>iW��\�Gw����dC0<Ɠh��~�~]C�rl*"4��{�e��|�ڢ�~�?@��ݫ�����ŲV�Q�m�N�wD5F�+h߽��*4��Z�s�w?�pk�'�w�<�i��3�Zsfvͬ�VY�c�lk�����,�LP�6��RJJE�dT���w�A������?���VKv�m̔�9�
������^�7�����4lR�6�����_�>�H��&���s����A�+����{�
f��V��L�e;̢�1�~2�U�(��켃�p��R��qu�"H{B�z��k�Y��->�&
耡�PDq'��4Tr� f��g״��>Go�+���w����x��.�΋Mm�`�5��RZM���r�sL�Dt���+��3�ݹ��׌��6yf�S�&��T+��W�b&�����T�#ta^_��b������ʮf��M6%�%�6`���ŭ{,}`<c�#	��N�_��������Y-����?c>o�>�7�Onn
x�zx�Gr%�W%�le�yM����L��� CKާ)��R�ߣqy���������s���g{�U��d$�u����jR�yȮ(G ���Ę����Z{gԻA��?tG����eUV�@���
�p���p�7�@�A���+�a��%����� �nT=Up�h��~�K��9���3�S6������>���ZJ���Q�!�┴.�w��,<[In�R��T8���qu}�T�m�R�˸�,����"�p��L�nbb�`eX��>��s����[am���fMז�m:��o�h-H��5^�?�������5���4a�zRn����'8��ر#f:T���;��IHeQym+}��	��n?��,xGg��.f���Q��In�Y�f�	)3�`1��;Xh����IT;q���Gvy/�΋�q���c�����p��v}c�P,�6����v!Z1O��!
�L<`)�Ͱv�(E>j.�8Ճ#�jv$ ���5^S��y+#Ch��:G�70�K�E�C��D��M��t�K�Bi##X�aa����BF16�=�����p�'���x�b]�\5s�7]v�ٓ�.�K&�=��Z&\�j[���tT};E����]��A��hB&�L�6���?��񘹄�8)N�����v�r�XTLg"�	��12�ѣ��,s�W鱕ʋ���n	�/�fb'@]�72zI<GS�p�&]�B:A�@���pZ^600�#g[SD�ַ��A$s���L����C)������@4��{7��n)��a�]��u�=N�T���%������ �L[v�hٖ�i��J-	-�4�A|��Z�{^E<�-rOy�:Ƞ�}��eb���#���W�`d��~@�� V>Dq�Ե���������Yd��51��wEz�:X0��0!�R��Y!��qI�����ܱs���X�<���������9fZ��W��������P��Gd���a�)�\�xR"��l� ��=d(��m��Lm`r�8�e��d!W!&Uy�q��%C!�t�M�-��ӹ�(�@�r�u�Ӑ��8̆OB�Mi<�zx��).%��EAc9�%�k�,i9�Wˮ�Z��$���.������l���	\�6A퐹�Պza
�k*F>�ohw5=��1���L�&V_P:(}#o����NT'E� ���$�a��b��Z���ќ���S���]����a�-<VE�=��B,bG�Y6ө���+����ngwa�Ҭ�ܶ��zktldވ�h⽒=�^r53�hC�ȵ�A@%B�L\�f�X��Yr��ز|���y�BA��<���ȝ���E���E�%���~+1�V�����
������,�SS������7}4���������Y*�Y�nX�@F���?BB��U�j� 8��ʋa)5�w��|If�.|3��x~��aP�H��,\��8(�{PJK]5:=�3dL0�Pd�_�I��?ɛ S隭_��S�2D�#R�$��WT�B�̪�<��=�C��-�Qnv��f�@�q����@���u�=Y*p�nUܸ<�+�a�/D��������+���.�b\�����K���5H�Z-a-J{��>0�P�Qܩ!}_<o�Ϣ�*��y��y����Lw�Ц�ӄx���v���K"7hZ5���Tx�=�s�>����
����	Iq$��>���O �L������,R�>�Z�aI:�5��F��I	�^zM�Do����lo��Q͑q�f�`��G:�G��2�q���8�e����h:�o&�C�ظ���C�������&��1b)�S�-�P�s  V�e����		 ����@����mR'��s�X�7��L�N;�������0w%φ�F�[�����AGJ�*����*
�+z�b����[��,�`G��IM�1�Q5�a�w�eQ]D2`>�OW<��ɓ���XR�=�P^<��٢q�S�/$�.na����D��t�85|C�9���}-�1?ߢ{���m�|��\����?���^�z��)_ɫ'��)ԃ;$�r��0�#se�����|nO�(��Gf7g=��&v�K"����=�75�	n�!/.ƀO�*��=jq:��m�`�8��l�t��!%y׌�苂�%���z]X��/2�����]Zc����kD08�-'U۲q���Qԧd�r}T'8�v����ܹ�:�D@��)Ե��S��t�;����zzq��І�>;!����(�M��%*����9��M���4(Z}�P�.ú>t�x�R�ɸx<.�R�㽉g�W�������87.6{P��6�<8ь��(e)�H���x�ޞ���*Q�,��L�i >yjgl�Rx{�T���q�Z?Dw|Nw��	:r���O� �>��K��Ug�ÃXh�]����O���&Ԗ�������-	��,렘�!��k�-34/�
:�0%��4�������[������g9��C�z�2�s�0OV밆e�6�E�)E���*>�K�G���(I���';�]��#�o�9 '��ˁO�OJ{x�t]n�T��QE�M@����3��XT�����^S�%}P�� %��]��A�0_�|��'�=g����kR���Rښ�D>6Q��V�bD���3�����g{{H�̑o7�,��&Y�o"�z�)i�*�ؾ�CX�5>c��o1 �l��5��`�b�#�p;�R%�@��=7��4Ǎ�2\���JP�u�A�Oߡ�]���p4F@vc �ɘ�2�<`ҏ��v�>���Q"���|B"��H�P�0`�:~BK�^G`�i]qT�h�p�RC��AV����#I�ltP���8Ѥu��b[�!S�@�V0U=�e����̙��1�L�Z0�+��^b�D�-��=v�Τ�V��\�3?�P�'�?�B��mg�A�9�Uש���O���;j
�;��a(���Wt~*�Z��<ۄ��%��B���-��x�vƎ7W���'���J�Q������3���l��_^XN��`(��>�z(��i^�z���'_��]�`��d���l'�z���D�/���m���S�ŷ�Ȑ4�W���3�{�膱�
�K0^̺�\\N��On��jLk��g��t�q[��pBL�i�f���`��?��vm�ѢT@A�)i����L�r����U�MPȾ�%��mL;�!�Bc�y�!�R���=����z�'g��%�dݲm�j
�WA��^�j�Q�qz���Q�b! ���A���bV���������[bl��� �H���l;z��m"�g	
ř͟|���'���������b� p�@�) ͎�j����M��L�>D�uP��=X �:���e`+/T�ɺ�;F��z�9/%�(��S]P`K�GG�d͖@D���=�*g?rj��7�5^��A���õ���"/2��љ��>8�"�F`9�X=?���jN�@P��'��E[I�ju�c&^=��Qٟ��c�J`�zn8�Η:�����e*'�H��y���ϹF�-�ʂo�/����a�ުn��*�`d�� �m��H��j�Aܽ���t��&iv褧z�#����v��@��~TM�2Z�	�o�詒D뼟vXAAy`�Z#V��P�]��v'!���l&���;��>Gi�G��h	��B��0.�m�5��yJ�"&[�\[u�Y�tɾp�c�R�zK�39�_��p�NW<�߮��R�n�[�(�]m����_˃!MOU� *�!+�}��4�q�Qck���d��A���HN%���m�iޱY���^�]�|%ဴ�%;�ۗ��>؂��!����.��<D� �����g�DF��u���h�n�,	�����je�,_�b|�=�tC�	̛�ܞD}��i������ǑM�;�lB�X@_�z]����j�Z7�Ǯ���)�խ��Q���Ƴ+��}JI>u�,�bJ�<�%i1k���R�� ����V��=S�8�^��i?��	L���Β��6���f[�tu8΍�zhp,��}/ѝ���֠sɌ����5�>���sT�/|P���2������e-v�2/��-D�爂��ʲ0�(Qb>�:�����V�ᥕ���9�M,�w��u�������κ�H{y9G�\�+T+S����E�����1��c5Z1�"��䫶�N�鋚�d��0�k�C	s^-�d�J8T�Y�@��C�f��j�* 2?�d���0^MO�t��[}d�c�����$iDU�E�ܒF44!c����+�9�����ړV��-��6�V� R�^�gz�>>Āj�A��	�R���<K��������LlI�>EcM#��||��4tGjH����od��TV�|��#+�%Vx8z��~j��ZՓ+�*�ِ`0��	�<��%�{�� �_���W��`�!?��n2��}����$1�|E�ì'Ȑ��=8����`�i�8>hsi� rÜ0�0�z>�J<i��)_(x\|!�6��N1�7��qLn��	C�n5�����K��t��n�˥���׬ju��m���"�V�A���0ut�K����c�BȖ�a$#N�$��-�)���E�1����9��q����M�G$��a� �M���g[��%#2���f¡>1�|�;E����r���[�\̓�5̍Gq�`��b��5���1&`�z�eȢ�~�������J��~=�w��J����a�w��N�N���rg���2ى������4�`ie���.�T%i�2?ހ�%��Ĩx���" �hߜ��R!���W��$�e&Ɣ�{�K4%�A��9��X�����ڊ��^�h�o�����ٵ�o�H����F�xb |_>M�Rn��ͤ�,��7�9�?НD�ed����I��F�w��wA�vzj�S�n!׎�Vr����\\ل�EP;�&�xh������w�]:ão��U�$vV���
lMޖ�]���7�3C�&������"�y�@��>:��x�G'7R{ɊH8��=Z� ��遨!S_�&yW=c�J�e�E��.�����֩7)��?)(������C/(��,	J�(������$\T����Af[�2W1����aA$��������X������P�q1#�GJ3nI�z3!_
��:�hZ�����{p�1��ψ�c�f�r:�g�������4�+#! @!Y�c=�j���ޑ3����7��h����%��q�߱r�Pf��/鄞6�q2�<�9+�+�i�R�V��I��~9�f*}�*�lsE��������VQ���#J�!7�VG�j���MG�ʀo�նߣ�A�s����+��ȿ��E=�0�>d��f˞�Β��ҭ�q����ݢ>�Jt��q����H�T��'0����[��i:������4�f�F�e��[{'n��Ќ�}�cC���}g �W�#>�G��3Fi?�D�$}U!��ab?ը��d߽�.���ƻ6�*;9q��8���k���V��u6��у	�o��4�S�-�#WGǿ���6jW*�Y�)0����
���Х� e���×���N!Nޝ2�;��ɻ~����.p�Q���R�;-�Va��f�4��U�|H=�?�LI]X����&Fi��H��`�;�1�������t��A�6�u�>\���=��O�^!s_�wH�۪�d����ٞ�>�Ě5���;��Wj��4*�>���;�Dx�T}�;OW�$b��G��{����<�K]�㍿�oܳ㘝�ζ����:�����.�P^,�g�;�^tg�tf����������%*��ᖑ~(uy��t��\��}��?I����mJd�z�W��GJ��`J'W�M%������k��g����jD>��3N}pF? ���ſ0��Yv-�D+�+o�*	x���u"���x�{�'C3���/��S��0��ۆ;��s��w�>��A�Zw�<����]�4�%T�*6NE����P���t3su�S'*��"�מ M]%��l���
��n�4|?sOb�����U����5��\��1�A��!�E��Sr�w��=�����gHw>�rx#�"�;e�(L��|�!�5޸I��*f�J�A��E��P�T��S�ɺ���0��Pq��84�w{bh�F)���4�`f��W�Z-�2��۔���["���<	��y���l��0m��Ƅ���bW�!E�6���~��BY������ ��x�-R��_��cy	�t��H���^�c��}�Ⱥ�%��t� �l�K���/�_y�;�������b�jMQ>�B�=��\����7x�	�#y0ՃX&���0p��ݩ���]g�@vh��i+�$�Y# ��#T�D0�{a]���ClG��S���(���a�34�I��u6i/����4��ע����[W"�i9�sd����ᴞ����O��v1��8|C���C�{�)lF)I�:���. *�x���X?�(Ш��Ds�@ vISȥy�$�
g����󁱸�Y����\���d~����Ü���C.O3&��n�s>�9�p><^��.+	K9�铒+�$rO��Q��/\���>F~�~
a����&e�P���3z�AT^�G��:��q���Y�H\;���ڿVC�ohW����8c�'a�J��R�,��7�ΈÌԾ��;�'}�^�f��S,������;y��0��2Ue�V���w���?=���W�d�	d֗���q��bPh����[7 /wBȌ���H�5���p5�^澲0��#��`��B#o6
mq��k�!�/�dj�UAA��5�ـQﰽ�$/ON��,����)$��~_�H�_��lPwE'����~���$^�z9eRC�hʤ0(6D����8�I�py�@ �h!zk��ڲ1�`��(�|��w]C���ř�J/�"��+�/�ͤ^�*f� d�p$�� |]�a�me���8��Rig�-xO}"���+������S�f����]�E��6�P��Ca��lu�,3�v�#c��n�i�)�������IOX��<}心|>:z�"��@�4�PDJ	⏧6��>�SU�1�������Me[H��fv3R�~2�v�p3[L��p�!��Q�K��#��r���2Y썑=��j��}�[=)�e@�['���г*#%�����=:�^K<�U6n|kl�՝��'ý�9U/�l�nE��ϖ���[�;WQ�	�.�[ϯ���T��� H�ۘKE���;
����L�/�\U�wx��Y;t"
�a���ڶEF�a|i�B�l}�W�Bm)�;���;°x�������L�����]n?���H���'��ڝ��b�����ߏ���W+;�a�2(�X�^�b�$.e�����g��9�T���<����`�r�w�Ģ��x�t��)�ol���(8�_1�hp���tA�r��ҽR��H�^{������ X��3-�1�%��K�'���A����8{�
#�=:�V1�Q2u�UȻ���
O����M�sҽF�雫��پ9�ϵ�]�=g�������9SL�6 ܦ]-l����Y��,�4�; ��^��%�]�і ����&YJ�3�j���	[���X/��azӆb�a��{j�%ԇޑ��:$6`b��B��b�Gk
Օ��=ME��؀\���,��u1������L�ܟbCx����J�]�@��%�V�O\I��1L� %X�U=��0�ڨ*7�#u�/�uub��\�9����!*�?���|O�J=
f1����2m" |H��\QG��tYI�����2Ŷ�l(�����z�����ܞIo�� ����h;\}��p1@��S���Ѝ�m~*���|Y_��Hkoe�"��Vs��������fq��
�s$K3��S�Z���IPt�����J������&Z�	���sts>;���LF�?��k%yӴ�$0���궺
���|DCG������bz�=��I&Mh�V3�������`P�«���R�e�;��M3T���^�ʋs}#c:[�#�����5h4�l��Y(��h�=c���r��N�P�,�0���:��E�=IA΋98���a��lQ�5/��(���b ���tؾ<��`�D�O�DO�-u�=�,F�� dsX��9s�k��f�*����rC����1�G$l]n|���]�dE����k��<�&W�0Jq)N3�*b����zᙍ����D��=��\��`��}bzm�Q�MsGa?,L�o�E����<t*���#'��Ǘ��@�῏ْ�y/��G&��8HQ��d����x�>��,��}(�S�h/)��=w����ӧ�?��E,w��1�N���H�@3/��ɮ&I��c ����֣{U�w�>TS(�F2Ŧ���Y2d}��[��>S^�L>�Ji_U6fj�V������N�GM��[�w,���fo۰�����k,#�Y$�e�oq��= ����n�)k.1tŻ�4ᘳ�τ9�󝂠ӥ}�C�M� .��t���-�(��X���\�QN/������X��)���:^�q��"$���xJ��J�l�Do�������v����=#�:�
K����W9l	=�2��Gf$g�i��K�X>�i�'9GKZ����M�WR ���Y�u p^휂q5<+Cr�Q�D$������U&-\{�3Q���b6f� �����Z��gz�1�H7�p?5�W77�}��#���U�Şyi���}1J�M����B��`��A� ��>�yp���n�5�E�?p��S��:��y��A��Q$����l�L�Kv�U>y-���/e����4Ra���7�;�-��;��
g6Ѡ�F�6w�~_k�J�'������e��N
�(ɟ���6[�"���vv��m�%+������L�~��Y�ad}vQ����\����
1\�U��`�g���_�f�j]��b�
�wE㏻L~�g����E�15�Y�Ї�m31�����=T��{��U�SP��# ����m��TY��T�h�r��!E���e��z�5�-���*��g��f�Zm��Y�����̬�Y��m��R
���,$��y�������\�Y�W�;��%�S�@^��R��2�U6�����F���4&ʋk:L#��ˊ)��©;y:x,"RU8Q�Sq���M���)�����F6�k�NY�T��᪹�&鷄8���F�]\�y�~�k>�>Z�* �2ݛ���;]C��fw�q���3|����Ɇn���2�g-���Έ~c?^.���J�㝚:C�K�O�)Rf12���KL[!`B�%��Fh?��r��M�e��{����lUOS	���0pk�2��\�K8p���8:JL����r�2��&˾q���(�&F}i�W Ϧ��T��'_@�"�=�u���9~#����f!�:?|#�����W\l��.hP�
�����/�p�qQ3�	��u��;dٛZ:��};�Ȅ�D��q��8�2
����w�"���q8���p��I�,�46�������Զ���
�;s���Wq�g��4e�K��M��+_+��>�N���E/h�T�f~F�V��cl5���ח`,������k3���2���t�^�,H���&��������J�Z�w�7���j�¬ʕ�����e	`���gyOɤ�P�d-2o���E&LF�j��+6ߡ���4L�;�J/�9	d�9x	>W����j#�s�˫�u/�F&O��Ӝ��%�ה�+�O%NݐlC
������\��%�F�u�5 &Xl�|�&� n!��ի�,ϔ�:l�ʾ��'Y��C<���*4/M!B__[�eb��(6�.ځ�e֔����lnփ>��3sp�nsBT8�Зi�Y�����v�K'5�����f���  ��5
yM4:}�L�,=�T���Y����^��3w�2�������&=��~�����*}��%���n��l��H��������82~Ε�7'w��)[zj7��+B�S�=�0� �1��v�s��R����8����O���2��P��e��8l�*i���%���ku�)�W5▝}��1����8�X�Yd�����|<�C��;���l���!��T\Q9mm��đ7�Rxj�F��$��7$���$u�/��kyp?�4e����
�ړ�"��fΓg᢭cC�FZ�	<�<�ի?"n@G��{v�ɗ j%{X3�7q3z��*.����x��#��v��cm3���~ J\$=��og{��pHV=Ԩ0~�D��|��4V�	-Q(�,�<�_S�s�,��(xO7����I\"!U3��v�y`�Ѻ�o��@S�!TQ��'�� @���sdr��3=V���?4�`P�`|<�d�o��LC�Oz�N�ܧ����怱���<����'�B�Y5����vYw/�}�5Ԩ�L��&+���V0A���b���np� ������1�͵���q��+uD?d )�3!���k>D�)f}��?��V��ś#,E��Ӥ��9I%�9��l�jWEHL*mt��lo��j6]���N���o�ߛ岠�1G1������*��� }�8̒n�� ����!7E-�{1�%��c��=L4'v�������r]c�D���A\_7��;�Z��>�!+�5�{��9���t�u�CՑ==ߝ&�JYoO��[��[�v���GO��va�)u�-��9J^M�ZIs��Gn$�Vנ}-b�%��*q
�G�eR4�%><��i�x�'e����->�^˂�,F�BM�Q��U�Z�`�"gWSK[h���.��Xn���T� 6�٢�EF,9�<}�c���<Eq���T�D�x2�������	0�!�W(H���{�Gq��rq�(/K�澍�3nUu֔	#SQn����!�FxY�J� ���*�j�>g!ըҢ����/����C���ǽ��sZj�
鐼4��R���A��ͷ&w4_����_޾Ed�Y��v�k���X�7L4M5���9W��I/�A���Ƚ�/�]��C��D�b%�Z���l�uʲ$'7F�[YI���v�~�=]���z-�9���b2wL�(� 8^l]d'����a'!o�w�[�h��j�Ψ��ۂ�U�U�;y�|��$ a�'�M����$��E8���%�!�nXؚ�y< JK�k�r
���T�����,�hu�l�����0����$��;Υg��d%??�^���p:�=�7 
3�q��԰\jX�*s�L���QwDt�*K2%~s+�p��mj��nB�69o�e
�yJ�m=6B��ɏW��b�����Ɛ��w�2^����<�|D�&��x0�ǃ��}ct�����n�<�+�������C^����H�����TFG�)Ǟ$�o�f!#9�RX��H�]�3�nG��bڹ�@Ac!t�.������Ec_�b�O�.Q~�W�;��8%z��	r�TUop�Ew���V�c��@��Q���c$H�a�)�
}2������9���xҷܤ�m�<i�
�&ᅵO]w$��.
�m�Bb�̴ٔr�G�.����We�,��y����S�~W����SWx4g_	F�BX6Gs3|�`h���d�~�Wݥ�a�H�@]���!��P��j+,ꅇE1i!�B�oݡ�!S���3�;�f�:t{E�(�8j�c�2o��H��a��]~Z.���I�P?Q�/�)�'�`R�M� [;��G⦛����?��˚�x�bFA�$7U�7�9��r�>E�9jq���NĿ����A�f�M+K���"�Y��&9rg�&|����;�S��E9�VV���������'s)�d
�>fY����?=7
V+|��j�P�Z�J����q�m^r��_k�0�
��ٍI�B~s��b��iT���WG��еĝ_�Ѡ�٢�'Y�Rpy�
8�:K�R	����I���؏a`�+KY���.*ڍ�~ U6���d����>g���ܟ��L�����[��g��O"�[lط�9���:~E���S�N�9��gٕS:x�~�p�a��%[��e�Uɞz������u!dn���m�ye  �C��=���nnƤn�o�vNgE�a�y\���2 Io�!��u(�+�f�?z��܂�6TY��i�j��	�/��bq��4Y��u/��<X4��	�T�=5�u�4�b��Q�әE�;"L#��� ��v�Jf*�D��qT���{�Hvu��~���Յx��"g�J�Ho@o�5]��E^��.Gz��նXo���;&�Ef�C��V�m���V��LTO&i>é����|�E����;���(�R�ؓ�e�b1�{nU��H�ۦN	l33q�/�ޅ'���MS��t��_�!1]�z�{)�c�J!�dU��)mu�·�s.&��d<���%�/��vm3�H��	o�Y���PC�&����(��}K�Z���zwcs�J	_JЋ�;0��s=�NW	� ْ'��Dkx5^Ts�Wk�9P��0�{ry�����h�蛜�Q�W
��n�]��7��c�� (#��C1B\��X���@�J�ϭ�;��-���� �G_�<�h�I�G�M��k��(Z���7K�E�L4�|wa��9.����- �w[5��
���(��r?��ɜ���ؼ��F�S�%8p����W`py�n�Y�W���A�om9���]ydj�c ^��Ӗ���cj�K��y�NS�&���<"��0+=�.���E�;J�٠�o1�m����؏H���x�B"�1��� @����۟�Ba���hr���������b��
6rY�Xj�]�/Oy��0ց�k��?�z�N)�QD�w˩?���;�[��m<v�fԗ���lιW�%��}��g��*c4|Q��G_登%'ډȋC/���t|u�J8 h�:`f�Wp�9��pvK˪�7�+㘇L�+�<G�J������*#�:��H�P
V�a�u��[�7\0M-J���Q�;��KN�mQ�!��Fv�%{Lr}N sp������5��]��#��	���<��Vw&&/Ӱ�>��P9�Ր}c�d(xyQ�f1�@���eǔP�jG�*��v�+#��޺)Ѱ�
+���24_�[��M���%������mv�J��(7'���������U/%a�	y��a�(W/�|'�"�@��S{4ѻ�K��!�Ģ����Z|���w��g+��ۉ.�'����JN4��	�i�i��a�2z�+D�*δ����'m�sߧ�]?UA< �����k}���W��M�@��--\�,(��T3e ��L	4VuP��,�e��(uD�N�a�I���o����\�|��U4�|rq��1���.J����e���NA:>�>��v�me�Km7��x{�[ƾ׋VE�IqO�u��Qat`���ؠA?k��摉�Z��h��������D.�$��������3K'����p��X?�ΙE�v���S<�}L�E̗�b"��x��y���gU�ci�Ə�� ��:ߢ��j���UvI�T�%���r�q���Q�%-�����Tr�e��D��O$`E�(b���CU�ٍ�8�+;GH��j�:���f���+r�S/�5Jڪnu��ԃ!�<��p%�|.7��:a'�F��t�^�O�Um_u̞Dp@}�,�.��+�!�uu��=s����l�b����U���&������6��A�8�+��A�y3ٶp<�)��d�͌4<
��9i����J��P�X:�oNhWz�k��f��~hĻ�?�¿q#q	E�|�w#qq�3���9����vU���ŝ�<��Z��?���'P\U'1H��02����Żb��i���M��Jl@���p��q�w{��pJi�_m��/���m�s�5H���_���]�u��9�~�p�ju0㰾�!H
Ӥ��<ƅqM��xa@p(]i��طX�qN	%�4���&��0-u8����`�C��Q�ﵸ�G*ǐMI���\Q�)S�c�
�6��+�0��B��=��y��(J�a�N�䅙�EE�)*^Ǌ�.9�1�=SkW��&�Ҙ"Cu6����v�ؽ���SK��~L�����B�_e���6̔�]0<lUY���Ӈ�e��/�*%����|�����Ii���o�2I[����8�=��]�.n]MH��X��d�0��65k	)�֑S��ĸɝ/Gu\�f-�`�R�����so�C�Q�����K�[�:�	I˽������+���PW]�,֪QrJd�6˕��y��#��֚@�A��*u�Voj�2Z��#�IL���S#Eܚ�թ��"�\�F���x�t4��UU�bY%�<@q&���ǭ<�)�6�7����Ѯ����$�p�E1|!IU����ް���Jt4�^jq\�ɲ����{W�R���+��KC.^���AڐR����I0�|����2\TM��M�m�� ������oN|Yv�/����/Oy�1�@��p#���H�YP*
���q����#ng�k�L�θ�*���O��ýM��t��殺6]l�1�0�?���9dmt����3߉$��.��or9��>��{D^I�lWc�6��,�4�Gv;S��4���wK�U�Y>����!Gu���q|��W���u�ﱅ髀i��E�$n�����7`W{vV~\p��&=�U1=��=H[5X3�iu��̐ٹ'�֯=�g�`K	�����Dtk�5���ljM�4�����k�|��E��M+£"j�%2>�IëA�e���!߃�A���%^��h��mo���v[R|���:P��$oY��ʥ̎���@<kѽBE��)�@/�?���� ��g���i�A�KX�Hz�&�w_��C|/��.a�ЕCf��y%�EU��*�ջ�])S
\X�9:�C �B=zVO'>`В��eZ'1�@#j������wZ&�p��(B�I���be,&��c���?x1��������[ׇͣ�Q�K<G���Q]<J��v��\�[L��,I�"� ͩ{��	����}�_��K�6�؊�07�==u9�����o�_�������1��V��cVcN����T�m9�J��6�u ����i|yx�@�#QĴʏ5�}Hu��
���_��~�`a��>�d/ γv%�a�|��O9�ŋ(x�)%[��:�G�i&�8ܜ�r�I]l����w2���y��C�~$�Hq�X�qc���B�M�%J��r���X�a(�2�W��f�
���1�y��<{��+=�$�Y<�]��A�"��J/ü.j�� k�-1�u� څՑb����W"�p$c~1� �_8�*e���U<���6*{���K�WB��lƏ-aA��R��;t�6�D���#4�4��#�7d][6�g�]%�~69�e���CA��"�F�c�N�8�aޖ�[�(K3���Ñ�Cs�TDEL3��?�"���F���_����quq��*�r89��g<��%�?:�
���lm#^K��Ie@cR�Z��r`��霞��K�d��8�8k9& O�*ceP�w
���׎]�c��0�9���A�2X,��jX8 %3��-�\a��42�`�1O��e�]Q-mr<���-@O�A����i��'.������G�4̧ �*x�V�e}෪EؑNO4���#@��k��==��j�	�s����4��a����B�oa�N̘�WR��h��P?Jvo���%>�.���
�H�)��4d���qf�C�ES��	`z�Ж�B7�y}��H�5[f�?E�e+��D���=��3�o��k��� �`�4�����Xf#�9��]�Ib�1x{��ԕtN�
$����{ֱ�Y�B���X*�78���IP�c� ��m��w }9Fyu7�qJ�yw�=2;Gjꯙܺ��h�qD���g��z�Bl$�P�����s���C$^�s�)��#�P��@�j�ܶ'@d��'L�ȯi�r#.v)B��itK�n�w�g����޷���M�����  �C"ڿv��{�	��r��2����`�r�ubU���~C�����Ẕ;m���c^�V"��9bd[�k4o 2������=g���]6�q�w�L�.�h'��1�+G|�_�b�1�"�1�P�#�'-g���+p[����e��Z��*�f��]����8�_iT%0+���Z��K5�C� ��������i����rY�����k� ��
@1+���/�F�t�$��v�h�&*˻{�l��$�%B�)�+JH��>�� ��­����"�p
6Gef;��b�4���Ng��=m���o*-'�W� � 0�wG�@��7���Fj��&<Z�J��G���ޟ q��U^HDAH������h�D>�t�i�bg���K��k�N�������� V����*�9H1>G�l^W��@��&�V&ۚ���po�i�D�ӫ�ۚ.U��g�z]�h��}[$Ÿ���Yep�d�5��к�T4����õ��<P�JE�pM����k��[�6�,��.��btjcV��������epOM������5FUی�x������kG-?*��)� �#�r�j�Dzl`b sJ�^�������aO3?Ë��W-�Q�R�Ŏ�-�67+�]�2�� �MR�35��Ͼs����n�_"�TM%p�p�2cN8�L!����U��C�A�|��s�/��ݚ�b�J�� ZXEGC�ĉ�E決�aL� 
��\ٻ�� J��;k�E�!�[�ML_��R]������<c��	�Ce�Rv�p��%�Êc�Z��-~]���#Z�eTlv��֐�t�G��8��{�/Y�����^Q��G���/)I���ˤ[E�LX@�$�X�S����T��t���:�߬��y��o��y��IaR��/~xvW��d(���+��eY.�4fp�y���."s����O AG8Xj���bn�FL1S2,����X�և�#�!-ikG���>�?X:v�r`���V �Ihg�M�Ѭ嵾�R�2�B����b���L)�=��!�\\i�;���o�a����cj��1'��bd *.~� {����w�lo�n�[1�.�X~�{@�<DGɼa�H�c&�?�S
0�w�����V��o���$3&���H��.�O�����/OV��-A�@��8���������X�q>����QaWJ*w:���1eږ~�Ef��=�~]�b,�u\k�6̔ȽO�
���Y�L���Ds�*O8�`�&h� O�cvL���.�����SLl0��5���<�e�/�(���_��$B����s�,�,i��n��7��3Y��(��I�y�o͸gbݸ�*��r� "��#�����lDNC�-%P7�BG���U�� }�-x�ˑ�V�Z�I"�{��\ 4���3�a�.V��]�-4q��5��:0�����F�zdu*Z����Ĩ�L=҈R��:�PY�^L"ZZ��Ugҍ�Uɢ��[���hoG�Q�S�% �?L�����r�5��Б�@�����8�n?6ֹ�?"k8�Մqhqʐ/sBobǎ�E������s��A[\K�!D�Eu[�E����s����� c�"��@Nь��3Fi���f��@Sl~.���ģ�KlH��:5��	_0}�S�>�����Eoo�����Ť�Zp
��TM至������@����e�/6��/�Tc��b�hY��b�p#w�8'��͔&�����9N�QN+�K<$�zQ�t�9M:)�]%�<Т���P2~ج�N.���8ux4���$^��0~M�V ����.��L��h8>9�Dr��/~k�|��5 �V�Fy������Ta;�ܣ��P�����U'm�|���-pX�؍����?
G�9#u؄
���l<��{'�7��p��d�3�x��0�X�O~~O�-#�{7࣯�NȐ�w�H�٩P�@�*���kL�ץ�/�٧��丹��ɪ(Ji�h^#,�[�@Z/��8����)���*�Ee3a��_���֤r�z�$Q��a8O��֘Aʷ�D��L*=%YLK��q<z�Pl��A_���p�jM3��A�@�cj$���#e�_17����`��+@W.��`����^�B�7�Q�mj���<Xe�JR����F�s���6��7s�p�W@���y�C������y�`D+�0?b�Ta5:s�ӊ�fqh���!g����|Fu���_5��e�0��a�$|��G�+hxV"����JP�M!��m�P~^D$��_B/�q��6W�b��(4M���ʡw�S�[�P
������^F��K�u����<�����䅛򂖓P�;���[)�7Ĩ���-�M�/�h}5=���^�?��`Ƣ��ɱ����׷�4*M��z0.�Il��?9_�mv� Iw>RDvyg�`��j݆0q�Krt��^�ʓ
�xf�#؃u-���6���`�Ջ�����1����@�;����FcZ�5��CW��B����N�v$�V� �Y&k[��l2�s�1>?�W8�Ү����2���
�����S�8�<a��F�/�B�ԟ�k�ak��攤�K��CV�F=�_�ӗ+�H��e^T��5��0��W��|���V����=���"vW��.�i��a�������i�<����+�o�[G���?���zR��,���l�H#�]��5�p�E�U�k^�����Ȋ={3=��g�5�c%�o��Y=c���mg:yY������E�e���\#��R��C��w�x�a��3
�K1-ߩ��ZHH�c݇���x~_���*<�P3N�.1�^�i�1o»��]%����䬡T�{g,a��[፼Ҥ��O�xPj�tdqi������m�9� ��~��Х�}��0��'�`P$��I�q&ѡ�~���-�u��T����{�T@�g��z�� �ح�w�ܮ�o�r����V�Abk���=�5�M\S��'x�ų� _,�Gd��߷��TI��M�y~xS�(�ș56R1��u�`���oç�b�u��Q���.8��4K��0Mu�b~�(~�iK��*P�/�_��|�ѯa�S�F��<9�z�G�mC�F ���P���`8���J@ �� g!��f�s��В��3"�s�H²:�6dj5�Eّ�s��k�eq�X�6���DXu8�<�+�r����r�S4F?����ռ��}RwE5�����
����3�y0��$4���y�>N���U��� V,�\�!�pa�2:H��]��*��o�����<@��`�6b�6<�vO���Bq+��jÖ�
k(XX:	�l��M~Gp��i�l��큾���ߧ�@H
�1D��Z���9�{�˻��
�
��udF���S�����;�XW[y�$��Rά�V���䳫־"1�.x���93�T���*����� ��c�H�FV>[|D�D%{Н�rXl)8�WEQ5k~1/��&��!���@n�g�^������q�qԶxS�4�x��z����(i��K${h����%�"�[Ъ��tߩ	���}�����A�ܧ��3���1혏��٣kLҳP��®�@L��ԩ0ށ���tQ����<"�����(O�����d4A$Q���e|Ap�;�ԫ�(�ƨ�,	y�#�����x�b�@߭�qD�>�4�����4�/�H�A��lI4t�I�X�[Ƈ@m�;U�4���Ϣ��M������Y��<Ӛ�Qe����(���"$��5�E@=�"*��et�H����_��:�¡�Nt�icm��?���'i|��=������W1؛�t���}����0�b�R���
]�z�R��Ȁ�VVم��yr�gBV�\����	OS��m]�ES��C��t������	����K��M�ν���%q��0��:g�2���{U����m� �_N�Qm�����l�MD����R#��(��Ih�CP��%g)���l�$�)�P�NT6^'��%2E��F���[�����Xl���3��ZE*��d��cb��T���}s�n�Eؕ����q$r� ^bZ�9�2������6�y��ȇcc�vlfԟt�	�/%{)Q��wQ"�>�ӭ^J�}�����_�.�S^�a��&BR��p���cN�X{�A�˲t��M�ӈޡ��W��'��dD�0���k_ !����"������
�\��|�1g�R�舾�4�}[λ���7�lX���|9�E�Щ��/�Ϯ�m��'fp:�{>�3�M��z4B`�j�A� �5F]�=QD%罾O���#���1�/6��n���L���7���a��-�U�!j�=Ĕ7����u����R�g�S�ә�IA��ec�{h��F�MNpMCx�d&j�.�M�}9p9�X��(L��lS��ٻ>xa�=Pq`�kb��RrO�d�햍g ˽��/�B�R��_�JӰ3��Mx�. UI��'��K9��P>l$լ';$��ia���v���ciU�Ϙ!h��q���) �+֨�l%,w&��b��N1��T���E ��MD�0���'����
�'z��+�F/���ꍔO>����H�Fz2G�X{i7<��l��f����Kcp��
xH�_w�S�j���}��K7�ڸ%���"�Ŋ|ǹz-0�P�Ʊ�H�i7h�Ge��B�F��wm�M�����x��6݀�BtG��h��
xѢ��~�7���VlIdؿ��������~�խq�v+���5��]�������w�R�1��;g]�������CV��_Qn@�dMM��q	Wn>�n)#�}Wo���~3|���I�*�,��R�����?���zij+� Ha�Zg��T��:����vet�����
�Q��m�l��G�D��ؚb�o��O�%;�c`�1����ЙB��﷫)��<�k]����}w5
�̸��Jb�����q*��_�9�d�:�+���$��Q*����i�w�K��R{;{X0��;FR�M����C�zYB�L�7a"�g^v p��3���L���#-1�c��}d�������d�E�p�4�Ј�O�P��
��ʣ5_�_(�"���	�J�}��j���t-l�`:NR�mN�Ϡ`�h7�Jb�{.�������"�UJ{l�]GМ�n,g2/�-� b���c�t�0���0u�#]���8�=�HE�ƀ��D�C^�q��7sO�ʐ:RO�����Ⱥ�x7D�%!d@�`���M.SoJwU�~yD��"fT�"Z@i�����KZ�A�v�@�<�0��܉h2i�^��
�*Ef"�c�F��A���
~���2�th��@��\0����L�ϏS2���\�q��*��$�=(k4��U�.oP�IQGg�&����u�`����~�� _�8���#p�����h�Uc��5B�J\�E�0i��ţK�ZI�%���#�3�K�}?���g@#� �rC��Bvo��!��l�6܄Hu�c�d���dԾ�q���d#:A�%��x���+W𲎄C�!Lx��óm�D�F-=���Z�}Tϱ�,lW(���p�h�_<hz�mP�'��k�����d�F�V�[M	������)���e�� ����~ě/ ��er9�4/u'b���6���Y�".=IM���F��?�<�R�3&wv�ӥ=%Ϛ=�zY�Z7#ԍ`b���|D��q��Pe�X�Ա�؜y�d-�S���x�\�NL2����;I�8N+	
tuR��Bd4�)H��e����<bSCcG˼���6�\�n��d�s.Lz �A�G�Q�gFG>"���;[
���}�Qen��@�&�O�˾�g�+p�����ըՕy/�[��E1�>*���o���HR�
,�v7��ȋ��G�d���i��؉�G����^3�3'O(̔Ř>ji�T\紊-S`;j34��B��~�!ʩs�:��S�ԉ������Q/?�g�!�mӤ�	l�>�癭���blE؊�8g6QU���aҾ�F���������� v�P�k�jr�r[i����G�GJ�8bCh��5�]�AW}V�}I�ts�+��J�I�;��Tc�bI3�D�����B�֎Π����'0�s�&��#a�.Q���&*N�᧝Ek���ſv\����tNX�nB����jΞދ
�H\�"���(b�,�k�W6ct�]�æ�/&���BJy�'�(�����X�M9Ťj����ӭ#�s}_ej��޽1��yO9<s��]1�J�c]ʉ)Zi��$���b�PYA*����!��clBʘm�M����)�\���	fz�&�NO_�,O��ͯT&����r?���ŀ�����6�%��0���v?��:��VJ�󖺾� WY��	�BQ�5ðr���Hǈ9�u<��E���6P����m�!X'�#������!�hK57��m�'�������i,pw���k`�;�\�yc�3�r�jC(�W��.�W� J�hȸP%ơ8v��5zq�tmpi��ᡒٰ���iyݱ����R� �;�IIV^�_�����*K���i���h�/x��t�`�U��{�%���_��:�6	t�b���V��~�;!�����tVg8��3�L��%�e��B�؟�d����c�5�؛��
�i|â��s_`Ê	B�J���b$��o{q$x�u�γw�GAtY�c�~���^��w��G"R�2�_�A�Ԃ5j����=�n��Z6��YX�1i�C�5�)U'�Q ��Q�����v�Q���K�h���ҰY&��h�u���p��T?�m�r�/Ll�g��;���v	��>Ym�3\���54i!TC)�jS����?�G��`9Z��ꈦ/|؛�}2/�K�����J�EB�(�<�������Z]#E�A�*��q�p���O�b?�,=����MDf��g!E.�af~�����bUaP.����^2�Wh1�v�5�����nE�?��g"��W+�ͼ�Q���M>�8�`4��$#%�8	:�Zu'�C�~�L��G�P��	��"I	���Z+rn����VC!tj�Ғٵm[��塅+d(u%U�k�A>���%�A���eȭXlߩQ��S�`jܫw����8M	�SC���Ό�r��x u�'�.Q>�uX�d��0�-�	+ͨ���#`�~h���Q uIuR�����_�3��#4^��i�?d�X�\�	/��w�(��*f�}lBXmV2\��` S�w���	\6���RT|���Z�F%�׈�[�`R�(EkS�~F�B$/�E+�R��ać~֖�P��*I6�"��R]���{�/8��˸��'yJ[�Q�Q����*GͿ�!�`�>T�i�	�� ׅ%f�&
J�����A$Nh�Q�T�h;��0=�]�9��,�����<^�rw7K?�(o��%�}����T<o��*<�����tm#�k��*�h@��A3ѡe;
קt���;���n�J2��/:A����kɞ�P�@��4�DxN��!O_Y�p�e���f�֫���������.E�����9�p��Ø	��M0�`�2����RG�P�4P��O�E�Pv �9kD)Ek���	w����nd!���!�86�5M��]������OK�0��U�<�Rlu����Ud�����>3���O�\��*�Y-�Q���R��2}�����+��M�?��%��%�B�a*V	o�Sd� m�@xHd\�P��yBwk�o��u�3LdI.�
����$���(M��U=Fş�|d G�K��n%���M�Y�G(�Vi���� }=!C:R9!o[�%a�^[����"����&��a�g O��s%��/���&3� ����Ghc��\�ݩ�.{m����V/霘�ҩ3"�98���X�	m����:�[��̿�(�x�LN�J��)Ź9P}������c�eI���6ߎ�J��xB贆�}fis1E%��ZaZ����Σ�jr��2�ʕ{����N�VfR�p�ytR��y=��s-.��7c��K�$����t��%?(�*|�\��@K�`Jʸ2a@JS��&�*�C=͟C����ߘe5+8B��M�䒲�:� �A�.g���׉zV(�K酌SÖ+6ǭ]��}�:������i�P��B��ao�06���d�Z4���R��};l��:\
����{?���N!?fB	�l��n�C�4��5B!�.�,�mdQ֥��i{��˾Ia�<>ͣ������PC�F������:��_�-�v'�g��;k�s�hQ?��2��?��_|�Y� 3���q,/`g�Y�^F9�Iq_�+�ִ��� 
j�e=�ˀ�]@�Fl��l~-�b���4�N���o\�و���ܙ��͹t0��e�ҥx����^���j��q�fZ8�Ru\�w���{ �*I�]l�P�;wѰ�Ri��qI��F;��X����������p(��gF^r�!H^�a	���Ɉ�x�$��W�%���pM�U.�j1���5gTg�L��$
z��M]xV'��ݙ�,���������Ee<)��қݭ�{h4=1a�q����Z~a�u��r�;w����am;����Q!���z�A���D��?)��e6�����N��sWi^��l�z;�A+n�ٵ�u���˒��N)QΎ
S�~~�vnW���e��\X�l�l5��&�4��ʘk
�� �X�n�̕Ce��e,n�ztK����Ո#�k�pnq"[ufC��J�=���jj<t�������'U�Z�G�	��wU���:<DȼA!���{�b�S��-��~�[����mZ"���!��p���ݱ����{�:�xe�h`���=��L{�9�G�Dn�G�;x� L�����}tFh�qYO�x}~o�nl����n��mه�_HU�2�b#� ��UN&�� �ܫ�@��^�ҳR/��H�{�~��u��]���@6?��U���e��n�(���m�������L�nsH��������F��`�0:U?�E�����]'�����9���K~d� �H�{w����p.�u���Ԇs�Jgc�o��=�*vV���Y��ʵǼ��f�Z~hC�K�NFvN;��K�{]fI��������){�����Ot�at΅�&�o��똗ӥ�(�6D�o�5U��GY�L6��aه楾���H�C5���Z|0��}��-ȝѧ�Q���٨�����:8}yvYy#$�[P��#C��z�F�f��s���<w6O�r�V�s"l���7f��vW�ltjP��m�m5�,k΁w�*7WWl��"�<��Յ�鰍�����A뭺�ΕGZ�5/�9r=�u␈8�����]t��)��7*ɪ3���Kg�l���@)ڶ�4�{�����@��:�/�~Ÿ�5�%�c��m=Ih��\3����D��F��Gķ�ܙ�))}@����������uN���Hy?lev��3Us�u��$��4�Q��
�Ɍ��Ļ��]n]M��m�nE��%�ۍ����!>~���jrg��h:���������}����+��1�C�_��b�L��7u�s5�+��t���a��I�_�f#���Q]�� �Kc�9w�����U�X��vtE���E!�n� 6����3.��PGQ�Fj��(vͳ�6�ZS�T���}�o��q
e��~�u&�mm�pǝ�U�i1��)_I�ە}�}aƝ�ߺy�����+�?ډbI�;9�>%f��&�)NHy3Ӂ���Š��zh 
��$��!��"��a��k��+��e�����3F���	�ۺD�0����٣����[gz�2dB�O�%����t��1���'LZnN�.�ݣϐ:}|cP���b#��W�S.r�r��Юc�#2�@���W��9�"b�1��j�o[I��p� ���{����T�S������S+*򆡛v�z�.m��!<Q!������9����%]���d�#)C��}��yck�k�\�5����d�b�r0"��˞��c��w��W�"�Y�0�+8:)SM���*7ܺ�n���A��e='�PV��/�'�����̿g��_��o.�N���O�X�a�m����O��vɐ�e��� ��d�E�f)�/�|����ۯ�Ł��8�.�V �{�rӲ���n��=��j�h`��w�� ��f��d�X��?2��:�s����y�
&8���:x'=�����M����"���^�2��g3��5#e$���c���n�3���s�ǈ��hR��K�]b�βRYiEE���'��}M�}P�2J�!�LU���X�|+�q�k�nˬ9�)W�=��GVy����e[�]8� *��!��n�m5Y)��;�	b��<a{�� �,6x��E�I�l@8�U��X
�R 7Y��a+h����]8%�°pi���,������)���f��v����G�n�e(�����[�p�#f��1����F�G-+,��4q0����h��ZΕ�<����up��wS��Q�>8G�4W0�́ �M؄K;�c�Ռ~�O���;-��ZKWU𣙶}�'!Q�0�v���aT�5�B����F��+�DUP
X��J:ڮ����E��i�gI�Z���s��H���I���(�z�Xi\8dx�Gm�n���)YsVm���@߮��V 	�+�.�� K{�YWCsЧ�*��b5�S2`wn?�~ѱ|��ڀ�5��	�g��4�z�Եt�������j����-�(:0�[J�m�m��m�sj��'�J�����N�$Ǥa6���QÒ$"�1o�P��x��g���ۿ1b��>�Ϸ�C��`�s�!M"�⬰�ZF�-!'��a6믑�%�69�y��U��P8��zh���G�3�"c^�#���kS���R���A��I�w�^�*��W����}�V���e��@"R�#�A�PpIΰ��1sP?\�r�f��c��û��ZA)I/1V�_s�Àr��z�}/ �a3 v����eNk3L`�*Zg�!�\@�#Y!^k�-�qOL�EIr5I޻��7�Yp��E��h�yawx�m���%�'i��\,���%agZ�|�\16|W�S�����
��,�\�*q���w��5�b���kӅĶ*����)�ьO|5��Ct ��L�O/�҂��lv��"��9D���!E��-.�QJ���S�g�,<_����W��DYۄ7R����]�8�_{*�|�"c�)'�V�|�nl|�M��ݢX��zg�t��Stn���K�[J&��Lw�
v�3�S8y4v��SR�K
���qZ�B����Q��^t�-�O)uK\n:_GU�����j�2`�ItQ�
��#Lؚ�֏�|�4$��T�Fx����y꫟V|�@wBf��}�Rq���ݨ�g�\�$>��O��5�]�~)����}�����U��M��j�HכCU���@�#NSi N�ߚ�y��"u�_��r�?�]��e�;��^K��nXs���r�.�g���q��1l�XC
h{�O��	���d�6����d�����[��& ,�%�QMM�`\}PT�*}L��^�?��ԗ�F�9��M�������}��3�6�$���~�Np�iv(��y����o�����Zz�9D�q�IlC�G�IM������;]��g+}�R_|R� ��uOH��&Ph�!i8ƫдh�s���h��$B+|]C�(+ S�gk����t���Fy%��ܳL(U�B`}=uPuA��c�N���G��Z�NN^��X[5	H�Z��,A^�m$FTPDO�ܙ+�a=r Wk&���sJ9��U�[�	\6h �������x������O��=��K^iX�r���/��6���E�O����s~�{��B��d�(��izj�BXA�y�#&�`yk�|7v/g��W9���&�!���QV@��k���©���AT�$�C
�K-�}��1穻��F�.7%h L�p�yW�OJ@e�	����Esɺ�k�9�LO����[�h�]�X�j�����V�u,7���!���;h��Ť�0���n�Po�<��c�7D��n�gxjɪ��v'�?��:��j2J���J;�xu�P�kIe�LZ
e�#C�H�aMI�4W�4�����E�d�'�;ڨg�:z�VFƝ�tb���׊ꁝ�KpW'���<๜�{�7�I"Fr^���!]�5��N �QPd�T�G&0��*�4�f��9���t�Ҧ+'!���`5�̼���W��r��>:b[�k�(�ȱy1ĭ{�����Ho��;��lVv$�DY���=#�S�=.6�Ff0�uQQ8ar�D�0��kA �A~�;-V��IZK�F�ɒ=�ei�s��G]��J$�qP>Rci\���ySI��EV�ȧ�5���l�����%m����	Dʖ2jix�&��Q;9:�G���v�v�*��d���(����-7"<+�������ɒ?�~�_$�7>��̋���Q��o}�I���q!�)a͹�吏t��1�O�ߋ��C��eE�_�ޘ�)�=<Oo�B���±�[J�n�fDVgϠ3� �F6�s��ȳ�P�x��S�t ���4Yz�-
�������\fG�����
CY+[9��ZS��ϧ��<�9�5��| n�ݺŹI���ۙ;�i�w��{T�TIgL'O�'cD�lr<c���&p�X;�vߝGh��8���y�;Q���ո�����F�5�A������V�l��ˀ%
+�j)Q���$��u"v����tc��A_�/:㾖�[�V�+��j��9b{u�sԅS�A�s[�y����]c0:B�G.4AI�����]�#x1�^��l�W)v���ۤ��$5$�/�$_���S�s��U��"�ZY7��A�j���ЫG&�z��-�~�p�E:<)��<i��
���h��'���d��G�4V����f؏Z�*��J�e-��o�a'BR� �� ��� K��l$��;����4g����}�lǸ�u��.�o���m(�S�xp��ŽT�uNvk@8��杇��q��¦�Ta&���� ���h����WsaG�k�����Z/A!z0J&�;���E�W��6�Z9�gm�aX�K9o7B�X�l�(�[��U��`I�%c���dG�g��7>4�ܫi	�|� �ul<7Zw�
£�^y\���z����f�E�LZY�8�-�0���k)V�._���Z��F4$��g��_��
P��2L���JY(��T�DJ���
í�5F��ݙ4ђ{!���tf���©l�������	UR� �O(+�*�o j�8Ǻ�b/MZs���u53纏H����)�Օ��#�U�u�E�R��m�W.[_D�Gq�X�w�}~�]��Ȟ!��B`���{��3�S�ˢ�CZ�j�"��O]�56k�*&�:�eDS����JY�R {	`Y7g�k望$D��^T��pI Ӣ�'�H2.���e�L���[A���'"�tF�,	��y2th�E��3�+o2��h`�.aO&G&�	Q�]��}7�#8�?���� 
�@Ap��P�:8в���ӲCPT���wU����.#Ѓ/x� �D�	�A��G���G��"�R��2p':ld�V��X�~�\�!�u:���֍�~RH�ܧ��Lڋ�����:�8�x����>5JA7nY��t�pr�m�k��p� "�	�Ke�s��6��֑z
Q���0Y�K%�9ݰX(W�c�!��Q1$t��]cv~��kZ�AI��+�e�(2Q��E(K�-�/i&S�/����i�o���G2$�����$��Y�w��<�m��s�4حP*q�l��Ĕ#m��࿕a$O��e��m3�wS=��K�:����v�#ц��(�����jbNX3�q���>Id�Ql��	1�k����h�a�٩�����00�v��6�X�Y���8^��V��35)�!�E�}7ٖ��<�48]7ϡ�%�1N_�4S�#C���d�I����o�7c!Z�Ll���З�:GɁ��l�|"�� ��?���G�R���e}F��oz��y�"v2��D�+2�(4�f��m'�'I�;����CdW���w�m]����=��9�����x�`��-L g��h�ڰ���᧘(�U��vZ��2L�I��:0K�<���N\�5�R���ī�2��|��c�:L�5퀜Ͷ�>�*��t�4@����U����AjG�͂2�&΂��Q~}J�ХqGٰ/`
�sqU�sǂ����R�PNĥ���dt_P,?w3V�����&�z�ﶴ���+���ޛx�偙��̊P�z��ݚt����E�X�1��~��C9�4�v�����c6L�6��0'�Z��f�E�n�Ӭ5G(<��$h��xǧH(�P�ZT�[Q;�G��?.	oE�U��Io�wJ�\��D�bW�o�+!YI4A�Z���'B/M�5b�X�ȯTr	�qm�ʁ��=�1*L�!z1�m��6H�T޽�b/l�IwM�*d�I���1a?�	Q�Lf����g=�y��q�G��=�����2L��G�p���P�
aՋ��}&ע]�~��F�6}��.1]^��4�"���B8 �G��帕`m�d�I�="�L�<e?hR�7�Ʈ���P�Z��>5���0Eyh�C��~�p�g*��Xj&�U����#x�H}D̏X���f��ե�����,��aI���Z�-���[�u��VG�'���&p�cK��Ji��7��N�f�)Oq��R���4�H�`<m�1/��K��^kh��$]kBdԽ^{�����C�:��D�&^���t����a��'~s�V��:�Ť��H��M �R^A�����"E;q5|�}C�]Ȇ-1n�M-����5�E�*�f��>
�W�o����u�r�$R>��E��,2j���r��+�_;�bS<s�e���mr�����Lχ�G�x��e�i���*m�Zĝ>_�\9�o��K�*�j��J
Cr����HO��}��4Щ����j�?w+������2��;�*�1A�O��f�����Li&�A�V}(c!�E�e��zZ� �jts��1%��ʨ!���QeU�.Hp��m��c�d����)A1lėhrxM�$���p�Wb�2H������.OJ����} '��ݭO�ar=I�S�K�'Mc��2��,�
zȞ����+1o<KInF�`uius�<����+F�ݳXkto��&��K���$Ӷ�R���y%��(���P8�Ѥ��C]��hQ>�P�w��STjQ�'ڿ,���ݑo�U=�����d�?�K�r�����^޼�&���L<�yZE�m^M������g@�t��g<�_�'��%�;X)��	��*0�L=��˱�0�����
$���n��fH��N��ے��F��������O!"�������`r���9ڊ���.�F޷E!z�8�`~-�Et��:����?V�Q�Έ5�%
jR�r��.�l@
�$-/�E�+��M^��^p`�Gj�)Ū7����	�2�0$Fw7��-ip����+��	e��	�,�0��;�a
ϛ�xz8�T��s�_��;?}��R��l��d�V#��CK���6H�~'$�x�	7���B��xK�)¡��3!��w&iz��rRы����аS������w8��)U�ĩ����jc4�]�uń�NT���fph�W��Uy��tS[��c,�Â�����_i�n���[� aH]�2�r&�z�������@,&��1g�<��P�]lێ���)��-XŘ�������8Ԓ,Fl;9�֥�p21&�_��ʍW��xM�ؕ�������V@-��%F�+{�K��%(k��2��3�{*e�r�$5S�9���y(��[N%�K�_VLibE!o[���ѠؒoKwM9�tzX��ƌ8w3���tC|��.�|�_	���C$ [\��2����}Wg�O,:��!w@���v�I��.�D`r.�0�xy��G�M���/�5�s�v`��tV�ź�����N�q!�G�ڻ����0�'AN�J�}K�c��������RI����<dk�{��pW:����h}E;SN"K��a#�&������[����}&@�r-�L�%Y��Dc�� )�a�e#�f�L��."�'�Z�~?����"�[yH��;ꤶ�V�(����^g���۔�bt=m�2���\����$�Rj����=Z�zՏ$���n2K���n~h�h���=��'���J�%X"��k�����i���x.W�]��6�U�
��7�w4�b��0~�h;������br�,��<tv�R8��d�O���f�����9>�Ѯ�N�L�UP��"a�]��ΐ2/��'�;�,b�D�#�&���$~+�I�Z��¦� �&Ϗ������Mm�@�TQ3���| {���d.k���a�@|p��\�/�=i��n�Gq�����|4�XA�6m�"G���C�d�����9�X�J�� /�I(P��V���Y�8���m�]������H��/~F���k�g7��	���V:)k����ʧ��;v��z�,|�"�	�y&��7���լ���Z��Tm����S]�7�"�d	�_�$?�v�[���Y���u���/l�r�P��lG<\U�zllW��E��Y�y�Y8��QkTW����pAJw�<ic��d�
��|NeD]�)����B���ýa�.�����N|�EJuF�Z�C�0��
տ���{�C�=����n�ñMӓ/	��g��������f ��6@Z�8*EV�C�Y���G��A˗sq���vA,
��q�L���&7Kuh�v�p��;��Y���'Y鏛ê��#ԛ��|��**Q���ɉv
%�ܳ�S�Ҥ���HB�`�H� ��,��D`�'��k�g��G�h�2�2>� 1�Γ���hS���u��}�W+���*�h��f�T�cYw���P��D�.�6�_��̑�`��`qȽ��ft�] ��2�9���MQ(H�ā�u�<G%7ٴ�]K-�؄�*Bu�qoK��"!�f�dK~�OT�Y��|�b�o�k臡:��nBS�.��;�9���ۼuj;�xP! �ܘI�de�dރL(7���`���"��k���fdz��A�F#��~�,����G�=ʛ��#f�΁Fz.%+��ȳ��BUP�GƾcyԮ'9j�KQ�j폆����d;x^?+뽶5i���q~��|�~�)uͷ��A�� ����'�1Ȁj)��@Q���ڄqB��_H�о��f�����s��YYH��s���!���?Ta�Z���(m��/$S����e�47^qs��D�f5R��o��L�P�=��}��:s<_SE�"C>��L�[����S��;%�o�eUR'��P
��XD�G=�j��q�~��d���-n���v2���|�~q�v-�_�Q��$>\�1�o�ALዳŦ7����A �����BX�:T7fz�`�C>��
k�֜�ɪc0�BxW��W�D��9@�bL]=���,}d�AE%TئH[��W�<yK�D���g��喚$X�_��T/	�a��{�5*l�tn��"{+ކ�qq���fit���$o����;����p9%!���XVP2�ÏJ�v���X"�@ �7v�s�c+ے<�fDN�V�X�Sl7<�H�/��k�Omi0�gk����d3ڒ�\��kA�C��T�P���x��Q��ޕ�Ѧ���5D��q��a}+;���AT�Y���Ɲ���b��-�y�} ��Y��8/%�D��n�Vg��nY���}V%9�C����b�r�"�\��ި���v��:'��WW��\1����-o]��G�)r���8y4K^�3���#yDM�|w֩N[O��7gG� �W�GB�;���d~z;1��^�Z���zX�1��e�Ln53t���� �����*��䤗8U"ut�gJP�Tn�u�00�T��)��!��Ɩ8 6�<Q���J�7��n>�77�j�ٺ߃��x�V;1 %�� �4�e��Y� \N(\�Lw���'�+	��C:��pO���.PYuZ�����m�y\;�����X�ײ��-��N9�k� �W �)��`|9(������"χZt�AT(7b�K�Q��K�LT"��Ag�9���1�o,��׍��LR�O�y*�R&�.v\Ҕ�P�r �1�?z7�[G����mn�,X�\���Nt�.{fY��Ht�?��s蘭��YF��O��<B�$9�6%"$!�Ke3T��Յ8�}��>��n��W�v��$�('a6�i0�hq�y������n����I�.j�!֓I�i};�~j�J�v�{��bX5�g��l�*e�O@�xk�"�Mb�Cv����烫� ݦ�:����2� ֟k_����w"~��e2���P�t���9�>� �qT&n 4P�?�FtF�S��N�#��Ϳ��f�1��(��4�����,5��	z @����m�3���� �I�T94�*nK'vh�s�vmPV�2�	j\v��g ��:l�>rN�V���K�H��v��$��|"N�Xݜ�E�B��/��[�)u�b��-� �r���]�8pC�1�hVL��+�*ؽM��f��&2�g���k��j�|,���F�,o'�WF��Bdv����E�\qA�
*˸��oP�*��k]C���7�6O��G�y�6���_�*���!����=#U����+=p+c���f�o����릓�͜�?~.;���PK�;3�����6���jB�T^6�a#��P#��`�,���P�����41�T0�w��lMvPq#}��k�2��� �v�bT���ĵp ����u9&O�?O��՛mGz�nh�U���:fe���bw�7(��i,.v�*�^���~	��4��|���M��B�T�})fC�5�����Dwl�}��"->����i�?�jZG}��M��У��Xbc�җq/#��0 򢛩%�r?o����7���O������0���b�*����M���A�G�1�Aj�mr�,w��?���T�Qʖ\pu�&˴Px˕���xV�?����;�	��=f�y��W/�L��A6��3Z�f��3�a��0���+ԋ�W�^)�M��Ef��ӫzai6,5�o���oV��N�d�>M=�El��zh�`�+�-�1@���k��w�.�_�P捹��@$��c8ae��F[��Q(gnj">�,�s�x�L`�师��Nw	����K�0UB�?6K�� �_gニ��&�2m�����>�WXS����.R�}L,w���
7�#�0����|�jF��SB���f�ik�觕����G߀������s�m���RI7@3�<��]��:!��,����W=�)%v� ��Ygu��k<��)R��bE�����A���p�P�� ����D��j��e�����e�:vGp���\�~ƂS3�q�*Ζ7&����7I�ފ�lF�pE1JQ� �j>G/j�6w�������F��爠�p�q�!k�
����4�}ޏNk��;'�|�
z����|x�6#W	�!=�ndx���B��՞3ۡ�2K3�?fX�&~dV�ss��g%�:�Ab�g��H�J��p{\qwGL/��q_�߹{s���.�s�P!��hp9�p4���LV1��>�Q��qx��y9J�@�6sYb̶�g�(@@J+��é�OI����rq�&y�+4�D��\,����}���l���0�5�H�% ֩�K�xC�B	�B���+��؊M���#����!��"�����v# /I8��������aP�4	��m�}�aSv�R�F=;PMz�6��š�����?&:�3\�m��B��� _�����X�gA�|B�ߧ,WJt�+'?`�R��u}p
�Y�Rڑ��g�k�3_��^� �����xO4{u*��5 ������<��}YX�ڋ)!�|8}O�.hy�q��"gu��׽(hN��^�t����$�����M��y��,[�4�m��NKhHZ�:K(l�J��y��w3,��G\�N�	_0���Ӈ�uv�Hx���d0Յ�V���<��h1S�.
���N�맮�x~���҉���W���m	������խ�)}p�.�k�K�*�p��ł3�Uw,�u��'�uR�(I��:��.*�p�����K�X��u���
��7k���	M��0�ua�G���8Z����RC�nh,� ��/���"p$���D��*�K6�R�`Y��FԶp:�-�}�.)0�'����{G+,� ���p��)G>�R��|-5_�[��4֜�,U����GL×���t��&��;ǥ�=�Jy~E3SO�R�p�/# 3�L�#��B��ϊ�*������z��\��o����ցt���p��3"Ǡ����}�ō����,��	�[�F�$�WF[��_��V���q�ǀII�Z� {� ��+�)���pl�6�b�
�������TJY�-�A���T��\���nHc�Ⱦ.��ط��p^�E�1���)R_�\�q�r�^ f<��d���k�7�Z��ZU[�-�)bt"v���<O��S�jvKj�"�%b܀�*��p���y)�Y��S;5��%^Dx�.-�z�_g{�:`'/�"�9" �� 纑���ڳ}H�
q��̕bp�RÞ��吆�u��	t|�` �Vs�8o��i�W%�ځׯ�����V�����I28�5��:um{
�W1���#@,5�����@���s�*�P��u�^�Z�Ɩ�l�q�-����N%�K�� ZĽ�W}�8B
�T1I^;(��t����D��K�m�D�0�� ��U{S�w����e�3��/*=]%K���M���ə{�\�e����EӃ��hu��N�7���+t���t������!(��%�
��l��f*�I��ke�(93�u�,��l29?`{5����]�tGt�����]k$���x����I�e�
n��������~)�L�d>��Z��g�S���D[t/�H1_�8{�:�#�W�K
�E�A���dD���W�.{��Lŧ�1�����l(w���f��O�B��7�SȔ֦�
5� ɴ������I� �oP)A}�l�.y�_c���>?�7�|Q�W�s;��X!Sb
0{˃,�?��P�:�6G% p>
�{!^���Y(���bEw،k2���wɗ�<b��� �e$��2�4 ��пc[(_�]�����\l�%�I���+��Z��A�xOv��Vn�3`?ˏ'����O�����H��R�ӯ�ߒ�}�9jf�z�ye�Y�͉򊅑�;*Xt��9��J��Z��q��=��I�?��D�l���p���ã�]�Վ��>��~hsG��{�,�A��?vdnJ����c<��4����C�=9��\,[�5�7��ۖ%?�{�)ʏ~|��u�i�LS�0�N+NQ���nUvق}L싻���Fq ���,{��:���Q"Z@T~��B�4��|�a
 ��:�׽�n��6��$�aqe ����($rv(�ށ'����q�W��/>;�eB/���0�@�G���0j<ݧ�q�&u�^���u�
�{�͙V��q�r�k`/>��U}8�i�S�[JR���i1���h"8�9��d9� ��9_R����|q`�R���oJW�$����U�%�8TM��<j�w�}ǉ���K��2�D7��z *jS������`���� mx�@ۗ��Z�Ɵ�u?.g�g��8�5t�|(��k�D�]�:�Zcފ��/a�%m3%��`��@?OJ&_�rMz���Zm0�JY���h D��WBp���3�b�bTjt��f/o>�z�iDV�42�y^�Ԝ@_5�L>���Eq��9@�94+��5�(p�����I��v��;�W�W=�8�a���T�\���#���0�ݖȣ�O��%;���f�h�ԓu�O��~���>��i��n�D���nE�R}0�浴���0g[�׬�9�0U*�e�?�a¼ߝ$�O�W2�np/9.Ev�����[&�����Lm7�0��;�FCS�f(�vL��uPS(�@���is�Se��#[Q����
��1r	�(	�a2<�edw�;:��w�����݃�s��+�9џTd]�7Y4N�a';\�4[��j�w���#� ���e�N�M�~�7�R�}v�ʆZ������B��ؠ���&@|����E�1(M�uG7	��i𠩗=�� ��7sX���$���(��k#Ϯ@YF��Tm7�`��>%�J��PJl�Fmo5���!��4�W�ћC�B�����k����2Wl)�8��j�G,m�h��*E�#d�+ZD_g�c����g$d��ѵ�=M��̙�1
�ϼ��.E�&=vzِ�ȳЮ	�����c�)g�,O�|�Ų��u$wH!\�_����8K��!/nR�8�d8<�gN�wm�S�)����(� ������e��3�=
Uu��<1���U<�G=連	�z##H��չ��(�{��� ��W��a�n�`U"k&{��QGBQ�W8K���v��ؕͶ�s����FR��0����������QX���n,���XM�)6�F&H\Y�q�]M|��B�q��%��/��ح��Ƣ<�)c1n2����$����c��� �}�`C�����)���������E0-�J��&a���~�i�J+>h��P�q1��1�'����ҩ���d:*�Ⱦ��#�_�E��w����� -�� b��%�>� |�_V1'�;GKF0�\j�*�+]�y�P}������!#ʵ��cF�.�v�ѵ'%�e���艀F�@�P��6�ٯw�L��#��D��&`~h�+2|ok�K� ����u�n�ӎ��o�D��O��7�T�=��߱�S7w`�(RL�p�P��4�ށK�M1�9�O�.o��s�SqR�S�t�]��.`�Y�
E�o�6$������1�=QV޲EQ�P��9��_��5u�x+�gsU1�����|�2���wd�-D�y;���vBzM�?��FU6�D���>Q8m�M;uuS�A� ]?�
��ߛ��E^A�θ�(�Ks3���?�WA
E��w���u�	Ϫ"��heB�:=�E���R c"Z�9��?�bb�R�l[q�Q�<�?�ֆ��ʻ^l��*_���~6Qy��B��h��*qZ>� c�  7�-N�z�cϓ���u~���^v�C�A�@2f˴������i�5�L��V�*�����!��1O,�+m�?׳��+o��;��0ڑZ2K��12������z��j�^ɦ��,;R�Ϗ�
z�bu����ŮK�^N�}��:Xq�J.�㶌�'	)o��ڎ�rJ!�gp�K�HDt#F/�d�yx0�t�>���d�|�Pm��8}��Z0��u��X ���f$�c��y���m飱�[�3I���K�������ΥQ��>5� t7�㷷��+���� ��No��4R�\y%�t�i���M��R|��Ť�5\����=�n��|��.��Ri�??�x��!�(Z+˒v�D
��WОJi��}Y��u!P[������6���V}s��	�?����m��[��2�J� �"{�|��%�.��-�0�8eLSrxH�� ;n/y}De
H�=`�=Qi&�Ó�V���N��@"�^��Wf~�+Hi0.XA���Q޿���y�g�%4p�s��Q%��S^%d�aY��(�&p읁���X��K"�A�O��R%6N�RCZv�<���X�q���5�G.k�'�S�+,qS�}">O��,�wV�jJ��x�H���E��Y�u�R,��c�aT�(��
|i��!ܰU����Eh����=0Xr� �@F}j�A��F��&���&9&k�k-��!��kr͞�5���8H��%�ޙWf J�b�*ܝ����$���w��̾��ړT���f���5�m����YGN� H���n!r"��L�d��J�]t�T%�o�g&�8�&��]�:<��^�0������l��*��g�_�NU�L� 
_H+����l�.��2y_M��4��vj<��E��$�P�.P��޾�����(n�.*/:����l��wO���`�i\�|oMQ� �r���(�w��rX}��r�Dl�N�E~�e�?o<k�;*a]nW��2��v�}gU[^b_˅��I��� �?qW꪿�w�q�q8��kF52�U��b�!lm��?���d��L̀�_����� M��<L\}������#'T<��O���A�c9Q�0Z��w#�D���*AP~�ZH���oa�(1�<17�6�z��
�/�=��1	�cZ�r^㵣��?��S�7F�h]d�WQ��&�Wn2mx�\��?W���t/�@��n���ҾuY������B��e"�	��a��=v]�'A��w]?�$�2Y;V�� �0�J|��ȕ�a�+ `�?�vq2mk�����?|��녛�,:�O���$��6$+�{��+ofy�>q���ɥ~O�����(a��5�mJ���5�P{n��m�@b���d��]���*��BO���̃&�C9�/�0��d|�/\��=F�$l���E�:��jѩl6kr#���W��L!����7��ת���^�Sn�/�L���V�4����e�;B��4�0 ����)oW�����i;�G�Z����t` <�������x��W�pqܗ͘�e���d�)Յ�G�Ƚ����wk��DcPO�)�]�b3���$䬿|��kX�L�;)����S8����C&{Ӟ����擛[��};(�?7-�H��l�ި���=C��
�ڗ3*?R��mn��va�S�oK���z��$� J%\�$��w�� %��u �I��J���d9�+!�����c��5��ID_R�f2H�Uf�+� �@z���J�A��D�*�Q݌��U#�\�4Ӿ���׎m��o�:?��v�k��GR:~����[��=.0T��QQ'��;�gq����d'�̲����}�YÍ�������Twp&:��ſ��0,9�p\@W��鶢�R��~�:%Sα�*bd<tЄ��ŭc�P%����FV��q�� ��Bܡ$p��~j�h��j"��/p��ڑ���v�	]�'�6�I���T�����
�!So�&M0�f�Y��!o�>�!��p���1��þ�Mx�O�Mi�cGdK�|)���a	��):�U��gT���� �� ����xێ��TH�z[=V��U��b!AH����+	}<�b:6�ĕ�� ����a3���k�	ʗ����X�>n�ۓ�LC��l_86?��S!s|��jm�,Ж�57Ȭ�k���g:q �t�E��\r��q����i<d��S�+ﵸ�Q�*�"���Z|��!p_$� U���<H6��(���O���7�=��
��	���Sy�ٍ����,g�׼i���R��0=ʋI��֐2� ��cJ#���>��\�nQ=jm8��U��wR�{)[*)JA+t[O�n�dp
a�͈����H�1`�A��rZ�`���C�B������P�+=�ɇ�$G-��J�VG�kd�[�N�@B�b�&l�*������1��[��H�u��ؗ���QaZ��N�b��l��,
������Ğ��+��N7���Dܟ��Pm�hZ����yC���9׌����F$��Dl��bv>�"滄*b�m N����P8b���'��=�N[BÏA?��|KȠNj7��<�E�w�-��6l��X���٩+�M�Kť �7]�5��?�2�|�J/�|��"��DeaAM�YvB�;��?�3wǨ�r�
-ީu0M^�C6�o;W��I����OӜu��1�Tf��x�"U��=����⹨�:�۬�s?�mS�ۻ�+9W�qP��M�/��ki��mM�b�܏��(����Kn�Z�|�	����ι�����,:�܁����Lt��探$�Sc D���>��h9I~N�������y�����PD%m"�>+��\��� �
��!$��%�\�B�&���W�z�K2���� ������dh�yS\�aZ3���</���M�`�z�	���{O��t]84��=�����(�)�O��V:8��ܻ?5n����>�2 �K�4���c$�5@"��i͔������Q[��"U�)r v�o{3��&��+�rmӮEL{#�<�f�n��xF�D��1�9' � � dYFA��e���b֒TE?��D/0]"r1h%�̺8����K�)b�+�����X�S��#tH��<�،��@�2h3���1	X_��B\�lj�f�h��7.�̓�w�uݪ�̨0<�^�=�I���Ŵ$>GG�HnC�_�(������P���p�a� H�8s.����#�k ����&p9D.D��F��qOg2�oݠ��řt�T6s
�8lyf��P�G�����T�}�ǭ3�7A.���r
�z�n��?�OV��c1�DuI�t}��~(������}ݳ���j�v���^���^���|�4#����T�XG, ������~b�9��6 M4�i���z�(��0��a9�ĭ(��s��v��0�D�n|�	B�j[3[�( ʸ7��-�]�'�)��K��$$��!���_-N�L������/�`-��>&cS����wf����$k2��>1=,���(���i�큮�H��}0L��i��Z�sMR���Y����g�k㫅$u�ݓӆz�w��\��|E���(�'�k��hk7Q[N���^���+�����?�U��$���?��d�p'jyN7���q��C���/�_�}�pm\.�8N��I;_%ۚͰ %�W��#J
��'C�%}�oT��1�[�K�LV�^�2���iߦ�c��bV1��������!\.��Y,s�k�Ihڇ"�[�!������^�p���K�F+�N.��o�}p5Vhѵ8�N);�p��u�=�^8���C o��e3FS�׉b��ȍ�mL�7���y�@��N�, ���9��_�sېS�3�kѣ̄�K�O{�yO&@H�� �R��ѽr���\OAzSp?�)�qX]�a'��n�[x�¬���\���W�����vH2ny��d�cJ�a)��즢�Jܟge�䔣J�a�tj{Cw����X�4�҉B{|LLI`�|�ХvV�S#�]I��F��L�<㉦�W���vȚ/U9Ap�T��7�Ԥ���,Zk�U4�k>A��G�X��r���o�)Fb�O�4�jH���P8���v)$����.����������,�'�2���P�\s2y�qjt
,C�Y ��&'O����z#쭪�;������&�6���?sdv��[|��<o��ԗ��R:�*� �@Ģ��]�^,
����
�u�b����	��ڽ���_���{�帘Ѽo.ځ�$�ŻN�Nl0�7�_,�ax���=|��T ������w�g��c�*���G�G�񍟱?:X�{�Ֆ��y��ŷ����9��|eq@Q�gH���]2b�ȣ��HM�:��3֞A��ܬ������!�s��H�4<��#���ֵe����{���t)�h�߅�vξl1�no����Ŕ�S�i��Z�k���1:O�wB߭��!�U]���i�0���L�.'�p��FJ'�|�!(+"��{�J�>&<|�X���o�1;��	�#���ڽ�p�U��Y��pS�:��=���ð߻C�Y�G�" ��^��+�	Y���(;6X����z} ٗ�h��[��{1:*������\��~�jل\����aΗ��@�f�}:��X!#�Q���5Q�Gإ�Gq�)g���S]�$l�Uu����%�8*#���,Y��Y�ނ���
[��,��f�(���1��JϹm;[��侴IQy"^�#�*��׊�@f�b�,uZP�� K�!u�)3gE�������Mum!�4���<:V?xlz���2�2����W�����d��k-\G(�^��O6W�^l�6�+!e���'�X�����*��@([\a_VxM��褱�H^^j��������o3���^?wY]���4��af\y�N���e�i���B?
x#~o97�����'y"���Rl�Қ��=в�,�n|sM�f��1e8Y�N�#�hT����;~��	�jt;�f�z�β�c���/���Je�{/޿���!@��H�ه�m�}��,rF�(lR��3�9�I�DcF�+�>�Y�#�Ƙ6�Ǐ��@v��v!�K�|cV��4Th�s*췂uvZ�l���1Q�,m�T�q�#.N�]�����C�:X�]es�4%Z����flv)φ�LP��CM�0�Ud��]��Jh��s�!'F��
,�=��<c*h�A�oq6��u<� �|
����Z����E[�v�?gxK㐬`�F�L�ו�X0����c&��dS�c0F�z��K�ۻ���K����o	����#?�{I����2@��p[���o}@:S��Y�>z�`HW�]ڧ6˘͡��R>����_��>n2�p��mJ��CD��uC���2z�f���k�_�E2η�#��R���⍵��"�i/yܴ�{���0#���D\y3���M�G��fK�j��S�����?�P8Aw0�w,7�1��	����ўJ�߈� ���cM)�NM�c|$��Mɿ��^�PɆ��;���h ��t鍍��22�Fb�*�W��]8v'��,r昴��Ihlc�����h�|������7���^9GM�Z�U���a���%�0;�2���RF 0��7�� �%%�E��~�O봧�C�jqR?%^�yB�^¾�B[>pO��:=����$1�|��=
�QQ���%4x�(WB%޾��y���xEŞ9G����D��<���'[�X���߭h88(Dc�`-�K�4�~kJՕ���ج�_��k s�T[����9j��g*�dF��"Ŋ%�B�7��*쏢8G4�HA��E��y��
��f�y@�ԭ���Yxhv ��=�?14<��.*��J�<	��q�������b8 �G�?�p57�Y��{�0O'�N}c�R7p TR?.�6W;�J91r9�7gªB�5���J��`��D��9��,���q�'D��7|��(�E���YrWN�g�Ǘ��^!�X-����./��ฒ^�΃$x�:E~[A�ұ���h-�9	:ÌM`�uZE��G�������r��q�+��bI�c��X��P�LQ5p���ފ�X.�����&���&ƚ�	�{��IKO�M�ð"���,N�J�����Ӆ���Z=����t�O9�m�Ќ,�͂�#�-��ZRQ�D�)ň�
QUEU+ڮ�I��y�.�?��4����xzJ���A��PG�.����޺���O�Uz'[���_1�bج��u&�uW1�ՓU�(���S��_���%b��q]�������d"gPMm�0��/���4�� �wMqD8��Yf�l��i�~ �����T��^�h��ݽ����d������Ĵ`X��(�ž����x��\��X�F�shd����� �w>6E�.�n7��Xt�\JGݙ{3/Цp�b������ҧK#�J�Eer�=��ƪkӊkQ�n��_����N�}�Pw��g�i�Dܕ����L��Y�����n��"d��/[wֆ�_�`=-h�Ҏ�����/���i{�@����26�pG}��V�	�h�s��H������(7�LW���y�C0л���Gt�;RU�� t��������ʗ�B(���o�C��9͈�����St�ޞ�E{@���]��K=��J��S�R�Y0�� P[�?�a�M�	�X��$3<�X��	Aw?���e$ƲMP��K`̹&��%)��Lk*�\IiAU���<�F�����]nـZ�}�^nX��l���Ê�Ԍ�!̛�&<�
௶�$���W�2�*2̞�#�0�WՋ�w���k���@�Kx�A ����&y�i4f]��~_���B�#+��{�%}m��w�ë嫢Zv����j�P��|�\�>�*��]�V���+���N��,-\�Ω�-q\l{}��ɞ� �ұ���p���.>�?>��b4'��%!�;���M=Й�+�)�KZ��;t(2r�;r/sn�����hZ(�������F6�=$��)X���հ�S?1����Y���7�s���,ָV�<�T�/%uW�q���렡��E�cTD1�&.Wb�Y"Un��D�����x0����=��b��� _Y��b��]�TT��>C�X��Yf&A�b�GIcΗC��u�[���j���4���4,~���Ӥv�s�Γ���fM�����\�s����xw��%;��t��>b;�L_��\Z(�Sl��6SW�g�~������	���>����=�&a؛
%�vdڻ���{�כ�����SD��!�}\d5q<�����Vl���Ǘ���	}�B�5�����xq6�gg�*�������p�,3Ӌ��s��%�����^�,ߡ0����o���h�a�5j����h�����䞬/5Y�՛��t�	���������� �d��zP�I�%Θ쯟�0?KOTG��\m�aEB(�nO ���`S)�Z[Y���=w����%>5�u]y������ 7X�&�+n�ivkhA4�=k�ij*�=�c,�6�9�v8� ��ĭ�0����Q`y�{�ζ�F�v��I�w�I���45P�I����o4�+=U��a��|;A�G�������戫�h�J9w7(�
��3,w7�u����3].Z�y߀�&�wݗ�?�|�d���9	?�͊�L�{��	�}��=��J����6���E���;�&�:o�[W�Ғ�i�-����_�Q� ����۴�F��Lj���Oq�F�D�n;i*��m2��j0��6��H�-���$P�}�m���?�����%؃��_�8Hߝ̩3��*R�+r�	�.��آ�ɋ)����|�{��mQ=f'��ʽ�:����9o�ľӧןn��uQ_g���^�L��{t� Ғ@��F�m\_e=^� ʉ�hĴ� ė���V����w��U�E��wF�\�{_ &s���͖+��.v7wK�0�|.*���$y��I/�b�#�PBb<��W�w	;$�n��郀��������)_ �3����Hj��j�� =8�S�I���EU@�}�|�F��}�+>6,���!�_3�Dk�����VMIBꝿ����-�,�;�T��W��ޕj��c�#�
�A�[2p@�$����#09���sw�6Y1] Q�C�q���/�Ue~Ń~�uq}��7/Y �0z�-l[�}��WVS\�fs2��mɞ�p'��>��v2q�S�w"��nn�D=� '\��|�W��q�����&��wD,!�H�$6'�!�m���RjH(wB���I1+I5��ddMO �I�f���}���>W���8ݰ};']gH�S\z��] �Hu�{��[k����V��K�\�*
| �1� x�ւ� ��S���CI�(ǋa0�s�,�w�c�7��+/���32w81��a�&@�N����2�1}29���\8{|��{�K�9)���P�|�1�� N&�2ׁ13ӯ�ՊV�8}S��3�6 �U| 3��&i0�e��"���y1���$���1ޡ�C��Հ���{� �HO�������2�*}���`C�:Yh�σ]�����F����{��!�������,�T�:d�:g�d&G1c����ފJ��*�P�R%�P{�X�k��!��?�N>�n����2�gHxqm(q�@��1,l:�r�c��5bM�è:�{ �MY=������S)��L�^�u�-��8T]
oƩW�"��)�N�JP3�y(ŐQ�iKA����/����K^���P�n�`X~w����( �DG;�4��;1��ڃ��Q�3f�i�٣9���Ƃ.�Z0��1��ߝ�ʩ��dd�O���k�ҥ��my�7#ɹ/�� FN�[�ص����O�ۉ��epg߸8��OAIK���I�[F�a��AB�Rh�%F��@��;eR�?�W�m������� r�}@�C�x�d��<��*�\��8��eW����H��U�(;`���WZ�x1���% �,~"bvϲ��6��rd_>��y���o{���W.�l=.e�is]��k	�t�Oе&�>.��r�
�$�N ��#�[�KZ2l��߻�8�n�h��>�Oef6�����6־�3���-#�?q����2�6��$��A� =V��z��Pw�h�(�9ۏ/4�Q)d��͂>��/���!A���)���\�c��/@���������kL����7ˤ�5u�@Ԗj ��Ëv_�x�����u�:�~X%����Iz<�2�=W(#~<6���g�*�U�i/yh�|֓u��؂�-?�/R��q�)���s�r���5t�Rյuc$*����A���p����o�#�޹�]�/4��8q'_uό��%.�;@��B3�����
-�X���e�����	�l��d�O��j�����Y[EMM\v�N��������$N�
)+�>@>+�R<���ۅ(���R�-%��;��8R..��/�On�SkAk�#4�����׹��*>��s���3<$3��'k85�׭�U�/����k��)��euF��*���@v��5��<�B�\K�Ԇ��UÖr5�9��O>��4%)x���]�8�ʀN�uǓ����XhD�)�r��T[N�D�U���`��\�J�����p2[N0n2"�F��f/��l|ptd��DMH�z�0K�6S����R���>��E�?�j���	��$r�fҗ��9Ѯ5t#���Q{x(����˨Scoj��7ͅ׉"
�S�*2WK�4;����N�����O��,Qg��uϿ�aЏSB���_?��XX:}4����bOVAK
�i�����'��MI0$�T���)N3�Vg���l�rƆ��O'�|ҀDB��,���Uz��1LD0�6q�2��TR�R�*�~����M[,5	��gQ����Pd!b�L��*-`6lW����h[O�#��Ǣە£k<�$(�f�a�M�ހ�Poj��_��?M�]Oa>��%��^���MwDt
��X�2'y���$ɂ�PmPc��Q'�)Ɏse�^��\S�}&���f=����e; ��_��>��2F��/oo�M���Y0���56��.�Y����2
T�X�����A[k���2�:�a*Ci�,I��*;[)��^�si���^��&�̴nٶy�-��$���=�fx�0ű�"Ƀ�;?~u��//�8����I���-���c�����ޠ��R�%k!rQ.-unh���t�0�*���l��B�=0sɧ�~�&g)���p.XV��3L|�4�������R7����n����i�]���7��\:Z��3v+�9d� �f�#�O���,�}���$S�t >��.�4m.^�Vj�?N�0��+I�t&/1-�݆����DUs.�x� 0k�(�5��z����v�Sʫ��j� ��tc"b��֖��A���9
I� ����2i��׏"��� e��8�Oԥؤ��c��z#m.�<���a7�d�	���EiO�GD&�I��>,i����n��8�7�}��B�a9@�<�����$J�
,��T���9&�#��^�_Fۨ\�^lE�KZ�w�v�6Q��cB����Kk�?'�����=rfV*)|�,w����I��K/�3ɫ���	��;���qW��_�z ��\��\o�`�d��h^���LB�̢�4+h�)��m�fw?��2��A%���B[�*�x)�3t�Q�{'�v(�Ni���ؾGT)S���?S���О�^����t�E�ۚRc ��sr,�A]�Az�Z���AK� �H��Q�(NEJ��Ƃ�Ep�{VS_x���~F&��o����	<,n:�T���O����Q֩�������N����3W�?XF��;��1ޞ��6$�9f�p�����/A��ɑ������"&�̾.��՘����L�xR4;4����`����/�Aofc� �$�	&�X�q)�Ct��1�Sg3@e��uN�~@��5���\�͛j��3K�t��R`5��o$��XY�m>���������+"E{O�淆'���tZ:m���BR(a�=�hɡ]a���'��b���C�>]��m�L�g�Q��2�l�Վ����9�
��i��iw�� ������XX�; ��2�@[�]��*�W>Hw�qͱ��a4�ҵnxJ&ɘ�J1���K���tD�Ƀ�]�J)Ie��d�n���؍��}x�/~�Ȱ�/��p.�T�sJ3�ޢ��Z�cQ�`�86�����?삲~+�%�C��� �f�$�'���i��#�wr����I�$�gʗLe�����-A�h�Kȷ��V;�2�O�pٍ��<�
�0֧��9�fG�Z�T�̀L#㪄� p�0���Y����ߦӮtF��$����F���d�(�ȍX���,&&����ѓq2e(��y�=o n������ /���J�@��p�N��8 �q�?��Xxp�)��z�z�Q��s�Ǚr~�b/�;��"�ܳ��CME��hh��L8m!zq�k�R���%e ���t�Fra.{,T��u�a�z`��+	�cG�
ɦ�v{i�&�p��i��Ъ�
� ��l�4[��
�?�s���Ɨ�d����ې�M�I4l��V�q�A4ׂH��X%��Bp��	E���(9�ŏ����/`~<��u��Z�n�Z���M%�c���z������Xמ
�4�xa������������z�!Es [z�<�D0��-����U���fi����Oc�k��w)�nnCc�}?�����e>�n�WX�؍"F��b��W�sx�vZ0����@$�8�%�/;֐y���8���[e��y��p���v,�SJi���d�g�V������)�j�?���ذ�`Jo�Ly���H-���V<�70���$��{f1�|e]3�T��YHܗ% �#�*��	"�n܌)n�#�JF����i���.h�Oї�i~K�]Kk�ĳO�4�E��ݺ�犘[���J>�L�H7(�w}u8��4�<�b1|�$X���/�����U)� ���7%�HqΫ8�����H��m#��+�?��efKt*d�uz�ܧ�6C�ۓ�O�J��u	�k�;Ȭ`�\�W!��5���D����-�����4M̧7YPbgޚ�∠�@U).��q�u]
OM�3h26�5�y���|:]�`N,�(!A��B^;A[�F��ո���:����vp�f�HM�ePMiT���߰`��ggvL!f�l�q G7��؏�*GR�Lne&�d�Ʒ�Y>�}����D9�
bz�����Sf�b]ȋIKA����<�^H����B�Ӏ(����bq�������z�SJ;�h��if��*qhl�6`?
ơ��y��b�(�%_�@��M-o��1��p	&�!5l�X�DU�n����8ه�=��}mrZCIgߔ���4�[O�+�9��0
�C=�ME-��),�����T���t��Tf��qɟ�y��E������7���<ޔ�Z�h1k�8�:���~Ֆ�G�8	L�¡m^|R!E���[����Qƕ�����$���B��¤���EW��	ߒU�JҶ�5��&sA\�o�g�$_G���A3K|����t�O|Ff��幩I_�x�/���0��	u����|A}���9-��+Xu�B
W	Ҿ�1{V�	�BX��W���H ��G���gp�};*��HD�	�cĶyL�&]��qz-����Q���8��3�	G+4�ڲ[��M~c5ӳ8�H�c;���$A����iK�B������9�,���-�k�� GZ�¥ ����k����IŐx�86�>����?�<�ҁ���$�f��8"bl��n
#�y�� �rkO8|>8�G��S<eiQQ	�
uj�r����dXs���Y	w��xa�7iY��nadrqy��O\F$P�P�?�hhĠ�/'L7�Ͳ�q\��=���:*��yuG�1b�e/T��0C�n�t�z�4�_��`%�muˤK���	%j�d~�c� ]=f֞Tf�T;���(zK����jQ�ɒQ�z�k�Q�q9{�rA���!�>��TƳ�?7y�����.(h������R���A���#�*PU���Ӏ�_��"D���~�郒���ĭ/Ý/��h�d�����l����f�-��h@��Iu^�rE��L�b&.���.�*�Y�G!�%�1Ӱ¢#ۚ! l:o��=qo��nl�7(����/G+�Q����*�gu�}\x�"7=-u�~\Ƽ(�'w)��~�j6
��ݷ�I�8��8+�o� 9�
��I� �lӡ����T�SG�韪r����=X��b��;*�Q �O��G�7H\�!?qKS��&*�
s z =�����g����fI��=�?�n�.�]'!u4��� �MV,�X�2�	V�l�����I��c�)�[���ES ���\���~	'�w��w�*zsC!���:�LE`n��DST�������R�?�����e%]z�]�K�+�N�H�>�4��q�J��[L�;Y��m��� [v�Y<��"��ȹ�]`����q�3��i.Җ��37 S�W"���͉<���e���:��M��-U7٩�:���`T�+F(�� �np�툀<�j3Q�e!�[���X����ٔ�RY��͖�}� �N���S�_��ݝ���g~���z��k�� B��
gZ"|y�.C�`��J����{30��1o���c����$t�w�!R���8tB2���\�9��]�c����D�k���N��*fl[����S�.Wm^�#�gr�Ĭ�(mk����<]�@r�q��P� �IV%���Z�l�PoG��?�!8L�/�S&����i�E�qy�Qʙ��$+Y&������/e���^֌Z�]�MZ����>A�ĕe�3q
�u���!�b4�:�,Bo�Mkٸ\��3�/�
O�@�m���G�Y$���/W�P�Ep� 5H�9��!�>wi�L%�=K=�G?�eɻh�����>��S��	�^t�ſ������`�����VM��N���H6��'3{�)3�c���K���h� ����]����d��������(C2�)��p���r��/��Z����$�/��{0�7spf�h�=���\V.�o�g��3RG�Xh�s�m<�V��C�`P��N[}���!u���O��f1�I�O��L�F���VH�3H�e��6��Ic�����:�Qe���3��H�e�>w�u aI��WR�V�]��u�d�hϕ^�7�w�}&# '��R (���l�eV�@�i�V��%T��T�cIt#�b/>��9��^�S�����k!���u@��L�Vޠ�ң���cM�t��v�Eϯ�4^�F�=������uN@�
k|ːiȴ@o���3�Gc!�^�Z혨> ���k��� �����##�^�mB%Q㬔J�ױ�[� ��Ƥ�m�>����@ ��>zt�x$P�8����Y�>���8$|:C�7�o���r��3�~q���6�b���
�Ч�;x�QVM�锴t׮�ڬf��W-��g�'�8���-��>z_�,�~yjS)lR!�a)��qڇr�o6��P�u���2ɝ.���B��{��74�O���M39-�<���z\[�-��N�mz��_-9��5F�|���ʈv�U�n�uj�
w����F���"����\U	�fm�z��QntN������h�Y��6���F����t]��R�>Nb���b0��력�s;
��LbT�n� S��+���G(�l���"�%��N^��;0u�f�Q����c$���^�r��Hf��2YI�;����\�o��nn.��Xl&���_83-u�׋����E��ƥkQ2�ݱ�bj-6vb�4AC��^�������܀9�����d�ck�R$S)z����;V�z��ȳv��d�dos�SuU3�#�=�jT��U64׈�C�W��m#ݭ�鋯�a r���nר���T6\Z<���
0�# ���m�ȿ�55GL��8����.��
qTcW�5���l��$"���g~<Ϸ6N<�L��^���c��9L5���x�<�2+��N��+q�]r	�y�mJ�# �i�e$�Z<t�l��Fǐv.ُ�һi�;�wzU�Q�Ig8<��K�{� >�C=9:��mM�_��!� ^�!���Sg�У�g&�I�-��F�������T�ɛ]���pkoI'���TOs=@��>*�
�OJ��Ĺ���q��e LZ�TuDʻ���$��P�R���
��7�P����_S���%��lϻ=��`��\W%q�p�j�'sߐ�K8D���8�h@�q�����&S�">�J9�|ƞ�m̰Z"��d��:	����9�Dk�?Tр��Sr�9��6���˝�t�3�Χ�GB6_KX�TP�����'�Qg�"#.�1������U���c�	@7֬¼��z����bh�am��Ҝ��.����>R#�̻8$������b�tk��IV�T��
�ր#;ù��)ϛ��|�j�~-Uh`�K�#]F��89.��X*������\s���qb��;���M�)ݗz����D@M���=�fA� ����]'fla��i� ��8�:�K[/]`�Z�����4�f�Ǝz�@����2��!)&T���y�8%��������?�Y�%�jD�yU�$<1��
��1���9tʉtsl�LlVoҧ����]�܇�/��12��cs�;tF�N���b)�}��h?��4#�uZ@���C�ڎ�5�S��1����=.��b�H�6���h����ԋ�$f9��I��ءo�X�2��@�"��	�?�f�qo��#��l�Z�.U|h9*���1�VF�&�az�'�66�t�6�4��Rwkur?�Sx�|�=�ڶc�o��Ɩ@�/w���u"2����pv��>V�L��͊_�5�
�HhC��Y���L������u%x#����,���K�tm+���l�^�O�31+}&���Ny+E}t�����#��w�}8�
u�M���"�c�B�j��]����/:Ql[r��u�})��^���Ex&����.] G:�ؑ�QF��%���� ������8��)��� ��&O]n�@����O��w_�y�,� 5c�+��N�q#�f��U��ͷKQUGJ��*n�K�=Ee��_I�Q7t]�3�y?o���u  �j-�#�a��ox�U�>;�rl`�dj�и�|R�'�u*��Ft�[vM��N����$x�=�!��b��w�1a��5�Xx�����脠�m����vz{�0;�3	�qK���92���a8����!{���������'Al�9o���L�m`�.�	��0�^����jy_#C5����H�0A澘��`�vwA�����v��r2k������p,�
�%?vq�o��SӦYs�ȧ.O���K�m6�N�E�1$�mll�ڭl�~��zC�߉(��_e���O�)�D�k�#J ;`>=0�"0�����=�^�.�-�y�Z�V	�k�mz|F/�I��a:�^��ۨ��՜�|�W+�,�~R�l��p��#�Br�)�k��;k�.����B�2g��Y
�+]�zN���2��_���=Q�/T�j8�CJ2 7���|�M5'�[����	���[J��f�y��H)I��D6(d���[�e������Cگr�T���o����Ѭ�X^�} `�J�`fIs�:|���5d�R���G#}�����'+�'*����'D �~�Q;�P�tο�F��i� ��B�Va�+q�8�k�I��U+`�e���\�=��̐4�(���阙�~&�p��QQ/ҷ��5z�����-�@\L[҅ !��� ]���AVv�c	�j�*��F℡-FGE^	���u�$~k�7V���=��x*}1�Ecuɥ(S��ሲ�9�4�J>�Y�m�m75�eU�.�3j�?�Z%���j��*bO�o<ؖ/��-�	|O|�6�d�N�����Hl�z�h�kzDzQ�� R.̡�W̸)���N�a2��z��D{]f����C�~���C��/P2�a:J���?px�����:�HXֺ6Z��"eP�FF�^.7�yx�����j��M&��gK��"p�4=B��|hdU�ŕ�Mm����"\��$��7I@N�)�'G_���Rj���1�zb�*��I���im��p�,���V<$�-8��p{z+��\x��o�ͳf'yH$�@0J�.���(�}��P�O�i�n�3oH��/}	^�BT�2�_�u0������ǧ��`YàoW�3�ހ��uyW,�j�w�a�
18��*R"T�y!䨯��Nݳj��0K�}��,!|,����w�I����-F"���3M�U-+��n��θ��ٳ�(��9f�ɠ�B0�����=%(�q���ah,S��J*�cH��2Ȥ��`������	A��.>H���)�ux�(������x_|��!��Dr��ƻ���L��c���1������{hOJ|��g���������ݹ�*��j2�Dj�i^JG� ��De6�� `�����c��o���)���!C�u�f^(�������k@��iy�0��Y�>��=o$k��m\_�+4;����&C��}��ֱLsl����jᙛv!m]����$f���$P�ͷg��ݑ�}w>���d_
�V)W�.����Z,D���kk��U�qg8�+y��.<�3D���8����"��y�ག�~�����n:���.hm'��~�Z�'t���
�+��,'r�
�0M���A�iòǜ향
��h�ɷ����+��$j�N�u�yN�KՠQ�u���YyǬ���	�P��`���O(�ф�a�p{]�=g��O�����f֗ш�J����U�L�(T���\H���,�m ;����h�`����5����`����|o,��
��Z�0��/k���l� }Z1G~z� ����J�R���@�����U�\E	�D���A���w#����X����T|���߱��"�b+U��^rf �C��܃���"S�}�Dnֹ��'�4���^�˦�����P��93�V�����]H!>=tKHT>�����fo����S��X��Uݏ0��g�h�MUɌ�Ҕ_���qG�2)U��|��̥�-Zs*L\K�`\	�Ӧ	�j�S���>`�W1���n꽃�(��i�"K!T�28ڒ
v>pGOL�F���1
#���\(r�p.������=�����R4*Jh�)m�e{��v{���n���Q�i�\oV �_��E1�+���G�_E#�Ë�s�t��}�T $1�/+���#f�t��t��4D0% �(Q�aˎ�BNR��ӂ�YUN��H���������"����m�@[�s�t���m�/ g���n�c_�B{Ƥ)C��FE`-oJԽ*3���>���[��0oM�$�d�NH�#�>L�XG��>F"�@�G��|%9̛s-�	����м���/Ř���f��f���$�LGuL??��v��)���6cM�/fڋFrȆ7Q�ֱ_B��.�p�!��I�ͬ���ZO �n7(B�n�u�S��7��^\�52zu�2�Պ߷<Y�� ��["ܳ���KA�b��b�;�CSC�|�,E�%�)�8��Y���3Z錣ɗuL�� v�^�F�M�u.���s. `Z>�,�]av(��2&�� N�����`�4t�^����������of:�O�+�L:�K�8���@&,���c��#��0��9E);\���@|��1	r�X
�퟿O�=V�C(k�Vl}R��˄S~��]_�(��F�y�H��:\�C��:��MRZ
���B���9��9�Γ1���,~h]f͔~!<�9�B���-.a��g��XK�3)g:��B(������y��bZ�I�7�}x���#A�}���w��o��{qG�� ��5�����B���˳�C�N�0��g�N�}�xD4^���&���6���2,�2kDv��Z�`�~����́�E��B%��{~�,Y/K��Q[/���l�J�,dS&��&E�b��G�ߕ�����>������Q�b����1��ƄL�[��l<U�Z�5ISTu�̙v����(Z�6���&9F>�K)�%���2�jg"��n��K&�#��b��I�
?�VLz6	��N�W S�O��{2�ݔ�4�����>[@� *�*⊬W��%l�֛���.�@���\��-z"(g%�	��Y�����=�;���(���ƣ�����_�xZV��S�&,K��>>����%��pƇH��!�h#8>�=`�R]v�:g��p�3`��G4F���7z��Ur�C����s�/���ԏ^//Ǻ=���1$���j���h��?������l�����}  ���Ԯ@}�ggIa�)R�#����9���G$�>'`��DGv��{ee�u5�9I�_���X��/�9���c���E�~�imˍ�{�h�M�G� 9�+�e�$Ѡ'�JH`ѐF��2$ސ��@/Rg��4�t�u�n�������5A*�KcB����mO��6&BB�k�[�ð�4:���+QXTi�-xI½|��ީe3�e#�J���Mר��V�%!yA�����_�5%�3	(�m��Y零�~I"�,����2Fs��ˊ�n� &��� �Z�A+�=����V�m�nI�+���|���;��E"�j��Q��h���9Gx;��V
.Q��O���<�d�96\�W	����~&�G����N{(�������0 ���[z^�4Ss�%�)�I\�G^�2I���������Ią+ɳx����O}-�3S-V��{&��8����4�c�h�sZ9-I0��A��^#�A!�)��,-�e������i��G��/�ei�6��9�R{�� ���A���8��.g��9�I趭�c��^hwjvH ���Q{9�kr��f��;QptU'�»l�RC�*�BZ��Ɋ��q&��&��RJ�[��$���Z�k]-AQL�S�!��b��-F>�u��!�9V{�p5�J�:R��d/����xYD�J͕O���)�0o�綬��w t�J�b
��]n�%k	�]	$�	�W4ٝ�0�A��U9��@Tb��\�2`W�C�@i����m��C�j{;q p�u
@�I���(�G�bwI�c���k��٫�'*o��ߚ��A�p㾒$�7i��<̓]f&�X�2����f���-S����|��˨���xs���������d�R���'���L�,R�֯�pE�%(|��*�ۘI�z���S���wi�>�h!��d�5���*��_t}Z��T���D�Uc���h�o4��!|���������!}���PV��y�Y�}��=�/<���<<�Q�3����l��8|�U����P�Bx��$��;n"o\�!
m�J �`u�
�]b��Ӯ0V����Z���t�p�k��>�w���f�e�����8a�	J���ǝ�T��c���K��6K��:��Bx��H�(���Gt���z9p�D���E��fX�gqN�<0���������=���6)1�֍�w�`8"��y��#3�]M�@oW���P#2G@���U�5Bb=�{����"d�����MeUp4z��'�aç�$��5�=$+�ȱ�	�ߑ��
 ˏ�t�i��|�1EO���[����GL�/PԻ�Y�����לƐ�ms�`�4��[e+`]Ѣ��چl�*��u�q��ɉ��o'��ɴˌ�{�%W7<��Dq�C���8EA���\�y���m2��B(U�`��H>�98�$d�� �L��O|ɷ4��A��ѻ6?[��V!��Dз�5�N��ަ��!9�+'��F��|f�!�43��iH$�5IE�tpI(�Q>Q!�ҽ_��G�9HV��W��_Ѓ�Z�h�9iK����6po=v��,978G{&���u��0�?2�o��c�i�5�~6}�G��(b�h�W+�<��%s��O��W�	k��6��%5���~�~�PkT���8�[�!8Π?X ��"t����AF��Q�Mņh~�s5Q����X�6 �M��5�?&K/����m�[%m��������\ƴ]	O���[�?�K���Q������R��{�����ʔ��
�\�����e&�;fBY�tg��D�Ӗ��(��0�,ʲ2�kY������h���%8��}d�	��g�UI�Y��W,g����ϯ�Q_l�@
���������g|W�Y��S~ӛ����# ������v����!��4j�����t�2B�nE#�EҚ�U |?^�*��{���q:�W�&)Ū�@���V@2>qF>�v������AX2*�
@t��o�I�й��`��+鋮���>{�("��Apgp��B qp�n�^�N$O�k��e���6�N�3Z�le�Vb���	��G��]�#�+I�n���U)
b��n7��~��<�8�l�˵�*���C=�;I�]�މgD�.�g���,\p�79�=벯�M,x�������!J�or){T�><��.�7u�Q�8��z� e�\v��膰�����jۄ/�帒��5���<����ɜ���O:���f	LJ22\)>>�?�k.sRݖ��H����{��)�H�<�i�K{q�W�������T�������3��\�<U�a���r�`�ێ ���@Ц �CIXu�L�}�H�q��K�
�_GAj�{O� m �j�q��4�z�W�;Ȉ4�� �m9)�}�F���Ω���Ε���Z�� [����mD]^����*u��%
���J���%��dг���ջ$��!m�~ThqE*�lՇ�gH��1�]�҆6������#���`x-֝�'�}��w���Lic�6OCv"�Y�>c.J��ܪ� ��|���ϼCԮ=��o��	����$�m����_��Q�:������ɵ��|���>feK��o�FX��h؃�6E��q�lt���������++�U���� �	�H��ӛ^���8p3:gZ���}�,N���k([���G!
h;=(9�1܂�h^�0��k�h1�xV�=�6���(O��-��[	�h9c4}��g�Q�;������!���:\�&�*�����~�Tzu����{���|.h�6+�y�;��ظ�S���)��~KB+s��8�E;RWǇ������~g�n�)YqC��~DV"������J.����HU�`�T*�a�J		+Z��E@���f��+5��(ti!���$���檬��oy� >�g�I�j��)v��;�x�Ĺ/mc�6�tW�\�=ue
���q������{`�wט�*�!���'Ik:T��#T���k��k��r�B����Y���$�]O3ҡ$�]�s��6_$����y��8�5Ⲩ�^q�lh~Գ�qLZ�<���O�&������gmB�d�0Q8G�z']�p��&W�%|�DJR*g�ܙ�6s3I
�S*#I�P�Km�����`�]*��`�����˛��G��XNa���ó�]%9%���e�6�U����
�����1�ⲫZ0�C�+@.��( U�؊�1�������g8�V}����M����6�(P���5�2�7��#YfEɣ;��7;�@�<�?�J3���&��?�|`��e�e�H|�Q�DK��x�z��F���΂3�� (���*JE�v��&[*Z�����c�z�C��wS���|L�/KP��WE|/������3��p��V�r�Î�i��� S��}0��bY������՟F'�ש6�:/��a V��a*4��87�5���q�i���v�~ಁ�~�(̄[������W:	Us*��P�:`��Vdc��3e�0Oh��/��S�I>[�O��n\���蘊!goV�C���e0��[D:Rz�_�~4��I�8�d�n�RN��M�H��Jx��������٢Z��
�=
�cKz��2�c�]���h�.��e����gcD���,8`?_�p+���m)P�Ŗ#p�gxG�G����q�77 �]0���`��X�!�Ul�^fC�� !��§y~���-;��\C�a��c���պ(�Yw�ɝ�!�����wQ,?��wk����/��X��;R<��g��~_k6]h{�����~�5"���w`h;���	�x���+?�_�U2M�f��R� 
S���my�wr.h_� C,�vD��	J��T=5�8���?��F�N���Ag�$��8��A�/��a�e�M?��$P��!�Ͳ٧��N<�x�3ԇ�Fk �R�N/y.��_��KqF$+�O�����@�!�d�7�� w�(Zl���ÀTL� !��.��i|��dۛ��-{�� ����.3~yUxV&��&���e����d��G�<���)�.��;fƂwK ���&'��$�?�JDM.�=���/!OW�s�+�-IBb � r5vS4��6�9��hǃ�ۉ9�W�ԩ�F�s���T�Q�t�׃@�^ h�z���SMy��KI$�O"D*��9?�ڪ�q�%zN��O�tA�Td.s�.����
jq�K����>ӓ��4�8�����K3�:*Ҷ����ޙ�G�ov�I��q�ۈl<RC�V����5
���6Ou�]h�՞T���)F��M�� �����MWB�b����i-8�q�n�l��Հ���sV&� O��<`��;�{$ߚ���$�a�\[�q6T.������ɍ�.Q�%W��:��NX���ŷ}c� ��)Z���¬��Mu#�tnR؎�Q4<�"�V0�}�Q�b+Q����L�G��TD�^a��EQ��a�Tm�خ����e����$Z('ޏg{��*�b�FU�'-�%s�{�
��[��Tts����H�#)#��"' ax�7ŵo7Xhͽ��̤���s����/8�/���N�*��o@�S����R4�J��-�������k��/Th8r<漒�|�7P[wz� ��$�v�S��OQ�%٣-�M-л������4�����f͎{�)+r[�~����ͦP*\,S����m�LE�����o�L��2�鷺��A�R��i=�o��E����`CT2�h����s��~��ً��w[x�ʫ�,�C�h��̭_(��[E������3�r6�)���m�K?)�3%���ȏ�m��D��h,/�v�ݡ���F24U�"�T�?�X<UK@W,���W3��JM�v���nbz����	�_Ln�������G���<ؽ��+�r������:h����ӳ����o��*㼮գ�ׁY��M�b+3(��H�X��)3ٓs�QA<<'��F�M9A�,kxi�K�E�.ȕR�2t#��%ꅓ�3wQ�#!���^6������j�7��u~Hs#"`_q%~
w�F����@�)�mRS/�f�{i�o�	.ë�w�th_�~&��w�m�N��Ff�߳�Vo�����*q���[�p�53�>nˋw���&�ĵ�^ߙ-*��:���ꎁ���s�y/���}��oɳ�ֹ|��3
��}�� ^
0��1��J�f�H����F���s��b��4�vQ�V��m����`�c���P
���z���	pw�&t�*E)�߶�tE�K�:+MJ�<�Y�B��ᘉѬlJ.�#���ʅb���n�'�� ����0�`��k�N�?��qa�j�em��nd1����U�$g�V�1�s����!�K�t�(�ߏ�(�_�h�]�!���wU��g���)��(<֏�G�W:\��x�2��R�����)wp%��>�d�9~��[��@��5����ط�*�r�f���0ތÁ>ߙ]��Р��6Z>����#_u�/�l�.�ҸƘ0!�ɭn7<���" x�xN���Q���_�p�9�گ�"��j���)K����e_:^�GC�x��`�j��~��
����!�o:Iu�C���Ϫ��?m���=�� @�u�r���+�5�����w�����f<dC�LD�{)2���@��Ws0p15�,�,���UW�4
ڥ&Ӑ�T�ؑ<�ǰ��j�k�{c�P3HyWQ=��b�H��v�����z�f	��A�(��zo%H`�er�ꖳ]e�GO�I��g�w%�yv���Φ("cfv���k�kj`H.
'}I�#����)n��D�YY���N�v7�NR�r+�f���KAt���i�Ng�2�E��U,T6_q^��R��1���OZ��Zsm\I2�=q�a�X��|���r����P˭i�H���rhՑf��8�����
.�$� �M�i�6��Q+i�5 �}�2��%UϊyJ����D������!`[4�0~SO*-C,a5\�._R�<^�|�8�P�B�
G�f�J����
"1��6��[�1��h�����+s`i@��L���N���Vq�{�Nf�"��Z@.P,;�9�B�ʠш �	���;1�S�ZG�i��9�0wd#�ͳ}�1dߍ��A�p_�!ϗ�OH�5f�8��z��ng�ڴ.�������4#:G�I���+��zo�|y�f2] ���&���Ș(�P��=�����-bC�^p&��>F��!'�����>�%��GTڔXۼ�ՂX��B��y�Ġ�L&˴����'��W*�w��؆�5k�wN���]���]4��6�˴O:�̱� |�CZoG��ҁ�H�Ec2U��	n��i\�>�u~�Uq=�QZ(2j=$��D�c���Ĉ��M�X�[�O;0S�Ԉ����������s١��fv�]d�t,l���tm�Ɂ�G9	�Z�:~:�rRi:K{���}%{d��!��5�����ޕf�(n"��0r���1���n�?z�Y��S����3�ˉ�f{gW�>cЃ�"wH?��Zݕ��p�I����G��Ү�Z-��0	�'��E����~����C3���_e��u��g��3x�rˆ���/�aJ0+&=`�E�d��Ƹl-�����TS�a��3�W���^u\h�|�^�%<�݄�]�1�2M�3���L��t�)#��؍¸��[���=�.�x��HZ���zЮ0q�^���ݳ���%.xH�VO��ٛ�&���lɰ��qZ9�[M9Ci7э��U��0<T�db(h�PT�v=j��C�5�	&n;U��S�Ɛ�YCOo�4&����ђU|Z��|�����Qm�ވZ�,=7bx���Y��U�MR�����z/��oKZ���UT�оZ�1مP<��H��H�;���f��Ы�٦?���3yf�C"wt��TQ��
ۈA]�.Z�����t��R
K졸l^l�4�z�G*=���H�6.�u�eǊ��+��2X�e����3W��uZ�MC0���Øֲ�t��=9�C�3�k�"a<��-�L*��/n��"��_�kn9ݘ�ol;� ���A>�B5��vk���K\�i[JjЍ!Q��3���L�x�z����2q�T����5׹>�:�Ӝ��N����-��A��O�֬c� .���z)t_�]�����N�zf}0hϋr���I����8��l��$��q� �hf1!_�y����$�͇C��fV�E�[؀������t@�c@�f�2�mPd�.��KgzŮ�_���+JKU�%�1�`g���Y`8�ڎ�1��_�l5킮��M�",����d�v��(:̓b�e�F����q��n��Aa��)9���k�|�����}��F��R��X�a�s� �#�3�� >-I�
���i�
��������^bM%gO; �mEXF�H�,��2�� ^�T6����L�j>S��.���K]}�9�ώD��g)��5p[+v���491���WcK���?هs��7B[�8��_�ʵg����?�5�/����M�ϑczƖ��wס��;�e��+x��N	[���|�J'BD,����p����#�.���5��t8�GWm#Xd��D������on ����p�G���$L���jk��|J6�v^���Ѫ�`� a�I(�t�eK�7�`ک��ŴA�V� ���]Pz:Z�/�Vu�$O�����EW+}
o�#׼���I�޵��7���IxW"$���i�<F���9D��U�?݀vHSk�m�ڣ\��L�G�z��#Wb��X-����&E��;ەͧY>C������A�3�����Z�%��� �4�T����Elr������E��ׇ�;�����Ѣ���	��ߕ����C��	y޴�co`��[�΂�0�X�p���9 M<*Kޯ�)I�RQ0�}�k��.v;@��T�G��"w�@|�b�R'd�N�uG���`�.��l����1�������ڐ�W)nT�pѴ�����[�ԅ�3�71HJ�-�IL��o��.��7�Mv߃̐��Y-��K�>T�� ���s`Lpm�X����/'�M�G�EC��!B�a셉"� ��u	v�M�)�T����gV�/x�֓+*�^���.��d�K�-����2������$��g�u�?ڈx5��,��y�}�5�,bM��i.b�.&D 3ז�{��{N�L���y�'�3n/
�d�Y�)�@���a4Gy+J�˜=��_(��t��C@Hv�Փ��5��&�����O���u`\��Y7-��1����V�ɦO�ë�����!Pa�<K4`�As1�my]Zw�s|�t��,�����'�Se61�N�M*_$�HI��0��bz.�z�цq�z&�9Q�9[���$�*��h��1��?�� 	�6��gU��rE��K��F(>ii�y��^뺫I�Y��[^\�Pkt���:�K|��2�|R����R�YNѪ�&���d=�bb��}ѫ?���}�O�h��Ю ��%�&�&�t�4/�����B
�zt�hBh��������6��=?}�h�'��o��YoLѴl�;��6�e�X� �F���&��z3��w-0�P�&,�����aD�,��ϵ���(�L�tQQ���P.?�=�~]�:�ecؼ�!u82����pR��*�1b�D�}�m'9�����ȫ�e�]���Ԥ�|g,~R����Us��P�4U���B��i�+˚^�,ȶ��~%���)�)�ʉ��v�d�3 ��@Ň�'y��m
������yx)1߫���c����#��ǔ:5S�d[�hX@05�}?�������9��p�",a��g�x\�&?�._�᭜� R-��ݜ�����.'1; i8�p����ӁB�,"^��lL�w�e�3w�����#�D�ӧMN�_oSn�b����+g���*��:��i	��)ES�~}Ҳ��e��vw�x��O&��=jߊ����_��������>e�"̨c⽲ȟ��W��[j	��{��|��B�N?�P�j;V��eߒ��޵�[����/����Ъ>��-��%��j��g���RO�C[�8���d�b̯�L�S�����=�PM-n���C)�5�A����~Cm^(��֫��ׁ��j���F�&���8i�I*eO-��L�V��T1=<��2�49�Si����h�5�K�L�K��|⍄������x|)G^Nx�Ho�&p�1�e��rK���.G��"�v+7m.1�Y?LwI�����T���U�d���Z�P;����#�C)��y.|�D2�KQ��_����ۜa���8���3H����#�ء�NB�����A�1u����{�0���P�P��z|��䫄�埏��[W��9�U��)�3�.�ٙ��@"k)Ǧ�E>����}��L�څbr���w� 
L��zʨŌC��������r�8$t�I��9h��n|_��$�Gğ��ч�i4Ly�R-gUD��)4�19����4��rҬ����4}�]W�"�#T�/9qJ��#{��f.�{��[m��㒃U#��||հ�$�^�=�f�Dy�_va&|5����_�<Xd��	zP
`�{��B�b�a�Xî��2>}1�@Od1@GIs�u
2�S�Ų������afW]A��h�ĵ��ى��~*��a8[*�x�]q�t1n
����g��Gh�*TE��֫v}"-t)l��ޮ��[ՋG4�0Ko�o�頩�u]�Ϣ"U����T�h�T�9�J�5l���K�ʆ��%�IL?�g�=��q� ��t�~Ǵ��=� ��Y��*i��G+�;��{��5�����y�����}�����j����z����\����u��T$��vɥBz�Ex�:��4��uT���m�87�ˈ�dT���V�"e$J9R��D|��vUN���C�����.
�zy�d�$��[�l��@C���]a3�D���DL2S-���|_ʡ�I��^�?��\��]��&-#�Ew�]��(!*��ڂ�̭��Hr=�u�2����	����Ln��u��|NM����N�O�J��:5�[5�LrˆE�Qg�9��`�-�C��6�«�ɗ���Z��$o#��"��S.X8��@�k0�Ñ�[�LJ#��W����_�1���̬��"�� qY�6H����5�&�[��2�!�� ��ۆC� 5Vmq)�ʇ/���C�mPQ��9����On�8:�%|��7��K:���ſ�s����"t2�#��II-~JWmD7Vv�ba=�j�Bb���a�=.�z/�ik�W����r`�s,Zq�����V�ȪFj(j����B��k�3;�}( ��0�LnU�� �:ʗ�b��Z���8�P�GeL� ��N>'�ؘ� ���>&$J��7��m���nH�3|;G��.��V���P*��%��Y�h�u�*�| ՎjN
J�8Qs:]���ݧ�g��������g�4̄��Ug��p� Iκ�9��!oK����?���|�:�4w(�r�J�-!�F�]aJm�|Պ�%~�GY��Z��w?%G��L�Mx�00�tjH��~v��6���s�2|C$`�!�n�Nk����/#N�^W�z�1���S�KS``E����B�Y�D.#}�]�W�Z��������VL�#o�M���j�F���ɐ)�E�0�<�,��-�/�%v{�@C_�A�%Ѵ�=/�7�^��=�N���㵵$��.��y�	����A&�O���b��}̓:�:/*�{)|�$J=m8�!�@,2@B!��:���+v�{�n�ѥ��1\\Ž�O6�Q��m�-Q�Kw��1����:��6��</V�7�Jy������b�ҙ�X�P���-��<�r���dM���1')#�I�O��ɨ�N�����n��.Ϣ�Hv��n��ؾ%^�3^���(ѳ�?U/ۮ๽��=\8�@�&�KP�xA���dAQ�s��@����c�V�j ��W�;�#w2�P)�5gv�7���#���W&]k��TWlv��i>��xSfJs�f��=q�k3UC�o1H�Win���B�f��WE�L�S0ق�¨R�8H��J[O�Z��Cw��#��$�w��9��2�s���~*|����o=Q��"��Kwj����~��l&�^�}�N�&����R�LR=����h*��0�-��e
r|{��'�� ��t�,�t�R����rċ�1l�ǅ2BE��Cؘ�����m�CƃI��Nq�j:�N;��"�=����@��Q�]�'e���]��F϶}�bL�^��1S � �=o�9P��[���|�'D���ޠ���S���%�cC�9��X�s��zhj¬�@��Jg��S�3	�@m)T2��}!h���Ԙz`83���e.�,�;[�mD��2$)�|u�'��bTB�䊄xmD�^s�cf�!
V��_��@�q�!	8�Ε��ZcǛ7bZI��t3�]���B<tx0Sݸ�!�
f(��7����l�2�L��K�3�N�O�v�'����V �`d�tB���S8�U��Ou�-��=/U5t��s���<�/AT*�'Zfl��K'	bdI�G�ԣZxֶA|BI�>M��������$M��<'^,q��E�u�1�)�޾�֭�
kھv����jQ��w�8ꢚ���Vp�����,�����Y
�Z��L�2��ʳ�z��w��BC�b�~&]N~�"��G��ufk�	�MH		��4So8�1]�s<�/ظ�8�Z�	,TӪ��{���s>�:[3�0ט�(���G��/�I�2872ԚbD��
�.X��b���T�u�iY�P���W���j0�s�%�gI����Pc�쿴������Pǲ>S�����6�flɲ���O�V��,�����>2D�Q�@�*nR$�����_����^󛷆e+�b3�f��/Fq��b4��s�H�\�no��l�1��f�rov+Syp����ӭ�81�rK
���څsƺQ�D|Fq�Ȫ��&���К����tѰ~���>	��`+ۗURͷ T��u�{;uҞ�a�>�T�3璇˹��Z˨p˞��	�@����%� ]Q%��o+rWG��f�g�㬧&̼d�<LA�|P�q7�9㖕q	�V��4v�-ƬU\O�FJ��jcX����v5���W(@�Q�'�'��st7�9NOF��:�p����v��@m�~Q9[�`���f��G��/��m/��<�e �x����N��p7U-T<�&�ǂ6fǿ.�����t���2��;뚞L��n8�"1��=e���ܲz��5���ڐj8gV����篎s i�Y�I���g(�.L��� �B?h�Vo�ɴ�W^9$N��f/��@L�k�o�*�ZKLw����8`�����u���!����Q�G4fU��V,���u�FO�'�J�j��EY/��hι�w�zS��C�O��X�<f8"Hş�P��M�lε+����f�AYN5X}?�������"Y�Gj�f�
���W�ц&8$n
~/������εL��/�Y(�	=iA�� �E�����z_8}!��j���3듫�.�&	�A�{�~�3�
{ 8C&�>T&�+�R&d'#�����8�(�%����}���w�*RH��r�[���ܴ慣�.��?�R���4����!��륥�XH�����U͜IhV��"sGst��.%��{�ac��mu��A�0QR�������>�?K�&��2߶9'�Ǿ�O�Ƴ�P�-{XHN�I�����ml�t< �B���hz���(��zx�D�%�~fOb��g6�N�C�T� $?.[��q�XW�X����u�<�i�,�&����nB<=��/�p��H���gP����.��B�
Ha���|W�gD �``���k�o��RŞ�s��E��+���֜�ߞ��7�
���������~N	u]'�`t)�#ec�Q�xX/}wY`�v�F�S��o$�dQ��,"��Ղ�����XJtrNIy����즹�/^��V^�����;���a��;�'6�X�n��:�:�H�f8?9���tr/�����wM��vb2迪��v@1m��0'�M�bC�e�ڑ��m�)�DOG�6�t�O((�h��w3��]�I2��H+�7��I��*�e��-�&� �+���z�z��
��T��D�1fB���?ϒ�㲚|p]������d1�'���3�h}[b��7��BV�o��6F�$NH�z�X��*���x�����I{������~�͖��	pM~c�7�n��ZN��}F��w�F�}���
�2��i	��XE$�h�~����^uN���[|\(��E��Ra�.��T�p7r���*�o�_�GL�����w��~`y��mO�a���O�n����$|�N����>�#�	-_�4�Q(�hC9����c�=4Z��O�ZE~� �J����SD��Ʋ����bo���)L���g��p�!�=� ���H���p�BlF�L�.![�����
�-}��߳���7TD��j
y\L(��hM�<�sN�䟔\�w�_�� �m��)?��8<p�	�r��a��c{�n�L@!�����Jl�ey���.Ⱥ_<#�!O�-B�?@D8"�\&©��Yģ���Yl �����n��@����'?�m���{���<%���LG7�4,��6�rPK����&)��������_U�3��u�R.Â��z��'��vл�/�WP��׶���>���_�H�1o��j;����D��<�kyp��+����}�S&h�˓���c[�M7�;c�S��49�Φ[�v*b�w�r�Duɲ��N�\(e�/����DI��I:�x�R"v�`������D)�%P��d|���&0���f��-�>O�+K��}��.�^�������N�?W�뻐�6�m3�\��C*�.��*��ߪ�/�`�JQP�h}����V ����F1����{PAXR��@����X�Q��IT�O����)`��zN����XVQ�;���45��Q�s֩ i�/
���~��A&��W���	Ȋ���?_=8#�#�K�F���J����%�V [��U|w��J�g��{�[�rÐ���V��F؁1N� N_�!_c�%<�����G��R/UE)�{�)�`ŭ�.�aL#K�^0�y�3 a�^Ǭ:�?\���G!68��H����Lz}������@�ݡ���
�#M��eJ��\jJ��/*�B���<�����u��GqzI�20�N�5�C��$߉��z+g�dLM�֩*���lS��j���W��'V��o��Ol#�e{!iԆl�W�Bk�d?w�d#�8]�̹:ѰJ˂"[�t6���J3Q<�N�ꕢE8»�T�/	"��WS6�k��;\*,y��X� ���u���"��|SI��!ܢ˦BP���}J�h�~T�U믟�Xj�R-��<8|����Ox/l�9���{�"c���$�j�rNn*�5��c�,�0��9�O�i1�-���v���<_N5��Z�\��s#:�f��e�ځ�N��_EI_ �����	p���N�_Ε���1=��`�������E\i�����9�Oƨa�9G��j����{b��|�$dAZ�A`]PA�j�0f0��р�ei@F�sw�HIR����X�%I�4I��H���W�ӹ�z�='Zɶ �f����pp���(���C+  �r>�jl <�)��[������F�.82�\��}j�Y��uڐ�3$�K*魆j��[�v�$�$�f���B�u� s�w�����ƩKo����Ї��]����dc#��K2� ��Nϳ���ƍ���$�qʫ�Q��
��3vC}$o�K{ʂs��/�a�x#����Wx+��ӄun�H;ɓ���V�+���ޅRt���,����\E.�h��KZ�����PJ�r���;t1_ꬎ���ا|���e�+;��~�4WJg>΍hGy��E��^_ہ��wH��wr9Q�ڿ	z$W{�]���I|�)��;�"����y�� �$F4P��6�^ �L�(kZ����������ܸn�,�sĆ{W;@�޳�9������}5Qr����KI�b��*�O�=����Xw؃�ɿO��8�_���Qx�H���<�����Xa7ѹMj9D=��N·/z7)E`�Wp�ї�^m7V3�ml���[)Hx=��z���;(�]�z0(CV����q�t�Q�[��=��7�~�T�t�qC� �� �{e��(ƚ�1�1��W	�>�7^�М����װ4��"�l��Fi༤�0�G�����6����	���U���iK ���=t_�`������܎n%�;�����_�8˒����,7��H�����{B�s��շ�'(�� ��Su8�5�ș����ez�+��r��|�t��iI&��/zA�e�J��B�k��ܠY�vٵuTv7MZ �+ۆ&��(E �� l���0v�7���݌L5�Re��'�x���p���a��dI�Qȭ����M�U�Ð	&`�w3kA=[�P�NN'B�H��(�~<���]�ce�*ܕ5���0_��(7�ӑg�R�*��B�ĠV���`Y�Rs#=��,����O"�,G�}�[����au���#��O+�v��~�xejk�n�����4����s��o�EǱ���}r��M���²�埶3� ��r�Bp�Tuܒrjv��\���rx��Ǒ�����_~���ID�#��^�Ds� ��H�]�����`c��ݧ{� ��E��ND��',O�2���5���f&�,ρr)��ȭ"�~���m����zr��JV��OȻd��[��Ԡ[F;Bw� ��e�ì�)GJ����.%�u��jf�&T�����D��Q��?���ym��ohۢ�-їu��n8WDLN}��:H�(����孑�4ʗ����-?Y��G���ِ������EN3�^w�Ώ���1jÿ&�I��hQ�n��ˀT�O(v���3!��R-��0����黡��9�%7�^�����Qd���f�hs���Q5���Bi;����}^}�Bd��zy�;�C��b�3��:��.e�w��������~}QB�@�D:�+?��'��uvwe�G��wA�op���)<��<0%3�����ޒ.c!%@�/��X��5v ߳/�Q��Q#d�/{���:�iň9>��_���u'��RH���I�n���D��X�CY�×�sxv���^h����rTIk�oAHG�^�<Y��\^xe�:��`��O��"#Cn�:t,�)��o������Sp ��+�����:�@���/�)s��Ԛ\���p�&��L��B����w+S��� �Rq	W���R� W���j��z����W3ʜ,~.w�=�_>Xh�
m�S7�Wi��a�xʜC�(Ǉ��	{�f)��j�#�|��}�!�q,�9-�- ���5��&�LD��}��bؿ��ۂ���Wû�&u������u���.`��0
�Ȯ�/�����Q����d��/p��j����I�*�ij�g���	���gy�x�
/�>ڛ�k��(3�E�>Ŧ(��+S�"�(##q[
k�� E+�ǵ_��\����^�7v]8�.�ԉ^[�'�8��v�{�>��h���4��i���o��Pj�c�꩹�;c?lE�	k�N6g�U/ ��Sϧ�O��Mu������2q����aT��i:��,�L2C���h?V~P���ӕ�qc䂌���D
Ln��&��EDA[��-U��bW�:��x�<��Ә�B`�\g݋��{���ߦsԔ�e|(��"��7ev�O�q"Y>q��|��a��B��ZD�b��L�Mg���f������������$�mk�{�cevF��Gye��sّ���Vn{Y�ݳ?��6X9L�G�2�߹���uJ�^��)C�@��%[�)�òn���z�*sL@��d����.*:Ǝ�/�-B���'}l����̭�y�_G�"��a,�p��Ńl�@ڊ���*���fK1�Z�bj�[[O��f�B��3/�T��3��A oO&��5��.��_[�(�țq7Є)Xc��C Hx��e<
#�03����Ee%���L��3���#d�],�-}&6�����`�9*8��`Q����f˰!z��1�V�d��|��*"d��I�"0b�N"���xp�O�t�2Vi��n�"��ü��s}T�+�ō�[�e�#$�k�I	���(���_�p�=D���y�9^�d��,���P���\av�`VDkL%>�5��na:)঻�!�����������&mn�8��*}3�*�N�B�4���]a�P!&���ld�F-�Ǡç`��%�B�o�d͛1]���6�������*�r桬d����^�Ѷ���,M���^z'9��
���N��>�WM�5���D�O��z4��%�<C�h�ɷWa�aon�]x'�^E �p�����ᣇM��[�D�� ���<f��q0`�;�\г����%T�"8gMS�Ft8�^ ��+�S����ø5�E�h<U�m�G�xa�0�YUzH�6&��~A�%��v�1nz�t"$��@牛z/E@�܌9��ƅ���}��M��T�߬ʭ�)����2�&q��Nơ�,*�������&� �Y�H�"��ye��.�S�z,�Z��:�4��Np��<�����u�O�(?���h�}s������a�7[=�׏e�2���������u�9�G��6�\��:њ���d_I#���K����<�ƷS<�W�QU�	CtU*�G�hT�l�hD��v�=��6�QnIM�eP��X����@V�2k�q�Lq�o 
���YN(�m���k�"��5`$GU0�MY:-����39яd�U�Sy���+�݄ʀN�b��I���]!�&��uv�A�6�.�(e����a��Z=	���Z�M�����GF���	λ!�)'y�r��
ŏ0kt�5�aF)�_0��(���9۰$�Zmjܱ�u�<�����_�>�ݎ��zA(h���<s�)�60��G}�v<���7��j�:**�,�/�XE1L�������66�*7%���ufB�qn�(�&��ͅz��v�����Ļy�ap�e��m�P8Ӡn�5�4۲G;t������b�������Ρ�1�?�8b�f��5't���AV�ĸ�s��,{ք�f�	�`��ۈ���`�hf�˕hl�81��VԞ�~|֣�����0ؼ9?,��{V@2��[j���C���7��,�χW�����+1W���ī�_���j �䟺�`�9J䷸��։! ��BY�����W�LJ<��Eg��b���:N>�����M0���B;����ܹZ2�B������fk�ϩ�
q�px�I�(x�F�DD�ϼ��H�ֲ�G� ?Y����܊ʲ��3p(�4s%%8\"敱��ri�t���]��x���O�X�'ݦ�1<��e}�&����n��7S��ȼՊ2��D6(��j�m�n��حF!�9�b�Z�ph�(o�,f�6�>��+���ݭ���� �P�� Dk�b$���!�0'�t6o�U�9]eQΟ>�}~N`�K��r�*�x��Ǘ�=����#�|6(�L��[��|	=V�0g"!@\[�_��Z�v����v$yy�����m�}���$�'#��t	m��ɛ]��ؑ���g�*��Tu����P�3Kv��N�R;Y���ψxǹZ�޸!������ �ϽsJ�y�ì�A%�:��j��P1}�H_#2�Eo�?�i�m
#�s�|*� �F� b�(`��j�ncI�AQ����~�(��lKn�g�Zl~BP��բ��AN�,0�u��F�T���M�%�\��JD�A��X���&�P�Q9�O�P�f�*�����"���nD�vMs5�K���S��|�-!�C$x�"�6�?��`?o�~zP�b�*a��2�u�Q�h KFR�]�,4��-�-���l��o\�Fñ e�9	��ƀ�����]Tfm�e C���#�$Sw:,s|B���јW��bE�Q�}��*&�Bo���"X�<-��r��}�q�`�������m�%UDeM���,�r��m����D/�2zF	w����":�m~����[�/s�yA+J";���@��@�(:k�.zl��62 ?u�Ht��^�o��S�����-]�kL���淚�g����+��Zj�D�cD1��K�E��H�ts��b���$,��Ϙ��js�K��R[-���ܱ�FcΠ��Y}�d��C,�a�7s��e�3�Q���D�va,<�%�o)ܽ9DjZ;`Q|�B��Zd��� Ϳ���2�:_��Т���G\��D0��C^@
�����EϹ�|�W[�^�&�0��������ǳ*}�y��$��>�C&�ܙ���BvD���E��ۺ�F��x|�_b7�5 ���--8��Y�a���O��FB���i��֢X��bo�nMvEP���9�g���%W��+��LҘ��/)Y���P���S�$�A�W�s2�}��t`AF�=�o�q)?Ac˒]II�d����М��Z�Nn��_��D����#YciyTA�l�T��bC���N�ֈ��\�Řr1ڑ'i�2o��Z��?#�M��HR�A��j���ŭ��~˶�4P�r�H���$��F��d��v1�9|6���P�	}n��+��n+$��,�a�ey�Yx���8�<Y^E_��&�d	=��ܕ�M�`O�˚HQCM��a����PTb���r��;�`^�pO��_F�%���TT7�}ąy�����Ev@Z�[f22�&��_�s3�L�_6KP �����+\�D�ۊe�7��M�M 'Fv������K<r�,���_m2��qJ�ՍG��.�.J��Dh���=8�t �c��(�n��|�'�%�c�M��Rh5��+4b-�xz=�͉��"s�^w|�����.����dk�\�UB5F��0AYI��`��0V<����Ioz��.jA�d���
2�v��D���C�l���w��Z�����º����Q���9���z��!��\
�}F��N&�pȊi<\Ǜ8�ͥo���#����bLl<�kY�VVzq��Ke���PB�^�k��W輨M[�Sk�;!�qz(I��Ys���u�)�t�M(���+Qwa��i�eߗ�6˰8��$Ғ&gW�/�m~�A6|Wv��M�'|��[Jؗ���
��s�\���!�GS�/�]�e�_�m[�7*�1�
��#E��=���e���!�fm�Ox��(݌�{ ���<��;�7���+�A'�;3��T,�O�|�pn����e'j�Cc��	i��tW����;~���P争���b�%��:¾8(�D^[#����/�=�G�-Zgw��M�5|�#�d*��T���Z#f�9��r�%v���w���\%��4c;�ԡ����M����?�L����~��� �#���	��^#l�ܤ�=��X�J�6����bX�jY��P���D�L��1g�"��k� V�?.��[��Z�QN��0�_!�y��^�F����:���0�:cl]�kjS�5H�#([��S4�,az�Qy�I�8�D ���A�C�e`YKK�!�P��'}� �";�
�S����$S�</��%{Q���������劅�7���0[+��X23�i�Sː�_������R6�0����Ny-�V] ��Z�e���wS �ʬLE��eD��g��d����)��1�u�棈��j�$�Ζ�����Y*j�&��=,w�����\�!n��w�۸U�S\og&���M`�u����G��3"�M�1`�4`DJ��3�;ҫBk��ڐʴ*�3������[/�ZZ-�o�R1B�xl }ma�'��9&�q���Bc('��p-�D�FQ��lQ�IO�g%��{�[F��0�x��4�ym�N�MU�3��:�{�ض�~�D�8�37���@z�_�d/���d��P��~�=��Ck����r��Pl�w�\�.�B��������?�r�84�]М(���Sޟj��(S��I[�oP1�Ԃ�z��X���J�J��U�F�O�.�BH��T�,Ȉ<R��R�1��M�f�{<�3�>��un3��VUM�YO�X?�ձx��T�c���5 ૉ�zm����!�"3G����y
i�fi)3�AF
c�sg����J����u�k!Y<����Eq�1`i�ؔ�$����i�eLR�-%I�kvm��v@��YFL\�M�5:��8q-��MK+���+K�|B�Y���_E��B)��:�B{�uo�Y�9��w
�{+}�������/[��H��o]�R�#�:>�l�ޛ�����^E��LⴎG�q�Q�g�,�x �G��ӴU6��z��A=���g`�B�]���(3d���� ^^GW�r��vqJ��Rh����7H��,����*�w�t�[2!g���UZg��l�,���	g�9��=��>0zY��8!�:ucS,�^vt�{�?H���}���}Xts����݀t���1Y���D3�s�/����~�vt��Z������`�_1�-�O��o�^2�7o�7/��j:6m�bڈT�E����H`�a+�q����O��Y�N�Q��-�l��r]I�I�Ơ^�JN�1��3�q	�f5���$�[�ę���	���:�"|���@g<"3����"T,:'�:܀�^�C6��J�.}�����#�%�(ӑK!��W�f����t ܸ�ѷ㴧����h�^�L���.e���u��:@E��Y���9������-�`������T9�� �9kY5=�Y��g�](�]1yYry��9���������_����J��:�10]���Ye�Ԋ�י��X��1֬���6��CҒT@/#x���gcD��V$�[��*���$h��}�WI&��N\ĸ7Jo�YVXz����%e��[�������{#�3ܦ��%=R�jj�<��U��B�#fnL,��**U`w�2�'��@C͑=W[�+=3N,o�=�%We&�%8�Z`�OSz:��d�v�1�Oѕ�P°M��'��@���,UU̖.瀖v�8��Qδ6ޥ}�����*,+��{�ҒI&pGN��A�Ŀ����[�P�}�k��˰kw�%oVϟVg�$ ����9�`����\��F2#�^q��D�T8�U&��5$i;��v ��0�6O�O��M��m���(y����,D���T�f<7�5�����#P*~���$���2�ϩr���M���������@�� _DcM����-�=��۾#�������W돪��u��7#9�e
��������m��B�� q�P!5�����-{�� �����yY}t_��V0��(�7�f42���,p;����g!kxC^�8&�H�0Wn�
����
:֐`�I�g|d6c����ew-M��t��b�y��m���=U�47*@��/D��ԯ!��ٰ���M��)�:���Y�th2��:��y�C��T<� ���U�.6�����v�F.<�[��X��9
L4��Z�`.�Lq�{���������>�uw�*��00���	������-m(]v_��+̥Ґ^�P�/>��k���W#��zJ9�,�xSb��tZȽ1�q�X����/�`�x15��h"�W��8�2;r�.g��#<�'�7�=��]>�@�'�<c{hsW�R����j���nE{�M[(�&HtCY$��.���E2�=�4pK�RqZ��\�
�j�(���+��ۍ�?�09���ۖ��;�b�!Ir.���(�}���hꀼ�K]���|Oڍ؞�Z�8�e�̀ⶏj%��/}5}�J�l�K��vm���Zhj�@�0���Th��D��7�U�j촎}w?/w�޼�L_Po(嫌�ȀC��O-v�����=`�,c}�	��+���ė��<����冦��_���S��İ�w��3l�4_s����j��)�̧�6�bcH)CR�Ժ��ƹp�*�c_`��T
b���7�~~��v��4�b�/�$�[K��R\]��H��a��!H6��:�o�v�J{x41��~��?-n����{A��k����E��B�>���5��ok
s�-�\p�����=L�n��.��q�T���w6�J�Ҍ�!�
��G��H�:�c�nm1�Ƿr��F�[M%�QM�"�����=�CA&b����Ǟ;��KC��ǐ(9��0��/)bs-�m?Su?��T�5�!J��s�851%���#�.Rj��J`��"�6�8�%�|��fIC&��IcHܒ�`�6�<���&o\�`a�.\�����C����Cz|�@ڗ����Ն�#7
�Չ�aoU3*�¬c� �:SY
�_(��t��=̃���x�;�$��U<�w�#̗�wZv��mY�J��W���<�Z���7�1��e������W� I�� Z��[�e'84��4�#�N��qo8��P)�DW6?��ꉸ��	އ/I�JF��IN�?��&m�u��AnU���]Γ��Q Iu
0��)��X�;�@F\�i��]�74c�x8�����������ϳ�{�5y��̤���K�:�N�b������0=ve� � �i�gJ$l	�^��'՘|9Ŗ��T�-�������	��D�Q7غ��J�#����Bp�]4�̄���sR�a�k;��š&|�(�QŔx7�q)����� �b�F�ו켻+6?i�;� *���[��{&��,iPt�U�c�D��[���9�g�[�!T��a�G�Bñո�E˛� �oi�#����0F���1����u�q�Б�E��r���r��6��Qo�2��,;VHO�iv�W�~�?y��w���Xӯ�I?g}׏�5����|&p<�M�r�����a�&�m��ˆ��WUX�j5���M��%���i5�/�4�0x��(�x�X(�I�5��;���W3���T8�MUS�0�~Q�Ф���U���������`���>Q�Cv�8
O� ak�c��_�c5��M�����z�WI���9{��\��u�p\�t�$9CԒ��n�2i��3c(ȯn������1 _����@����$�U�є ��7�c�^��-TqٻT2�Uǵ0�k�u��.a�SҼ��4m;����"ZwC�%�c� ~y	�Sb'���+Hs�{w|�5����IC���Ǖ��;�b3p���+_��7"b1�z���d��^�e?&ًL����4�_p���A�������&dsZ�v�Mjbt� ���v3e�Ǳ��2B���8�����9��X��@�%�
��x�6R}���N��-���9ʕ�����������B�
��N�/���c���Tyq�ּ�I���G�6%3r�:ڏH�t$�W���a�3���7a)oG�K��o��؁\6�1c��CMT�tN�\�v����ԛ�OT�f�fs���?A�R��@07x�*w�<C7r��$ɇee�L$�0An�	'����a��,�؁�	83\�壠-9u�^g��2�*>�'�M�y�� �cM��!ȓĝ�ǻǟ!�;~��A1�����
� ��(��9������<��w���������n3'6
8�rb]����`}qb'x�?.�|Ro�v��3X�����Q㲉�C#�d����?z�ŗ�E�@6�R�ߩ�}�1��P�-&j�-��%*�$a2/[�+_�oL=$@Vл�F;��h��5����.S����N�������H�.��D%\�*�ܦ;��|�����T*���)�S�'D�0�8c�2Ew�nQ��5\���qZ�jϧˤӟ����<�!@��(��Դ%'Κ����JE%��#����g��'�Ë2ɋ!���+I��A6�T�%p��m~2�NB�T(�x�nծ��{2�{���$�)�D%P�_�bteD���*�q&L.�@ d)+�������z̧�t��!Iad6u�V}�+6�+?:��\�� �]�{b�Я�Gv#�k���n�C�ZyD��H��
��x{rcbؠ����v�)�@M1�2�VK������9)�q�u&�~;+=9���7��I:B��C�/e����/��Ͳ-ε'�#���?�I��)^��EpV���u�Os�7XtvU�m�xU#l�?�^o&����%w�0��PC���U�dݘ�.�A��1����a���*~�k�|�5=���wT��F,�,ј�����o��;��&p��W��+��)P'�H�B3/1z�V[��	��$��
y��%(sA'E�r��h��AF����0qQͪ�w-چ�Y y�ϵS���с!=�%ۊ��*C�C��n��Q|øL:��8���	��Aé����< �B{��ҍ=x ��n<A��?9�[����	ig����$�cP���b����!��O��Ĳ��6m&hp�æ�YƳJ��dP���2�М	@�I��P��wk�z���4`�5禞Hx��p/�i`����T�Xd�d/Ν�c�٨kB�q= "d�0�B����W�#tKٔ�;�D�AtZ�4V��5@�g��!Yf���qdAN��<�Њ��x߫�a�ŗj��� L�/r�Py�y���>6f�������*�𸢳�Y�>1����9�W��z[�0X"���蓓;�\�S�ow���h��� v�"�� ��+�_���7
ۼ��#�'�u^���N��-P 5L��w�ԾP�eҖ׿*��pW�>� �3�,�#��%)���W6?'���)�t���@�\��kS�G��wR���S�@����RV���/�18z�}q݆�*�_���i�Z��v���R����Nc˅�~�Sfy�* ��j�ء�e"gZg3j폒��&�!a%��[��zK���ꏴ2�|k�\��3��"��;D{S"H`S�4"��*���_~��CNǍ�qp�6:�g����Nڜd��8O��\�4^���k��y�׭����U�}��4��ג2n��枞ꄒ�Z|��P.��E��9yn���,J8�tଫq��iuW����ov�#3��|��Y4v(���b�Hz$�m����a�t!���Pw���ǡl����*썝� �}�NK�i9�]O���!3�W��G�y�MH�x0��a�?RY���x8������Y�fռe�Y`F7}GశZ�Y�����?��8��#޾]�|Są��)�t�%�x)Nu/�B=� ,��C��X����S�Vy�\�l�
p�Op�ͦʩ��(z����`�D��	ԒWD0�_"S*]�Lx��')g�YnG���mçLSc$B���`��F�@�^Vݪ�z�-LD�oInK^�6"�|@X���dJ�ZW��y~P����*�@B���+��Pms�;?B����͡+�"]G�--b��Ez�ӽ�lƠ6hi�\m�0_����k�1�eK��NW�ׇv]@��)���B��k�o�!���#��y��3ʦ�(�_l�^�<m���n�2[����l>'�y�ʲ�u�V$�}ް%1L<�����֪!��<�?Q8f��8uu<8"/�dW{�5�g����p.�k�O�ӕ��>��$�L�Va�2��������E���T�!Y��ѕ��ϯ�i�v��y�ӚQ�'�-5�TQ̓!���wa���~�E�?���{C�ɑ{!zkG��SS���a�%A�P�qU�p�W�<v�yk�����AU���1%�� ʖ����nDK��+`t��dt���q<Z� ZqP��j�t��uڑ`V���-�|��v~40�X�v&����{P��'�H��9o�a���z���A����u�Z�.55)������O���ݩ ǋ�/[��!�B� �5^U怢9z�H<lR����l?A����H5��� ��[Ad>=H��|��	o?hя*����\�5�%H�%�B�	͌߭�ujNyIL,���!^zX
4����VV"�!�DL����*�3��r&�^0�~~���=���"<��3�q1fk��Ǎ�g7[��,�����^	)����ڳߊ��~gW$�=���Q\�Уh�ڗ+R��;
Q��C@[.�'�����S��n�12�v��,��G�ߑ�H�<�`��w�Е��"�5
j�P��_cb�W)i:��Nج��5�5���&\U�Ʋ�ʒq�U)�s�?a����פd���N�WGʿK���A���ر�/}G}9�	����`��^<�j؀��%�ߍ��i�����wFx%�t'��]��(�	�kun��U�5Y�Ts��`"�@���v��3�r�L�:��a�&y���n���uPW��!
�gd�B�EG��f�a��M���a�t��h�_t�+,�Ih����G�63�9Ņ��>%�������[�X3���� �CkS=l���NvA'c%�9X7��:���&���~�@��Y��R���P����َ�S�X��!�C��BM��T�S:��)-��9߼�HEO��� =K��+�^�ag6%����e~c�}$�����f�y�ڑfp��L�~B�f,ǫ7%�~�7T}c����8��	0������Lr�J�}�"�P�N+�&� ɨڬOl� !E��v(��+,%��cA���ߑJO3����31}l��!��u��M�ѡA`�s'�\���\ñֈ�ػ&��{�~K;�P��P8��p+�]����9��PH�QC	NO�S#�}�*�zȖ���Ts~;`�OU��ۢ�]��r������$��p�Ãm���s��_dR���1��^���գ�7�؄="�JFj.\�a���ă�eM� ��[����=�dc�<�&ͷ��q���;ne�����X�Em�N�`܌���)o2k����8aHH�̡2�d������8x��u�6'���"L�[
��lʵc�0.�;6��+ ,V���ԧ&M-$�ٽ��[�q�F-����l����m����r�e���[*��Jp�B5�zt�"{�Z���'�p%��J��G�c�Z�-鷂�����b��e��3�W�{��߄����^y������x~Q���8�s�k�� 5Y:�k���'���֛�h���C��Q� �*i�7S�R��̆T���:��$B�Z�Nk@�8ªoJޝo�����W�y&2t"�| �N�+�Mf��I�uSsTC��~z:���
�r� �U >�P(��S�~D�-�/��hC�6�<�[r >���o��d�+/�;%�xS��znKX���h����2�̝R��i|�X���E�0+zc�E�մ�{���ke����֕>�M�q��%{�>]S��[����u�	���Z18�PM�BV�yz㏼�X8q�j
�����2 L@*��$�O�p�L�����%���NbN=�����
_\�џ��axZ��k;⾼���`v���3�<�1gս���d=��Uc�Щ�i���N��%~�ž���K:��Š}:I��V�U,G�b]��9����t}�(4�����ʐƮ�'��Eخ���C����3>M;�-����q�׺L��B�}O�2�?��i�l�az�!�Q���Oğ3�TY���m�<�T�j�kj`k6�[���\��]l(�1�N y�؇B��p��� ,��/3�B2��	�-.��V����韽4آ��*E�d�A��ے����p���oJ{V J{I!¡��tKx��s��	
���6:h��p��r�̯7�cT��L��;+�SmR!����׼�������]��0�W�z%�`�ctw�������{AO�i�G�sԁ.=�I�w�+����'���(�Z�a��7"_��]��PzQ$�"�I���̸���b����KT�}D�떙���Ag�}����0?����|EQF�|̐(���U����ô��o5��7�'������I��/ͅ9�v/���<�@�k�S��g#v5V�x�h,�t�>2w��������$bZVb�_0<���{��K��Ftj#�Zx�9ow�)����dR3l�����6�'��&-ߺF��;¶w�_�J?� �C`��M�Oܽ��A�����F�5�Xѥ�b�Dn?M��Pp��K�� �y�"P�պ�Q?㥳&�̿��KAگ�P�n�&�Cn�X3�A�����t��/�/|m�GhA_ Ԕ׋�j�L��@i2��1���B����(�hF���3/���Ǭ��a~�����Cd �aa�� ���k���+��;�U���7��_=+m��:��r)ad����L�T�wf�Qb�!�ǔ�y>!
����fL�N��Oݡ�r���A����_]�::O��@?&D�{��Ν�(�%���_�*]*��]���_��:-�;����&��:(��ݩm�@]�l�t�
���2}���[�P%#�5yw��ё�it�\C�#���0�G���׿Ó�r�l�!�5����}>�����iڐ���D�Q
Hu%Zp�ܤ�>6��������R�(]�H���GqKtwX���of`��#�(�ev�dR|�;0XX�lP� �H�N�>zF�STD�����w�`�hGl?(���^-3�ܡ8���:&�6�[)4��y�d>��[�ei�.��cT��pF}�/�ep�.�G��*�����7 ���+bG�UΫ��[VGR����~i���/���X�n��;ٿ�t�(�J��s	yw��Aі�՘�'�0Zo�S� � \�Gu��GW%S�K������F��*�^�� �	��L���E��� 6sHrV3�8;��H"Wߎ��q�ߒ] ào�?b/�О��x�C���K�"����X~ �)���'�d��Dc�h�dV�>��C�=����KU�9[���I��T���3]]0�.�@�U�*=��b��
_����Bb�	D3����(g�R����ܐ�K�!8fส���3��o�0�Z��6���&s�+V F�"fk����DGh��O���Gɦ33����Nc�FZ�|c���L�O����	��:$�J��{*B�:�%bNH,������6����2�������.�����>h�E�A_�zE�6�,�̨3����d1��- c�b�ב��r>�������g��F��em�u�:��Lrhy����l��������ĝ?��J��{�t�Pn����R�� ��v�Ɯ�#� ���,��;i�^��^�罘�(���]�"�C<hS�3�z����}�j�A���ߑ�Ѯ:��m��o��w��^p<W%a�븷d��*���Z�$*�ӽ��������LJ�\�`3������1
P��)��tu�"݂�E�����s�iޠPdc9��T��j��@���V�T�4����,���\q3[϶�����O(p�P�ׇXVY%����z��ܦy>��'��Q�m���O�y��Þ�&p~�)�*��mw\�A�;G��]Z�ܭ�4���xj�
hm�D�'�n˰D� 	��u��/�F�����};�
�7��:#E�BZ�Q�[=��mV�9��Е�����ȓ�3(fZ��v;��#��d�T�7<�h�� ��	��o��}�h�<!'�N��C�"1�W#Gq�
��z#�n~5�i��ʞ�{�G�edϱ!�b�P��7�)ڹ��9����s�e+��P��M	'�E ��t�%t�:�VFU?�AzaNA�g 6�3M�U��i���.x���-@4�Nt����v���}���Q�D>kX�lؙȁ��}�7{t݋zሑ���d�l�8��%�9ʦS����$�������m�G?P�� �iT����?=+%ſ����0��dR�L���ڮB������!�¼����;oPdj2��ɱteūg��FZ7Co�AC��rfX\@X���`
{���K��&{�n���%�J�f��Ӭ|�N�3�:�N�
�Z��A{+�HT(^�b0�y�25鮰I�;|�2ƒ��'Xl?��@��,<�d�U�袖�R��r�H�ț���/�:�cO���9���_?���˻e���A�-m|u��bW�.���/M�Ɩ/*?�{�8��"GWI`;L��g��2�fe��H����[�N+#���l����x�5�vVM��L��+;�Or�}�]�8Ԭ�������{��3
��T�e!IR�_?ܴ�L��Mn'��dD�D�6��ŭ!۬�����9X)����8��1��w([R����S��b���	3Ǒ�Z��;x�ը�_2G����y������	������ㅟ���ƚd�L8&a@�e��C���R_��=�� x�r+Q9�S��� �&�S��T��PC�G��~)��Rz=�ǋ#�.o+X�?Jd� �����tz��z��ӯ���ځ��'m)��U�,���f����O�ϢkL8���'��4���Q騙f�3iiS���m?t��"yV�,�v����V���?t��$������K���e.��>��K��̀{��/��eI(���|�+�`��3V+d�~��@V�>VT�z[�v�2�
ߴ4EY��Cg���$�c���{�v�&q�m�̬�EN'�i��|��� �A�ѫ�_�hK�ύ}wP��8��	@��n6D���N�ӣ�F��{֟
��B�r�OI���VQ3+���g6���+��cp��v�|"�	��y�U�R�H���Ϻ=�W�D��
j�
Q�ru��PKHg���E��/ط!�0<˧[�z�QI�zǂ�Z:�6&�����X.�ʲ�5�ѝY����t�F�C��*��2u���[���/%����|v#�q���{�k(��ū���!�-u�Dh�6�;�TD�2�&�l�sr2��Τ����#ٜ���a�U-V����r(�Z�$�	d���b���{��>����(9��X��|\]
���x�CAҌZH���0BX�ŭ@")��"�3�c��h3�2��o���ן8�3����+?#��b[~k�v5	WĠ�Đ4��x�0(!������ˋ5[�l�t�&��J�ʺ	�ܮ��,Ӭs&���w8��HaaA�:F`@��4r'������נ�9�G��$d���n��V�4����W������_9J��ZeDHs�oo���ހbe]��|�5+�X�~}��Oܦ�?>�o�r0�Wa�4��6�}�$�PE�I=?v,k�2��}��ɒ��i(�����3Z�����Zќ�' ��B,����u����]2P���Mv�Đv�[y/��@|�<��������Uj<dh|���9Y�^�4
�+u@�yt�2�m��C���r����r��
���.�T���,�Sd+xo�ޚ6]���DxX�쉀Ukg�
��\����'�ԁ�ߧ�������^ �V�K�&�Y��F���p��gp��S�hLw��R�Ǌ>̕o� ڥ8���� v��"|g�}�T����_��M�%���F��)>22]ؐ�(��z��W�vcA;#|ȧɒtȶKj��<���	Yme��b��`b�4�t�ǩ3���Z��t��(1��J�� ��	d����Lȇ�\�3������2���-���k�p����&��1x(Mկ\a��4��E�����?o4S��y�0�x`]�Ǿ���9���7�<�d0l:��R��[< @-ǶI�+@�0F�vH0�u����D-��c2ck76R�<����ͫQ(����o��	�GA�#���3�4�Ħ�i��4NgI�m� P�����{�b��@d3�;yx�ٝ,&#�/u��$��l�o��%H<�S�i�K�M�}�C� �N=�tg"������㯮�l&��MA��!J��M/Cj�#��f�Z&� ]�$��E # �:f�� ��|P�v�z�dO����J��z"���q��L�]��t
 �ʪn�Lv��HaD�8$>�>�S�xӎ�9�ئu����MTA��V�����?@S��= � �--:�(2��u
r� �';���1;48V~��Q��wI�S���V��@7R�!�"����k!�.��j�ezN�'V��AP��\�80*2��c������/M�ө1�v���/���!s&g�9���H� �	a�kQi!h�4�fe�y	l���3v�]kZ���^��ܪ�V�u��B�R�iM�{׽���w4�,���imGZ�U�uHW�D]�a[�r_���q�$�����E8di������jѐ�s5�fȹ�<��'sA�Vi,�V��0Yi� ��}S������L��<�\/���� �\�<gG��̸�LB �z��B[�]{&��?��*��*P��Fs����4+���)h Y8:(0}"�܎�͌���FD-X����0�g�Rx~���^��9[m�C���˄o��4:��rC�<��.��;ؾ��j�?�ަ[����N$0qp��y�*+�o��+�/�F_BTn$�Dp�P��;�������^��к��?��"���b��cJ#Ukq-����������\�@Ys�_�$�x�atO�c>\\�Ӛ�҄\0��U�M^�'0�)hB'@%��D,����P����R��֧�`�ۈT�I���,�.����#��=و�ĭ�x�>|V5�1�p5)[��,1N6�W������:#(��%��0_*��n�섄�W�VVUM���u|��Ne
.I���Ǩ�\�$5���E1�3�b�_�sL{�%y����Q���C���e'��	�����ݟ�i$������L�aQ,�ˢꘗ,Χ6f3�^Hҗ�<g@���fW�ZsYD��<N���l��	���k��a��:�ɟ�]�~��	l��#ϰ�N��J��	nm/��/Ӟ�*���iu��<w=���2�jqB$��8��8���)�2P�S�_���_�2f�5�@M���v�bG��:�����8Y�SЗ��O�*a�dz4�(�&
CW�`݁ �x*�M�u�R��A�+�k�Wټ��"G5�~����	�g#�ӟ�@�Vj ���H�0OJ�0,����W��dAIJ��)��m��~~B��\�у\�d���U���5���KR���ŴJ"�J�:AB�V���A�;�LS�9�{j�W��	��+�b�ZI�0i��bP����4�M�㖽���rviM��K��k�c��?,���|����1����Q�R��DO����s(�K���X��r�}s��ތ �����X�dx5=��wR�5���Z�xfE�&U?��m�?�	����`Y����~��VB�3�Za�����L�07��U2{<�!!e�ɋ>oi���`�P2_��a�,��c}��?�&�R��9
����q��G�����]����_\�����0�X��)F��N��в��-}�RM�o�>�Ӭ�-9���N~��jC�>�2�74�����i,��C�ޓCZ ����T�<�����,lQ Z9�,�l����4j�1r7R����|�����/b���{ƙ�w�����.!$�<V&t�Z5'&�v���^&�l\v!�J���^��̪� z���\T)>�s�v~<��ô�Q���wEJ"cA��]��7y�ң@�P�8Z�/(!(5�4<:�;�n�ی����|j�))v#�;c&5Y�&�kߙ2Y@��1�����B<Gw�(�����c�N�4u����rE1������\�m�(e��m���u5�A^�ğ��i�̺>����r|�9q�5��D3}}��3�d�>����x��!E�ϲ'���ZA�h0��\�a=d9�4���6�Gm�n������>���|�9� �f�-Ƒ�����$Fd
��G2(�X�|gW�gS&������ڔ���w���q��Ŀ��kh>�����F�S�^{뭠α���
z߫��3�\� �~����_��U����I����)�J�!ٟ�XN@S9���8��5�¼xr�6�������~���!�Ǥ�J4ޝ���nq&�ud��M;���ݩ�������ȁ۵0�������/)�OX���K	����2o}cm�� �^Z�����, �p8(�&7R&��o.^����B%�9� E��
���
�H�[�Î����A)	aY��k��L��U�1�����	��{�"U���z��xm�� F���B��M	��ܜ���A����[��@å�<��낢[�Y���t"�v������0-w8���5�, �{�gHLfA~���̯��J��x�ߦ���R��k�c?�xB1���h^̻�7wad����BL�K�M�E�'�I��r��icNn)����u^}d,XCm�c���R�,�����FX�Q@�/
\���(�*|_h�c c2���Ϻ��`@���.�t|��?�� �T;x��=!����Lų:R�=g�ض٥�/��wD6L�M�1I��
;��TK^��*V\� ��0p��p��o����{M�WL(�{5���gkZ���s;i��}�W7G��{�~�,�m����\���gxqyL�N�`�KsX���jn�>k� �G����g^jT�gȀ��� ����FH0�q9����F��L]�'y$Q�B;F�@%\,��+Śq{s�dG2fX{��ئl�g�c���l�s������E�i9!�!�c����f�vyZJ=�Z}�����C5W�r)�OXu<���ؙ���)�F'����[B�ra�
p%�=�F���?�rŝo^R�@�*g{ܖ�2�ntn#��m%Y&��G�i�L{_5a���SG�H��E��G��r���?�m��X梥ޅ�}XM�EM�$Sʹ��ey�_��E�W�d�XJ<���ቧ���ş6�f����V�?Z����!P뽧�$i��$q��ϑ�b�2d�F�U7m{�����'������%g+��W\���4�����+T\g�]��xN}U��#[�Aj��RHK�>���b���Z��ޤu��_@�����ӮV��!���N�WTkNH��q��ց?��D��(D�(M��jR���5�9�"�>T�d��{p�r&��Z_��K�8��@3��b�����V�X�N@���}�J���n�I��8�J%uV��&���L��s�YU��f�%��l�X�� �.;�Mg(8���R����R�ו�0���L%�� ���4n�ؚ�)��/�F�C��4|�rQ�qO10��Ⱥ)�@v�\��U~�Aw�7�-�[@�6+�uP�>�!OYu��N&�,��kE"�$���F�Ԃ� #��m��ֺY��*R��*-�j4�UqZ<�e��A��f��r������7�7����a_��t:�7�*M*bYY2��]h����� ��3��2�W�bc�"ΌC���z@_g��ϗSq�I�]�`�R@�l��!\mP�dBu?b�u�&b�y��Ϋ��n��i�����Z֘?$��!����o<F�<d��X�Ż�!�����U�Cb�����c��"v�KLMUb߷�}�ruRAN��e?s8X���@g�����<3�(���'i��	(-*$<!�A	�}@�����`�t��L�O�f�	�Jo���d��i!�ux��������*��	0�zU�7�����1�)�na6�5t��������}$�"���s;&qZ)h�t�AAE�X�n��0���~�`L�bX��c�;�c3_����<lْ�?�F�\,�$�;,�?��@*ʾ�@�)[����%������'3ik.KW���F/����V�"z��� ,W����߄.gn�X��$<v�y	�\k��AVz��&�(�ΩO+�'�î*��]�0�E���[�g[�,M#�m��~^D�t�X�($���_���,2�!��	t��M�o�G+�N� �Z������;:�`�,�JŤT����k��v�u�.�hqќ���4]flE֒�hk�2�Tkz�~���6��V��n5��&k�6��V
/�s�Jߑ�ںˁ�<|�K9*,ץ|���CV�c�\d�����7����*��)��Zt��-��:���X���L��r� %�Q}	�$Ӆap�KR�2��X�>o����k�%�U8W�+I�F��E9t�<�O�� j��Y�����)��������1����i{w�|����^�
�%�4���4��أY�n���� ���L���W��* �^&_��G�+04�ل�e��ܜ��c���I7�
<����U��l�7~�@t�����r��ٚw�C5+��1Y����<gG��Y�T�+LI2~;�� ���˻����N!O�҅:��
28��O߅=�EY�B*�;�p�< Z�&�#c|��<�Q���r�O����O(��2�ʜ2v ��ƉW���q�eMp�;6��8t�'��(�_kɃ��DOfE6£���14{���+�^�>>U��P'UJ�K_C� �����m��f�j���=��l��������5L����w�^ˑ���?�����oz���E��q�;ؠ��X~ÖҮG�)�$�*���s�n�y��H��I��V�'*ō���1OB�g�3I��Ƌ�h�F�Kx"�BEa5ͽ(_k��<�{d6�O4c{�� JDe�\�Iao�c�>��E�v-�y쨫�Z@��=J�Ȫ�$L&\��W�W)��L"�Ē��� �B�j�P|�A� ]耻���|VX��z4��{�]�������wl��[UH��3߼K�E����kԎ�2	�O�����C?���HC'�L�S��P�Z�-�k1�����q��^I�X���N.����<�"�~��$7��V�7;��Yݯ� )�_4�-؎4����V^Y3�t��b~Uɨ~��<��6./��à b��4����Wh��"�?Q�иWQ���yo0����<�6�t����e��[m�m[�(w=�C�R��o�.�-�H�`k���73���G��bQ�4u�iU����!��Py|�ix�I�>R��-��o1t��*�0݈�0�N�
�FM�R�����\r�9�Z��h��g�A�g�l8���g���!����"�:.<�6:�JJ�b_�r��(�-�U&�/G��!��DDl>����S��$�׵�$�TQ�8�ûo_�b�<�_����s�Lq��br1w	e��ꡩ��E}���ց>�Ȭ�E�뉺������������Ń�dHMH�:�;5IC+��ۉ�^E�ȒW-.�sv9�<����������;�8��j���l!).N	�w���W���� ���5@{�s�`�� ���SXW�w�j�6��?�P��� `l��s�O?U��H;L���P֋+����YS|az��Ϧ0���{xw8�����t���y+�|͝8e��~� �g���}���\"�`�;L
c��ۖJ��z	2�����Ф�ҏ{Ԕ;���*�Y|&K��v�c0hnd�`O	���p����jn��&��g���X�����p
H!��go@���`�n�T���3��_TR2�y��s|E|LӌВ���;�}�0)�J�Ӱ00?u0�@����S�#&�}�Bŝr �(�d������_0%W����;�^S����������X_��Ф&Y��|Ix�.�=!�|�~o,欮o����9'U��R��h�G2������~>
� ��9Ӱ�XgJ=϶�����Z�$B�׫q��	:���/�+G����iq0!=1̮cz ��Σu�����9HJ��t�z�o���/�����������O���FT.㩪�?�0��I#ʮl�)ɠml`d�յud	�%���*	�Y��J=B���O��2V;r��k��R��qb�@M�0H� ��ѻ�)Z�pǧ������p34�1��Q�rݪ3쭯 �Q~�r0�����E�C�]���AEet�C�idrÞG6�������W���9n��̄e�GGj�6ոxV�B����Z�Y���x	d��wX�����Ý�x� ��~Vk|Ƴ:����!�83���u�k�eЁ~҇���d%җT�CD:.�*t=V�:X������=:���Q���"�'�AtVr�`1��P�c�')qΠ�,XR562&��Ɋ�ۀj���)�~P��OH�ȇ���EHZ#�J[]P��a���݃e�Z~` 0�i��l���"Ib���=�O3s�*�OcP�(+7v�suh�ZV��R�4"��}�ÄUz���I��.��4�{�'�{~�w���z׽��c$Z��׬n�`�ڟ��G֍{�ya*O0�Ѻ޺��wzF_Gh��Tu�B=�@�l~ D��}�To/Fh��`����MG�5��5���ƥ�+�ɥ����R�Ί�. c�n�?�?ۊx���Ϩ�}����R
��Ҙ�ϊ��U#H�� ���h�����dM�$�),������`���"�Isи���t�~�|���3�
;'��2�GV��pM-�!P�S�$�w+�<�?��S(C�813@�Mk�Gh�V�i��~C>�$XsP8��������m ifT��C���_]��3W	6츱j�A|�tF�+^V�:T�5gg�.��{��8k�"�Շ��=6�O��2�~������U;桟Y��<+�e�׽CHx�G�Һ�G���Ab�0�I$��^��+nԈ�W3�k ��CL�y�[���b�����A���3}��"�N�U��jZ�n�A@ͱ]��=��b��f��'V�֒��&+�0��@$]��*�7e�.�W�����?�Ӟ�(�|�P�6��	<(��^ �O�\�G׉ R[�=
w�A����mm�VPi�h&9$a�M8.���߲`�����Ki��*�5�?!��7�.�)�ӫ]G����-bl�.D}��	����y6�Y"�BzvYt�ߠ��t��PX8��K8��C�!B̼q��	6=�J�G'V��ۘ�?�����2O?��L8��>����$��B{��__��Ku�����^��"�o~Y�8�� ��ߔ��nq�/rR���-7�&�)}�xj��s ��!Z;W��y��[�}�*�2� J2�����0Tu}<�z~�"H����IX�R1�UK�,q�s����W^�8���
(���y"��t\TOF_���$�kSx�9�2����d���q��4��|��Y�I�J��UL�m�ю2��
�n���Ch�}�'���՘О�\HB_�wY/�*Ք�Jjk� ˝�թF��o�Ȧ��3�I�AQ�������25�W�D�'�i��4D�D�wsg��O��߽f�����[w(O��{w��e�Ns��F������T}џ}Dpe��_��ģ���� ��Us�!*�L�ޡY0�仰	�J]�E�4�p"=��W+C��f�O@ަ�'ˊk)M�����}�A������<EE?02cOc��D��x/"h�`C�5�B)jYL�7ٌ��(���rs�����M��b��_&9�%�F��=s����������|�LaN���!`��;�١�4f(��ݠL�!mٛ+��;ĥ�ⴈ@8�3}W��Hǵ�'+�ݫ���/xhn&��ќf�lJ�33�b�jױ��E(v˯�v�D�{�L�������g]�:no��+�c���Q<ӹU�-ɠTT�(Y�'2�?*}H������9*�@���X�|F�^_�}ۊć�YR��5��ô��Ǖ�L*)Z��zbz�^�7�(@�3�ebe����[���0�z9qwو?ƊQ�XZ���r�\�G���?f;�(�C��\����n4��tw�.��.�#|�$0�=BZ%ܒ~x&��_F���ca��#8XY�E{�z$m������C�\��^"���0	���mB�"�0�4���|����ܫ[���M���>����$]��΋��t��b^�5�-�r�)yתv���\�Իn����Fިz��
�[�OV2��x�w��C���Í'ݐ�U�߯�h3�é��T�'����ګ$�4)������P�{Z.�3\DÈ�]���]�M�>�6��澃f�
��3�����j|X�.X�����)��� ���ޅ+�ȣ�fJ��*<��oW�c���(�G�Y�j�=?���U=[�yr����]��U>(�4���#�Z���ی� U�z�Y��#0�=g��T�F�ք�Yy�;���(��J�Lo�t�kJ?QF6���5J�9���^�e�t��HM=P۰B�<�^���RvW�j{�GI`+=��Ƌl�B��7#�"Ə+�c���4��V0Y�GN�����q�;?H�Yr�<9�㥉��Φ\U�?�\e��\>������л��y��s��0WǊ� k!�*Unp�=)�7u~�$N��z^W�G`9��u���!ׅ����������D� ?zK�k(�I��_�\&��f���G2��x��Q;��{�-�Ouwl�V��W��gY/?�G���s�'Һ)r�z����K@����A��X���O^��|_����	����ݐ~�� Ԃ���R;~���E/A(睈!r
ݬe%�TCt��B6P}�~���P���3'�,�u��+p-�R�ݗ���u�#����I�D�̷�,�STz9D�
7XRr��Z��P9�� w젌��_�BE��~ґ�˪�{�[����؋�� ��+�i��(���w�g������Mj�N �<�� ��m�N=����/ihkJZY�Q��XT+��~1�ߨ�֭���'�ƠO�Lh�"�^g�E}��-���7�:uI�l�^ѧ�3o�*����-��&�� d�čt(zCp���б	�t�����r2� ��k�J@�)�^��Gt�_��|E��@d!A�+�{}?FL��յ����b�S�'MS�wzH����H�"AKحGT����f��S�Z/��elQw������mu����+`4�p���wN�l����<�~�u���/Z0K�Eo��l}p�cbnj�uT[T����VIS���|1�ڔN��o�7�ӫ��"��o�j���a7Y��U���*wXU"7B�0���� Կ��ҋ����w߀�� ��P�.�ϋ���:s�N�㚉�6�qo��4�Y�	�W,��x�����^\�%�;�U��}�^:d>h�OH%aV6���ɕmy���2�1�*����ء����x�տa���Κ��OޅbS���;@�%�5�T����-fO})դSe�5�{���9]T�D�s@����6y��kjE�Ԍ�K��֊��9n�[�?B���� ���ڰYR"yX̶�Y{D��r��D�8��x �%��¬����UЀ#a����2��>E(��OI+�#�S�y��(B[#�����k8��Z'�B��a���<�\e�?��R�Qi���6�們�?�+Q���[���
���/�>�|�խ;�(�l������M��\`��y�*��e#���H���+����i��J-KKҡ�2	=f���<���]D��������	��2^��y{��� �9z�L�ߧ�z�j���@�Ɲ��~p�h�m5�d]΢�|�����[d���D��EZh�-����V+���6��]}�>�nߵ,?�`r�Å����@4/g})ݲ׏��-��K����=t��'(쒭/��F�g�q��!�����=�(`$ȧ�Kw�[�y(c��U��B��!���~܈��\�!�!�������IG�,p �i���`�FX$�F}|@��< ����V��� �H��%�ڙ�A���ŕ'r�J����+E��☃�C�w}DY|�(��!�� ��iP4�Z���x��&�d��c�ƇF��N�ܝ�z�M�^nj�"� �, Y*��>�$���:���ewe}�k�g{̣j�y�I*��%��H4��lik�Ɍը^�e%g'���-�R�|�,�L�S��-ն��p;C�tH���<:���L@�V�Ը3�0���U�>i^۳9�BCÒO��p�Orc�z������Ʈ�!�39��Y������pT\��Y���"x��p����� �S��d���{!�UxF)ǃ���b�B��)1���!��~�M�֝���oHfZ�e��K���.|n��M����xt�C� u��C+���m�7��Z��\��(i��B~��������[�!�Hӆe.�(�LyV��/n�'Mׄ`0���L��C���m�����[��~��a/��d.CQ��ٷI+.DG��
~�GJJ��<��K��$"���������A����_��������$��}�e`	�x���0E��G:�E16B�̙^\��̎��S�zm����'���.�u�y��3�Ѫ�G��'�F�yo�9c:x�˟���"����O΄s8�}si���
����7�d1k*В.���M-`W׀��E��}}��s���]8�I���Λ�Ӹ����@����g�K�Qc�#�Z·����Ϗ.�}h] Q�氍���v�/�8�cS'�{}ف;[_��ͯ��Zd�-1)�o�����L�{
h�wp��0C�d��d�\e���ͩgU����������C�xqyΰn�t�Yn~-�ϔZTƚ!�o�_����E�iq��N�)��L�	��=�6�!�mV�����M���EZ�>��̇�H+��K�����~���U$�����ǩ8#�ڔ�W�Җ$���"8��A�GK9�!_x�x��θ[����Ǹ�I��] Sjy]F�\�������g����M�>�ȶ�m)B[�K��/t����ȹ��c	����筏J��t~UøA�2����$k�����-� �٢�ݾ�װ@�����GI�/��4�S��qA�'����NWFnۚv����0e<���ni��SaQ���*�ϭ<鋱}l��]|Q�R٣���A�	LkG�����֑[���&�/��6���.�s�{��f��;������n���"\�/P��9+��c3_�F���Jd�ZG�9}u�:#ۭ�'�G�QT����fp$��h�h��
.N�̨�h�� 's�27W���y�11��"ԃ�49p�B�"�ݼ����Lj}�l�~W��v��/�jFD���dg+��s���k�ӣ,Ņz\����?��Q۞�r��=��������j�Yv��i��t*�h��w0��������&�+D݃h��ܤj��o��-HN�â�!s��7D���VY!�|����l��&s"1�~��ߥ򮁼-�&-_g6I����aT�7V�+�d"{�rq����	��C�	U��*f/x��@�;���.�>ԉ(�^7�]Z�|����&*"o;#��Q�R��H�wz���֍G�5C-dr�n�2Z���� ��x���W|�c���"�}����+�}T pن�{ ����/�܏��]m?>�g��g ��ch���U���q��a��x{�I�w��D�f�!F�i���rثǁÇ����9�?Q��Uqܩ�ltX置5�LsZWM�� m�}8ZrE���^�Er}d��	X1�\�P~(|���B��y���"�3�X�hm�훰G�R_��I�اA͖<�[�����1�{�^������Z��K]쫑G�r��J��ѯ��4��~�x�u23Sy��Z@�2������N��
���t<�v�~V��yo�?�����J��۩�j�2j��c�A&q$�M���K��W*��Y��S�[������OK��{EE�y��C�c����M��OI��<��P�^8	�f��]�<퍅�1����*�D���'w� U�ԗg�.��ԩᘒi�?+���B� 9�K�9���l�v-��r�w�z ��/{�X����!;Ę�t���g&�R�����N�n����^�-��>��2_�;h�g�������f� ų�F�ש��_ʸ��kD���t�pDp-y1S�Y`K�i�lu#��p�}��Ŀ�����y7?H0z�R�↸�,1H�=�5�d��#�C"g��]��۴쾅?*b�_Ʈ+˞�;�H���v/�К	�����A��V�(�\�5u����s໾0<t��X`2I�B"�~���6�.�����*����M�͔��rzj%�]Q_���ĒR4H�����K���"�F��:8F3����̴�lf�S�k��j@��;&����fH�,O:�@�k� ���~;�qmA�v��`֌��%[R�9R_�@m�	s��^ ����+��R�U�١"?�A[e������}Y���r���1�\�t��&���x �;��_FV5{�iڹ]מ�/�Gc�P��&��[e�9�����+ۃ���.�y�)i��uF�s�ڰT��Y�B�9�uѪ�[O����*vx��1x򯛘I�.>0=-�.=m��S���Hޔ���:&V��O��Q������V-(���%�XaR`���r0�(�H�M+)V�Ⱥ,Ճ��y1���F0F������T�vM7�X�R5?f�"�J�������>%����eg|�Gq���q䓽Z�V�z�cG��O�u�܍ڪ<Y׍h�y�KK��=��*7{�����[���~8)����Sm^ѓ7%��a�\��lf��&b|X��Y[�3��3�W�T�F��i���T�	�h��ş��Q�F���wBR�:�G�Oa�U�V#bg� ��Ƌ�BςC=f�5�n&�!\K����ۈ���ќ�/��Q��C���k�[&�� c�2f� ��Y&��X@�)��C9�h6�`q6�3�Jc�f(g��Q8�L�y��� l׈�;J�j�S�Su�~wX�_}O��'�^�i��=.��#�� y��}���wjx��R�H��_'�Ó����oq�qSn��(8�i��0|�]����$�ȖF^��h�=�}��T��N��h1Y&~Ѻc�K)Q/��5n�ަi���N7�_O&�Wy��=�#�L���ɮI���g>XIu�8xt[J��^/�ÿ�迿y��$�ԶZW�ɒ�S:E�i֛K���q�yC�@Q�?�>jh�'��C�bL�,�ڂG#�s��S���B�w� 0�^&w�ə�	?4�`8� E�|�Eu�4��j��l��s������%�<@όub�T��i����:���e���.Р5����\�TS\��M@����_�{q�Q9��q����y��ϕɧ`� ,�wQ7���kQ���T�K�5���I��1}��=A�H���ݤ���$Q���#�`՘���G�0��-{�|v��I=6-�gq>�ap�XS��/�l;�
N�~��{��f�7�)�{�V�hEϗ8J�Hh9Y��T��p��6|aM;���f���	����L��~��:#[O�Sq'xA���)���g=�n%����x�Ǘ��*IHJW`!#�@�\��\�
��&�q�	��������=���EL�+�'H�:p�pR�YDl):�+����&ObWu�+��jɆ�݅Q�������^�rnF��������6�
��'�5!��0�rJwyz�岼�!k���|�.��#5#��r�ݱl�mG�ݵ'������+g�����2[��b�u{)����0�-�<h�m�A��Kr�罹*��͔·��0�v؂f���[�>r9�%=�����Q\�z�\i �f�'5���!���?@{?�?q����.��C|{��\)9�ҝ�p.�G��R�|��b����^њ�8'C����X́����,_kKC7?,	�aA^2�Эo�2���N�a��C��>������l�ҕjn�3K��&e����-t�<���\/�,;���'��˥��ߔ�:�}>�[`3�C��!��b���2û�<�~��|��_��n�v\(��ed��{*��ٓ��gn�+ }�����Mq��3���S�v��Y�O98�YsF`���~���.���=��W�J�<OPs<��E���˼U|��]#��>�Ww��w�O��{�x]���~1��8����[S�w7��z�	������(b�)����K�1��(��.��]��k���荷��i�y��H�ǛB�j
��R��%P`��Jn:�+_�K�X�[��c��cnx���X��U�I���D��wg���z����D����9[��`�|�q�	2��)Q�f\��CD0J�\<�� �V�n�!��<�$���˷���4!�tQ"���.|�~uo�¿|)��)2ұ�+ΌKI�}�O�?��I}"�s�k�$�P�Kr�������#��y;FQ�GP��
]�Q
�<O������>(�v�9���7$��it�TR�@gt=xˏ��B����_*�j�o4�LYK~�� ��fMq��2<ÐH�mfk^�(ğā�bᢖ�Ȱ��x���U�'?�g��
�}B�@7��[\\�O�@����8�m���5����0�ze�lk�0s-��@�}b�������߮)�/,͒��R�̈�0�Jjr}�(��L����-]+��1�{����O.C��]�-W�wF	%26����;�#�B�*�jĻt�\[n}}e3��Qg��
�cF�\k$:�,�+=�E�#岃Ҥ�д��Rڢ�		��� 9&`�ش�V�R'Ơ.C���	��X(�5�[]�}\o�\��XԱW.�)��n��>t������5�_1,���e�]�
ho�kUy��#�Y�Ƃ�\��1��DI_�!�,j�[�j�Y�+bq�Ëw��(.'rs�:qL�Y@�,~rJJ�k�X�\Vi�Y�saL�����f8�;Aad�#Hґ�IJ�wk��?p�bj�cq���i��_�u5���0���c0���,�����x
z�ڱ�<zm�q�!�yG,´��(��.p��Na�J��'�:��Qu�/a-��/r0�1�1,ԉ����]c�ϳ��f��qZU��u�T�l�Tu"�a�$:{k\��S�`L�Jv��CյT������S��zk�jT�q.��p��!�����Rq�	���$�1F���n��sq��<�L9X�|%;U�,�;a����B=��*%�A��6���O��Q��!/���4}��H���A�ͫ�T~��	_m�о=�f�ygQg*�\*��/��'���<�>�6�O��2E\cU������/��V#���,��!���&����f ��P�j�Z�\�2Ѵ���9�Ζ;>����2�D)udݻ++�PQ�f2���
�u耐�ŻA�l`�:|�L��0��T�ʎ(�B0��T���[ai����SeQ��W��Qr�����~ꃣ��W�s� "D���-Z����5�.*���v
^���k�����ً�g3_�c�ڄ?�#�v�dX�o9{{O�a$�v�K��5�F������O20;�${����{�������F�-�DZbċkm]���E�-9֑��N��fi�*Adt��^oQ���S�Q�+]c����r�J����ĺD]��l9�C�ɻ����;ւٌ�%He��>%���&����M܆���e\����ы8}������.h>.X�s�l��$@%5ư�5��Fv�~���7IM܋�d�!q���ll�'v�XZG��c�1�3�J�����Ow���9?�i؞�~�-������[�?�i�-}�`7��[���vˢ�8��,�!˔I-c��*�p�	J�k����Zr�0����3���~���ryY�8����o�����0#$�@_X�ݿ��P��,��F�D�������`�ݤ��Ş�|x}1di8E��|ߞ������l�MĶa�uǆ%�х�ɠ{զWp%�Pl�r/wOI��b$����ʦ��L���m��|�o-�u|q�[��JÀ+�k�j�.�NU�K���Ź��1#z������cM5�}Z���Pv@P�9�8(4�!��z�n� *� �7��o����v׈� rP�Xׅ��i_ 
��{�n��z�1=h]����>��'�K5I�o=ed�f��&5�]�ڥ�I�jd��ȏb�Y9`�+����Ԡ ����6������D-���xn}�jyɌ��&T�Y��=p㈔�Mr���^�[*�%a:g~B�ț�Jo��Z��<;:`D��V�U{�����J��?�Xg�(�߉ۇ��ql��[��3��}���6�����o'��&.�Q�1{���o�+��L���>U��e�w��AD��z��xÓ�k�� �a�̛�����CP(�0H�S����:��e�
�)���+Z8-����As��S�<J��!G��LB
�4���-iu��Ho�����S]���x�~����X�;ۢ7�jN1��6l�\�Gj�*��Z�j];����������bo�9��{y����M���%)7oKr�B�GBS7�s|�w�X���R)^���UP=v��	�ېp�[V��|E�r��#�ŗ3��6�f`}�4����,X�]�J$f�,�ܜQi��ݸ���d�2�31'ё;��%�t� ��53��!#侤ƩQ����\�J�<�^�hJ%�
�6)&B�H�<0�Sn�ɉf5'����s��}|՟��#��Ĳ/h�����-΢�Н������8�z���?j��p<�I�q
�Q�m�c��ay?1�A�������Z��6��)�kEk�����9��^㉦s���j�ޗb%�b��28��E�3������`B5�{uܮ��!&x�ڍ�CSlm#ԅ�MY_GM�eOs�}J֢TBU�2v�Y����(a�������m����"�1���mM�Y��YbS������*-��������n��]B�5&�v�䬪n[elQN�y�euV����
C�����9eqd�//#�,�h~�,��d��NϫV�����o����q��+h���l�o)������K�4i�9ԝШU�:?)g=:yt:|z ;M'R-?V�����r�1��}�J|����h���G�d��,\EM�������	p"L�m3L��m���\����/����,�����WE5�x�h_����{[�����������y;N'���<���	'�֒>+�h;`�Mw���-����B¤�u��֋(�c��������+�x�F[�PH��Q�gɽ:d$6mpz����u��}I(��+���h|G:<�f@^�y�s��wd�x���,��5�{S�}��P$���_���|M�-��z��p|7>x�k�?*�7s�����[ܰ�z�;���]�3�ߓ9I�:6��0$�/�EO\ގ��2��k�0N��oH'#)9j4	��o�CQ
�A�1�T��Zf�g�ڑ�ӫp1^Bv�F4����{��b���#�)$�T� ��ujU�;�0�M���Y��1AJUu��("��@�'_0�e�z�h%{¶��Hk�TAH�u�V������R�4�.`Wѳ:�7s'K�J�������`O�~�:� W,Ҡ���'��X��z!z�x���f�y'���R�Y�f&������G�ܳl��p`	���	ld{g�Ud �'�`��0��� :e�5��Xn�2��NH0B�~��柆���P���A�AN��:���=�|VSx
��Qg����MW��W�{%���� }$�gRC��7Dy=��x��
`���/fT}�Mc������Ċ�E�v���\ݳ�o�k_P�h���$��p���R�w��U,g�b��8�_@�T Y�I�W��(�A��8�2=�U���A�n�s��D�V]�lK|n!�����)`���rj�Q�H�Mg�E~�<v���1r��5锎ܩ�	CT��ݷ�O��O0!t߽���wp�_z�K恢�/������M��(�bF���7`�.�S��^�刹��;x,��QY�>?K�m�y����Ƹi�_�|�nI��B��*�����#�i���l�5��;�6�z��P3Ъm�w���O �_	_,���-���T,���6L܅�-b����yg��8���Ðb�Xx�����+�B\�f.8�>�^�U�\���*�kk �2�2�!�'fN%�|�]�c��s�O{�&F�Q���`jG���� ��(̍��z����a.�C����r�M�����L��x����ma���eھҷ�=���1)��\g�2�s�m3���/4�5Ǹn�������(�I»��e�u?��bz�v��@�RZ�E���kV��Y��C)a�Zt�5� ����2��/�t�ёj'��T�w�Lv�!ÿ�# 3l5��G,�%��g��F�v¢���*�����+�}�Z�W-3f<5%�&,)�v�0)��5��OD�+/����c�ح�*W���,�h����T���=h�M�ܖ���|�~`	|��GK�d�g�Wr�3�� �&T�YN2��R3��v���Kw��U��:���A�����$Q�}.Fr(}���kR��0�ؑ2w��>�J��ޡ^���4�6s�������P��a�H7�֐��G>�K��a�l�s����۝��%��VWk���l�2�JQx� E��5G\���f��n��}("03�1%�����$&pV.�S|���Gv,-��3��@P�H���Ti9@���Ni���w}=Q}�3�����Fu!|�g�&F�[�C&���v)���!S�q�5�4R�V�t�A�L���0<�:z^��Q�B�|�����O�![�����'|�v��t���X�&H����N��]֍��b9A�{���v�{N+��D���)���MD);,S���A�0T��i&�$3�R�b4�P;��k0b������ѡ�m��gֳ�[-��dﲢ�l��J��0mG��s1B�uG4i��2v�ޝ�'��ɻb("�C��r����=��O֒έ�w�'�d�=siϯ���y�9 ? �lj�K�$������h��׏��� ����hD�ni��g"bQ��1Y��M�h.��Ցp�&I�D�k�!�v� e+��լ���p�HTR��ɒX�"��5�X@X��O�d���%4�-��FwUi�i�M�a@��^��f�����~��/k�l����n���Y��f��l?"r2�B��7�}���r���)O�>��h+����p�����"�|��Rﵩ�67�1Tf�-E;�J���F�ec�W�[b�RZj��!�����_{���p�y�[phnn;��~��Z�/��7��pN�������jq�5�ٴ��t����Y��u����t���׸�s��g�4Gӓ�$��P��|ג�x�D>A�R�~q7e�r|�w���Y���_	���/�E`��7��X�ңV_�([zb��F���i�
;��	m�ƱÄ�-I$�j�L¦��MT��U�r���}u�d]3g#$�P�%��j�.h���s��~�LO��%�3����wM^�v+������hM���ه��
'��$����=�_Si�Y��6(�A�cC´�93[�1$,�%�p/��uӤ�ՐE���ݏ�XuW��z�c��&�oɷS�X��Y�����l�.I�=��<��L����{ۏ2����XA.�������_Ai[VSZ��2`B�dS�	�M�)�@������0�ba^�yb�{2�}
/�,�G�1$���<[��ZC��F�Z�W%BLn��6�����s�<h�./�gnH���-��%�g��LO಩��gs��\��&�[��Ep�+~�"V�Nx��]V
�(O�0���rr������1���YdGa3
�=W$��7�t�;�r�H���2{.B�Vׇ��ip(�}����_sPf��\��h`6�c����*t���"vD����pZʥ<� Gp#�zvkz�
�B#黠v�U?9��h	�x�"��Sg��Dq"�N�^�cr�	z�˘a�4����E�t�+��#n{�q�����S7FG>��殚������1b�Ojۆ635Y�ȼ�e�.�-ug|����,n�ʭ.U����&՛�OI���yOe�za�zzU�5��l
���+���� ��!w�,U��#��%���;R���_�k��� ~�E��<!5�(.�zeRBE��{�*P;����k�N$K8�G�#u����]��R�Q$�V��A؁Ex�ߡ�F��Zy;a*g�D�©�T�H�r��)R&�E��n��|I��&�8����$�+^�l~�yJ�`�*cP/%�,��N�U_!^'ds9I�<1	�� ��a"\���aI��qֻ���&څ'JT3�
��t�@Cˊ��u��OWZ�蜻&��X�Ų� �݁��G�^����J��e㝾{W�DE��X�Mn��*(���_��|oE(Jl�$+���(tDU~�nX=HT̊�/�3M]ܮxu{17@��`�Og�mZ�D�ݙ�fӰ��M�����ek����'(Ƴ�n\��y��`F��OA�aWX�7��2�H������	�D�.D^"$������.���Aӽ·`s�/�5�T�O�"U�n��!�ɲ�`R��qp^���T�vxdU��u|b-��)���h�v��l�Iӂּ�����v� 6�vڊ�`��/t�ΩU��'�󫆴#�h��y`BO<�<V��b;px�D��K�P�٦�{�_ c4?��ܠ�
YZ�����Ԅ��2���bW�赥�vb����J��!8ъZhb%M�o��jpA��}[ݚ-]�?%�*}�2��|�����n	/j�^����SL��#�;yr�Ե�-90��V���k�c�ѝ� *�-E2��n-||�D�-�A�F˫�����=_b��h��׏"';>L��,���;E؂��xHD{��e
O)g%�����x��=��E�����(0�X~u��?�N�R�0�d�8)Y�����"P��t��gV�s��Z����i��勜��V�r˥�u��,7���`q�T�
��Ϩ)�p���Yh ����FpW��}��;�o�����}�J��ǖ4��H��o�X	'chv ��Z�AO~�Z#�*
��Ç�)"�s��!E�N��iֹ��O��[+x?oLp�(V&��h��F9��A�L�N�O�"�jƐ��oi�}�P�Fum��$��^�9LZ"���n.�NL��ͫ���c�p)�W�����b>޶�?�>��_�)�w���m&q��n;؄��2fQp:g��b�V�A���ԱRk�����C
�RUh�%�S��ߝ0��0id]�d����N�:�ߡ��\��]f�Yї���ˏ���#{z�[�sع6$�ׄ�C��=X�Za��X�j����V2���M��ٚ'8���� �J����2&YY��+`���w��h��.Q���U�L��ڦ��I�5�CӇi @<����Ƨ�CW3����#����4 Q�]z�L5æm�7a�]���ߜ�nނ�����ܧ��e�tbF4%��1S��ͬ�:bB�O���)4f�|�v�Z� P�P�׽Ŋ����2�9���p��JN�OD�M��%\��*X��	,:�Z�~�Iy���
���0�>f���aw(	��)�㧦�  W5�遯�o1�<��}-a���}��t�� [\��
��^�����h�,�k$�:C���Û����Ŭ1�����k�+bOF���@�`��'VB�w�>�N�4�~�dNC[�����rb�M�����4	����W��gm2'�*����Gv"���~ac�WG��y��8LE��x8G��A�Ef����#�,�h�82xE_��|=�Ʋ����Z$�.�HP)��aw������D��"G2,X|�9]��Wn}E)�u<�L��˶��4�1�]�=�����6$�$(��+f����W�O'��=�UM��m�4���9�h/���yN
��W�E8ۣ�h�N�t�����F��E)�B1���b��V\qM�N����VV�#c�y�rс��}q	��іZmL&{�mf�_��xֽK�����#�Mc)��骿�#tj���H�-��A&�	�l�84�����jt���j�+x�/�Y���ȕY�t��5g!�!�!�k+֮찈��c�P۴�At�~A;�2�1_1�R�\��$��-�r�(B���8q�t�o���=�i#�{���0������p?�pv�����Y>y�K7
qy:�VA���C3��<ӗi�ƶ ��ñp@� ˂w߷P�r�eS�4c�E(L�,��	��Q/��4a�&�͊����ya e��SJ7��q�j�D���F�鯩�]��do�K*�<v���q��[7��t�j�*��(�3�[|���ٜX��h����3+B-�*g2����+!-�hR���џ8�[���e�{�O,���E�D�������k�п{-A> n�|�S*�؀R��L�'��S�}$՟Rn�����>D�;�?��J3��d�%��Fg.��&������Oxu�*mM�`h2P�1C���*´k�TZQq]����������㒹��Ȩ*k�3"e�ܙ>ڨx�VH$�09�$\���`W� 6,Hڢ;���������>a��FQѴ_G�|{�	֫a:��_�RPV{./`�w=�"��P!r��Ҟѐa:-a�k�*�GV�gjؔX��9K��q�9S��=��Qй�w��N���?6�W�
�zZ��;qLlPVrf��>A�πL~H�6Uxa��l9�i|?[�Q~����xUHH�ěA��\Zד	����g.���� i�d*�;>\+������I�'����nX��U���q�Az�"D�b�����Tg��`��<�,�u){��k6
�]��j��v5�8�.��^[D����Џ#�8YAg�4Q�"�e�.����TK'�=��E����D{���}�sk�S�N� �'I�U�J�;ܿ\����Q7Z^M���aS���k��73����b�T���,|�tG��4��X���e>T,*`Ȁ��>��KLt��ݿk	��*���nI��7u��>���S�#v�Pm \������]�_��8ZB!���tD��9<#J�r��h|ʿ����W׸���ʻ�~r��� ֑�?N�����Q{S�(�״�B?���ve�{>5F��㯧�F��>�˪uvb�'���_+��SA���Dy�����eK��$��Aé���x��7C��[��e�F��j��숷��@ʕ���m�$�PQ���J1�q��\�d}���%�S%d9����V��gF(����d�7���B~�{�Lw�@�H+�uD+NQ>��9��-�X#���lE����z�U���379�Ȭ?9/)7.�DӒЀ��^�J����ߤ��pd�i��NHS����nJk��5����4,���8��eAno=����ww&}�ۅ���r��:R�xk�Y��]s�eP��gf��Y�v�	#a-H7�2-����|�J}���y1���m�L%C�u��,'><���6G9W����G$���ATGzV�P�T��Y_'�	'���F���L����r�VuW���.�o	_p��NhW 1�DE�˄4g�y�я�1dyܕO��bS�� �o�HXg��ٺ��v��W
�q�ǜ:��ibO���"�!t�ȺH���7Zͅ[1ɐ�%�C,q����,Y++yya/�xjz�{�X�:��>��Ӽ�&3'��[Q5�K��^?v9�Q�����W��D�,V��th6��XE��GCN�}`їdPЙW~$VuX	OIx統k3^���_*�(9��6(��
��/_B��4:R���"C$Q����t_��Ҙ�ʼԁ��TSW|1��`�3�r�������`��A�p����6�Q�*p�L��7���������L�{����� xjaV��黔C���W����]�~3}ʩ�P��	�r �p��ߺ~�c�����_RlM)���ڏ�Ƀ%ҟ���3�t��?�/��+'��}n�5#Q�E�m>�>,{t
���Ef]�Dz�Y��8�m���"�`5ů�XM���	�yQ��Kg���| s��G�s��[�D���š��{�`�C���g�E#`�N�����`�������̥���M2D3�n��6��\Z�,��,ݝ�U��+Mke>�O�����d�J���w*sW�ჱ�̮O�`��׵��}��Q8�#�ۓ��Lb�P�,_/>΄[P��=�(�V��J{:L��W���d�-n���z^R$E/�&s�F�8ޤޟ��`��}Ɯ[��{�C�,\g�p��\���i�S~�B�-Emvbܹ��j��_��^�<��M'�5��N�4sj �2����tNO�ƸN`�<m�K=L� �zԳ60�}���\*IX\"�BC�CL`5D�02VZ��<,P N�wUB��L:��E�߸A��,E{G��T6"T@w�4�$�^w_�� �9�˚»��g�b�0���o�ڋ��{b7yk��0Q!��&������)�z�G���M��F�0�H��Uׂ�ICX�[�G��u�#�њ' [�t���\��XqNI�Ee���o���Cl��1ڞEf�M2/��~�mt�hIqD��� U�T�H�n"�]U����ԓ���`h<�Z��w+S�M굗=0c6E�#�9í��� ^�1;�9v��dm�$-�E;ި�	��O��P"��F�Z�wM'3f��x	�Rv�,]� }��q1������|;��%��N�6�����ep:A��fY�\�py��d��$lb���]��塛r5� Q��P��_���� `w�5" cD��9�Q5Xj+�a�)��d�Y7��׷ߵl���L(�Sp��K�ދ����/e�#	�	ʕ����������H�ת��4)H��<z�n�=�u� ���H�V���S�|����e�Y8J�^������_�t6���3e>ԍ�jC)-_+X;Q*N��:o6#�l�2W�-?P��Z�IV������7�um>��KuJr�XH.R?v�-���/�{沈eq�剖��%���=�Ţ�������[������p��G��9/�5�r�*�ˀ�N��R�e1l�1j+��kC��l�팽��᱀����~�Lg>1� �VXbBXs:��
��lٞ�(X<�&��J�rd!`v��������� �b�c9*���;�C
R��)�c��T���ě��n�2����t�E����7 T�G��G��=*'��v�IdS=���U�\�g���.��I��	�Ih��`���%������g���M���,T��z�э��� ��+��w��4����IW�����j�n�Z�XU%y��P��m��՟_���|��b� ���HI����:h�Ʋm��p��h[F��[�u����PX�Ժ�_+ʴp��¸��eF���-���0����6^nf�zX�1�a����8{�e�i$;r����|�?_n���[8�l?���A�FS�OZ�Z�&�Wq!zh;��"�P3VYq�)�$��]ʢ���"�W��\|c�����V1�.�Rs�V��Jn�!+q�H��
�by���Ym����?�J����J�;U�ڴ̀��~^Sd�8K}��,R�*�k"`��re`-�("�9J���=�1��9��M�UWX�'��h�a����e��鬶o�N�᧐<�KpƨQ�6j(.�֜kR���@i�$֓�����#�1R���ߊ� �Q�2#|��A���?h�|� P�������=�,_���X��qV�?s矯�th��+�>pt|��כ��Xjz�B"f��[cV�Ы�h�yA���W*,��v��_ӎꝦ�r��Z27��������L}����V�"����a��õM��dT����g�(rZw0����뎾�ԍ��\�D<���.�%S�s���8фt�ӿ
�R�_��ҧ�զ������אy���˯�T��5�g�	�07�?MA�f=X�t�c����X�8��>Jx,��c�>kY��=�"����Z�N�� ��ܱ��$����N��D:"��Z��Da���3�YI˔o�<��}�2r*t�Gdp�ym�)L·���sO�7d9p\�uE�� ��m4�І�Z�>�K�<Ta�kb&.�4���H�T`%	:���T �7�1��$V��?�G1 ��bW��̦v��tTR��Ҹf!0��G�P�4���DU�@yG4��>3q}���c�jFy���� �)u0�-rV�^򼃆}��B���v(�����S���~�Gʀ%�e��C���q@R��i����9��?�N2���f܃���'a�~�"f�4<oЈ�,S[�����-w�����W�u��N^�!��	!�r�9��{��F��vӍ~,���ީo���@�r���#J��b�Ǘ�-���L�=�dx��LVk5��O6;n�#N'Rz��Q���H���s�l����>p)���J�V���b;�e{�1���8eaKd�J��7�g�
�TP�S� N<p�8|$atN���
U�T���Y����(��Z�P�_��zyT|p��ë��唜�c�d�����?%�FI���ӡ����ҋv�b���'���z��@w���F7��*_�h������޴<:���
ZB.��dZ��$|%$��B��cd1�"oh�
+ߢ7�|*_/��.p(�(��'Ӄ�h9�d��`��qK���s��H��_S����� ��e��-�ݵ��Z$Į�ѿ���]�@_KR4�W���i��w��?/L�� C��c;p
�j��^��ԒaF�6Q�?H��;5�Ҧ{	��u���hb4�A�4�ˢ)�����'Y��U�`�5��?㶏�Q�%��2:ýj�f)Z~�<�c�y�j �p^�&޻�q����#ȳ�R��iב+�r�u*+d#bS�0jWRm�^r-�"d��\,���Lhq����B��t��y��*GZ[�}����/�?ʧn	L����K�F�c	,��A�;���q�n�3��GNʹxG�8r��ܟ[��7@�{%��^`iwݔIxZn�3#C��n7�h�0.N���!��#�LGW�,3�%�i|����w��Q?��L}�P�kA�'�m�Ǳ �&U$�u���)z�����H
��g�o��a���e!~���bF�H3u���A�Z�����i"������/�r�t�n��m��r���G�����TcH�k�����h|Kt�Z��a:�{�QV}�~dNQ�0�����H�D�l�X��b���}����$����lE2�%�H���ˎ���Q¤��KC�U0?%�R�^��
�N���b�ƾ�������B���/&��|�)񞃅qr�3���{��DO�}����o�FH��,�z��]�ǂ�a��Y�e&�+�e_�h.+`rmw:������k\cs�;��[rB��޹f�x��P�藗Zp�,�|���4�S�;	��-�2�����êʋM+!:��e�2煰%tl
l�eE��㤝lr-��l��ϓ:7"�:�~*�i��7�r��R+Rډ��[/�-KQʍ���i���|�ŏ�6ɸ����	��Wb%�~;���� ��v�1�"O+��iӓl�,{��)f�{(mvh|}]K_��)x���6��\{�lB����^�MG�-���E��.��n���Ϝd� ���9�.?#�D.q�ߍ�'�e��Av5Z�b�V	�*KB�9�Q� ���Ea��hx��l'�Ę��Z���As��#]c��m�R��Kѱ`d���&���YQ�+5Spb�Ac��o<���Hu:�WG6�S��5�O�����l�_}io�4Ư���������畊����N�
f�B��Śq'���Gs{�Z����0��W�R׶D�BD2% �MOsF/��6-V<s,��;:���������"�0����������c�SQ��@��3KHk��O��S��V��;[��-ʭ�k֑t:����LK�6b���Y�xfp��6/\��{��F�=r6T�=v1ǟE&5�an`���ݪ�5:���x%�8A��:7Ó+'���<:����-�$~t�����R����~'56���'?3��^��@셗R�x���]y��})&��ԓ��&�$}:'}��T��j���i��;��[��&��H�p��tgw�-�����ϑ.X�u���0���w��U�����ݺ�m�5Qw��|5� c�kJz�ˮ
��k���|ZGw�6h����N�#@�V�W��������)@��A���;�/��5�<�a��o"e�E;�n�o������w�NJl��?%�	���a�C�Q�5���5%���աH�	�;o?��]�� ,�kXł޲�ź�4�T�����<�4O�pV=_�&+�i_h����GΒ�&J!���Id*<' ��2���Q�^m؞�9:�4��1N�Y�e�:�t{t17�� t��L�����V���W=
#Q]��J$���=�0�X ]��1dugٖ�f9��[�7������������I!�H�&Cc�(�������z���e���d�D{V��^��r,�7�����	d��ڭ��U�%����M ڕ������f�"of�D��޻Z�c�6ҁ���RrF�R+���9"K��(��ft�'�I�5ͽ�d^��<o�G$�:��p��6�����OPV�Z��a+V�g���p�ư��,�/ټ�M�a���\�F�0��J�0^(xP0`������v��VՃ���O׾�lfWĻ�����"�<7M�Ã#td{��;�ω]kv޼�����G�_�@O����6ҩ��Ι�@e�렂���/�.�5���	����=ɐH�qR�%�p��ی���b�!6b�&ڼ�wJ�Yǯ�����or�;�0�� ̡|Pj<,�q��̶N�@UPH�*�|0�XG1N��u~C�x*�R���2ؿe�����I�Qe�#�ww����uq^׳���7�>H�$�Ē�d�іi2@���d2g;hd-�b�6�HCG��K@�I��qqo����J�|&�o��`�j$�f�V<e��9��7O��ܕ�>��{*?&�"�;��v�&���;H�Wi��%���+��15�踽]34`�~��N}����)��{OX���\�W	I+���:���m�tH:r���=��$�Zˏ�����t3��m�R����{������4�;�&�d�B0�,��� �����\��0�g.��9� F,�Oe�]�^�IGɛL���8L�ر�[Be���+�ԩ�m8�~I��\�� LIvj#2A]ۖ����D܀��@�E�J8���ޕ�[jυ�l�[��4w;��3��p:����J��h�V�ߙ� ����⸆�*�6e
��%�2�ɀ�5�'����^c�|Lq�2�lj}��"'���w��ϼ�mW��Yky	��ޟA����,��xP�\���0�U�N��2���s>+r%�=���
}�����`
��ɩ�#�|�	��z����d<j�i�W3�rk-%�f�	I�~�n�[��O-x7T��pk~��o.��n�D�_�m�K��C�i<.��	6���7ozb���Y��r����Å���AR�)|^�g��؛鹛��Hg1��M.����h�㼬@��iP�KԐ�J||;��_.����me�.B�f��c~CjU𚲽�̄9$��a��\�9J�6w�5�{��̈́����l�+�i Nz�>F�U[�i�;�����f5g(�W�N����].�>O�C$��*6�l���e:�ԅ:8��F���@��7��>�ns�`|��0O��
l�>��,�����oZ4�u<NJ�[L�ӳǘba%`��D���C���	SI��Y�(m��;�z��2�yǟs*9>����`�^�YUW1�Ѧ%v}ђIrh(OѴe��\t-��
�ES�w��3�G��و����gT�����4͈��s�k�vHo��jth�F��{	1M ��N�澖�t�Ś:�,���3$d��:���Fe/0���LY>l�����jڂ���YB�z�̺���ڙ@���l4	K!��x��ه%�#�0@� jqL+�{��Śk��^L��,-9_��SD[<�Vl�]�v�w@���5e���l��������{v��z:Z��!,�2t���Q��ͣ&M��C�@��:�eډ��n�� ��u�Vz),$2�zgϪ��é�LYˮ�#��B���
s��-t�uf��0�� �����������s�������C}����J)z`(�"E|'�����h�ԇ�0@���c��齾�z�K8�q%�E��3N�D��xA�}w�^3�����E�G�X�=]�)������Gïw)I�$������HBL���뺒�J�|�]���:�Ľ����l)��r'c����兌�(��tF4l�j�[���=Q�ч-ٔz<;��O��F�^K�M���������|z�g�X;��R�E����k.)^PG��*&Q��ݱ��Y[f&��D��9 )Hm�7�IXt1��@#px�m����[��>�ٙprI��B�=�	�&�'�jIH�{�� F�5U��y�TPۄ�B���e�[�P \~��4��Y��N���2�ah=l��L�]�U�����/�4y��XB��h>.���kq��[ܗ�hB�w���>����\��΁��qb&ڛi~R��e�����Ȁ�<E!�_��2��V��n4�*�̡��Z0�wz���an�l��!o���eĦ����c3+�4˙�;�Bf�F���oS��SrKpwͬ�B�B�.�[�!�Pg=�[��6�
���?)5R�M���𸉍qHѦ��in��k�cn$.[�v2l��4q���w8��f�U��.@��"rj�.��G�A�����j�3�lX�S�"ϰZ�L`��+G��t�o|�'�4�יϺ�Ϥ3�P�G�R�̀�QBN��;+s�S{V��9��֭7���ڜvz�Om�=VF�:h�;v(���N�Zm��<���"@�)���؍��Ԕ�ԝ�m��0�|��2��|�\4��6���E+Ժ�,S{�\f��p�
��sk�J����ʾ�Ϲ#<|$�Do&���'�dn����5���E@YaR2/�}\/�9R��l2mA�w����sE��Q_��wN'�:)
�������P��k��Ì%���""�C�V�f��3�qb�i���M�W�|5��8���8�v�0S��c'T8+e ��.�A�\��	5���6c��]���AN�?��ߩ�f�Q(u�U:�)h�T(�}���th��V�$�<��
	}�&Y�����ǥ��T/�[��"e�7*�a��@�aD�o!�i,�b���%X�Bs�C'U�
ßg���ͨmw�af"�j(V�Ga!�h<�}o�S44GOE�3�P�jA̙kj��~M���w�����{"���a�D�w�AdqQ����� ��kR�Կk3�h!q'�)ė|�K��dv�Z�< �^z��1��&ͣ���?�)�FU�,t�[9���cCċ��I�x*�V��%H)vʘ�!��F�����і hLVʀ���鄝.�^��` +�&ep���Rb�t�A?��%2Ť��8	D����_7k=�w�z��䵺�]wD�[���g4xdUgg-��M�k��.g
������Ap�Wx}+��;���c~a�&,1� a!�����u�HE�m-)����4KP=s�%Ǆr�/�B;Ɖ5S�p�d�)�Ֆ����[�BYC7 G.�p��\�o�un�'>����W�����Ҷ^o#���N��~dK����Dc!�!ћ�s�R�j9�{��ή��<�[�=MR�W�~���('B����/�Q�f�Ͼ�)g\�쑾K�3	7~\��C���"��!�!�}�.��=O�$�#�.<��L?ӵ�L��ԙo�=.��b��V=ƿ;����/*��b�V�E�������u/ѣ�Ϲ�ԝC<�J�/�i�WBvڏ#f˪\L3r�a��k��l�Zpt!7��U2qYTq0�CU�P._A �о_�^������8��b͟��sM ���'JM.�N�R�g�7�|�b������|�	������^�n�}�F
�N|G=mY~o��Ȁ�Wp��;�������J7�Yw�pk����6-� &��]��'j5y��M�>9���<��=U�ȋ��Dz �O;���b!�q#�ݎW@UU��D��ǃ��44,��*�����|�-�ٓ�>h�����.�Kg
��.���d~> �w�_�P�g@v�Ss`�B��U�@̏������R������Mq��WHDp��n֨�?%Jǈ[��0ge��#�*��"�WI����xf>�nǒ����� ��f�Ȱ�ﴶ�	�>{N��n��72g{�\V�?k� ,���PL,��z���%	X��|mS���������8t��>#rCۺ��-G�{XtNZJ�����T�fj�<
-�^ⓌYG��4�M��Ŋ�\�RR��W�����'x�&в����[7�u�B�zY�"��Cqw�2s�IMn_�龇�HX�-7���|&��3�x��i����JN<|Gnk�{&N�� T>d�!�=�TpAi��utͧl���^��ŠSw� iZ�ͬ 3!��?������Q�#Z����A>7�����Z� �=)]2��̡���
?"�����{�ۜ�o��+����*װL���)=<J�/�oJVQ8%1�@���ׁAM4:'4�^�ėЫ#�{BӲ�:�k�V"`��G}JR�= �k��DzQ��QG8s�����b���!�Q�?�����1O� �Z96Y��?S� ����oP�������R�����^���:p�$Yὠ�Lr���e�h�l�%���t"���h�dS�r5C��r�b�܄(�B���,YHq+2���cc�SQi��~�~�Qyv}�!�@�𣈭�8AϾ}�bk����v*��S�|�UB�N/C[2�m���p�&�Ƣe��RL�#dSx�럞�Տ}޸ia��'����;`�NBz�k��!�\�~�,�DZ�*=���#,��Lc>���|��)�uY���77��+}�����B�uH�m��1�Y	u����j0Yw�Nc(;��	�|g���uy8&ʲ����+��8��)6����]D.{�q�YL�CEHA�j�k��=a�殱�A�ϻBT�0/L'ih\k��q,[�Wjq��}S��<�>������d�����ٳ-Vp�7�ߝ���*�(��~ �3F�^� ��i�i��F�daO�,�6���`���ja��KlP�ΐ�ˠWb���Y��ё�U�Ȏ'��Q&.�"�|���.Q�53�lG�W���-����Gu�1� &�\�=;�HG�B�+F���gO'��,�JTVRZ&�և�)m��Ao��u�����ۅ���,�3׊����3�w���5�Q�eZ�������VXl=�$�����ts49�lk��̓ҕK��|���T�K\s�����e�X����!'�F�"@�9tG��E<�E�2���&[��ovR�u�a�-��o8���sU'���e���$����޿�IE���s��4��H4��X�E���3u��>����D@tϳ�\43頂"z�1�r0��K���v�v)Q����-���Jp����h���RU�Y�t� ;7��g���j��uTO7�~L$�^��3�� -��am�=��7j��+�}�ː����'sR݇��eD%����jv|���&ٙ���%
r]�RK���ݲ����o��R��m�?*�RJ�Bf��G��[��6���=!.&��E�4�-��΁0_�R�C��9��x�.�7� ��E�5	P����Gy������,�!ɻ�qNg5��{��u���G �<-6�]G�2e���Z�*$��G� ���7�m4Sv'V�7y�@�OF��O�Z���°>U&��K~��a��"���(iϥO7ND'R�Fwi��5Lv���|�@�g�;a+@N���aDSx�������4�v��W��Ps��u����x�&f���l����{�z���?[^���0D�5�S���;|��86\�"ś��<?W���2ğ��б:xg����\˪U�d�u���D�z��m�sӔl�U�8m�v6f���g?���ɾ�wj��a�2�@�&K4UT�?A�?vÔ��'�as}%f��>XE;P[�c� �?]|B��g�h�=v��f��=��K��bk��uq��_#�)AC���oR	�v���#��dH�侖c�z�l
�j�r��?��d���r�$k>��Mǜ\�G��g/܊}a����H4����È�O��sԾ��Z1�hU�dQa��1b��7��$:#�o&��aR�������ਫ5V��}6�]�J�B>��u�XL��t�=�2	�OјX.��L�n�]i�qPN�&`�҂�����a�Q���dJk�FY�x��4�݃>%6�9D,v�+z�8Ы��[���6p=���d�7��zkj�ͦ��%���H@�Y����j��p�\�S��֡����)N�l!Ir��u�o6z�P+D(����W嬂�Tr��<D�������/J/&N�|L�pkT`>D>2��q�孢m)�lJ�� R�Ư�D�&��yK���}��>I'B����Ƅ`|n�/_�B
[fBz�VHR�b��%���dM�S�Ru�װژ]Ia;Y��s�JwЋ&:NC'���$@�0��8Ț9��|��V�թO��u����ƳI�8���kD��)�����^�)r�N����ȣ��#�|�����Y5LO?�dI&�� m��z��q��4'6灑���}�78�\U\V�T�<��P��K�G+�xSZF�Wl�)e��RU�MHҏ���9V��a����#Dy~ϬxG����Ynr�m�/\���S<9M��r�Fwy��yC��!˕�F3�������h��{�Nˢ���0�z�U^�"�6��e��Y4�2��'B樞X�)�"%{w �[-W(�S�$�H�Tg�@>�4��݇�I�H)O-�OZ��W|D]�8����N���!ն�ǋ2�()�a�Ѿ""B��w�"��04#8-���D~y������
�a�L~%�=��9����TG���$��8su8��\Fq���p�m9P��YH��˵8�Evg�Ic!�b\�S���Db'cb#��.w�O�J�'�D�p�;.�k�^.�@7�j����Zg�L�{�B0,���f�J����G�HYM�|�/��,��nx�P*����͒gO�����^7&o� ��/9����+�l���	����pb����T-���k�2#m����G���/�7�NrL�_����_���^,N�U݈;L� `���ȐB��KQo"���%E������I�-l�4n�&�&
���m-��XC]�2rS0D���1�5;�Z�	@~IWI��ý�S��eR���qmL1�ǌT����øoaM�w���t'���<U�@�S����#g��dz.���(7%���κ��엖�:�?�\���c�N�w�#՛#	�:&S$\��+$I9�7�L<T��I$=�2��d#O�~�S�;�����㨑@���V�X&z��v\�o7���%�ӌ6�rh'1\sۅq�F(05I?�	D�`{�i��e�b||uLF 	Ù|b�ؤEȣ��3���Д�G���+���v�0A��A��i `�����C�l>�g�ġX�ub�����ga_���
9��'Tv��5�.�CɣT�þ�{���na�V�y��ȉC��F>O�6P`p�T�x}.`7Y$�����n&�N��a���p��+���K-��ٌ��)&C�Rbq�_R�����L��zf]��� �m]��^�5gd`��PI�%��s��]|3[�<��uVN,��7�0'Q>�RX�qd���|��ٟ#��#ad���K�M������}��������S����O����S&���)� ���i�:Q�>�����U5j���s+N����3@#��	�!$�Y�m�������@���T��w��~�k�m(L;w�k�b�U��g���CQ��\�q��g��a;vF3�4.��A�[#��)йLbݭ��s;�a��+�A;��eQ�PL=�wo'l�狆�����ԗ�,�hW~"k�R���Ċ��?gpƥQl	c��J�v�F�_�J���v>�$����V*ӷ{�1���$��Y�ȡ斠�:hJ��z~���`��G������b��k�M,��(:E
;�8j{����kE���J%�x����դ�`u[��2oH���-I;���vkUó�����@\)��~���P����� ��,�q`|�gұ�D�z:��:���,�@��O�PZ�N�Vak=�%M���W>�fؙc��M����m&w����Hp"�����p�S����a�j��%��U4���x�X�7���3�{�gr���s=�Ĺ�q��^��0�a��]�~�%��NѤ}sg�$�
�b�L_�-��9���r��<���0�7lY�?a�4�d����Y�hVH��:ε:�C�#�CB�2� ���a�nk����U��wш��M�'�.�Rۥ'!>��F��#��e\�+����S�%c�r���T���2�����`v�f�/R��(Yͩ)t���>�m/6����rP��%�낐WJl&Wٮ�U���~�K{���S0��(O1H�B�EK9��7N�F��E*�1�IM���g?>��U�cziuQpc�D��u5�e�X�� ��Sǫ\>��` ���\5�ihg�+�-4��2��{-��x��'J �ei��Qv��#�#��c
3#S��Nm�ni�xظ{;�ϸ$�Tu���R7�}�(FP�e�̅�Gu`�9��$���S�Jk�v�428M��MŶVny �iM
5���@������Ԇ�?���i�s�K
���h�,��KvV�L�9U�'��ɗV�	� BN�:����"4�����{,��֭N����=�8ǜ�o����1wu�'m0o�VW���s������Mɽ��f���m�e�b�|u�X�}��/�	�)h��ڿ6�{�9+��$
���̲�Y�������Q橎�'�FJ�Xz$���Գq��)�I�R�������!�\�VS�����׌4��A*θ h�
��:��vO�)�W�qgnL�1G�\b$�
���:���HI�du�=�v���G`͟F֔�+�sw�O�@�_EXw`�l�yژ�Y\�ae���Rj����O	5��u'�{�,{uj�����)�f��\ '��v�ZQ��H�H�g��ܧ�h9�<ӌ�d�?еf�A+�
g=ě�E%�赶��*��Y�Q:q a:� ������3=
&1���f�VP�%����Dl�D�n؆`󢯹Tsc��ɉ\���^�y(�7�U͈��/��u����@:Kƿ�"�`�DP\�������1�	 � 1뭭�[���'�߻�p����xD���[��d3�e�sW��:���?��К���
���>�����Z\as8C/S�)'�6��b�l4�E��'��{Iմ�Md^!ra�p�MXkT�1���.[�a�{(z�J����B�mOȠD�IÐpV���������΍Ȃa?�e��>���'r��E�q���6-=�+Ԫ�Y���"@�v�y�|��z�n4PI՗{>t���f�8���YŚ�
���u`�n�d���W�x��$�ASbv��NY���e˱�{�c �����W�AĘ�ɭ�ٟ��q2څ;A����t�����s���>T?re���Io!�+��QƸ�jk*��n�#!S�Pݓ����}[6��7n�]ȉ?��G�ؘt�b��!4��,�Icw��;E%�����D����*��'t���	�di߱�g�$2�;����-����:��h�хCm�9c���Ć���f�c�����F��-O09�:�X���tw �Ğ������N��fڷ�PA��:%YHX�"E����p�U�=���҃�$��
���/[�'��i]��c#���K��L>@,�G�!'g0�n&z��w�3�	��	Pz�Ye����h�0��B�>�� ��>�r��=i�b�?(���[�en����tFqנ*������N�cW�G���h��Y���;m�s��`���1���T��z���^8��,opI9~��y�!]<�Ζ�F�^�7s�Fc� �+�V�&�������r����f�y3h�i�9_&���t-����4�/�5`�w����[{�DƼڹ58|CXʹ(��-�W�����OƜ�5��`�n��MT�O�2O��o��̬≝���!;9ҋ��������@��%���� WG�Jv�t�����������ϝ�_��'$�M>8X�H�])����OckCV٦Qw@e���K���&6�*w��)|%#�}�W��=<&Tk�U���=��G#�2zw	����U�C���i�Ҕ�N�[�~ c�W���A:��q�K,ܤtN|Ai�w�~:�r�B���7��ܼ�� �_���#�(��x{�J�l��3�=�`+��,8��j*B}��8J
Vz�����(�?ٮ�G"dd\s�7櫕j�z�w0��z���o�E	�d:�` *�w|P#&�����Y`�	�-�^�j]��R����p*I��(y0J�j�J�Sm�"W?(R�ƽ�5�{� c.�)�)�������k3��&TgL��6�!jL.���,�b�"$j�͟=
�=����t� �5y�+@G��@j����SC�7��'0��t�0Wa�g���Z�M�����[h���\�!ǡ���i3q��F��Qx�1�c�\��>�<��W
���z*Z<�e�^Q�<�V��O�ҙ#��ܱ��V��14#��(�o|��6^�*��y�X���U��?�+�og�����<�{�p*J��c����>�3� ��.�E��i�1ms�ST��<ל'��*��Z��'?����IB�,Ne���ͫaP��e���S:s���O�W��ί��cu�Jz4�`�ŵ�w�F/�GN�K������ضj_���������;8+?���������6$����f�D��U8��na�T����fM͔_�׏Ft�tQ{�)-�G���2z�����ю�Z�K����I}wo��3��	w�XC�ԣP�C���E 8.}�`�6�⣤4qH��O^)䃠N�7���!���'w�`l�-7�����N�Y�j�'�Ҡ��[�n)���������o�Ϸ�}Rꞻ}t#�qC$=k����	*��]!��}��������E��������
p�Qo D{0층g4��˛}�c�����j��t�4�Ur߼ 2�E��U��eX��0�B�4�Ho��b�h��n��j <�s�׍��*�����o�l��P�;�����[jE"�[��ѥ$�ڲ�1�$��>��B��a��4��K��8bB��ӱ-�Za�ӵ�-��]�8+��߷�z0PW3�f�0�@�V�V�lbH�+s��V.�� I���>;�j��Wq�w�x�RWJ�ʹ��8�[�Ƞ�	�f�Ww��/"�����H51�i���n�5.�D=��� _ښ˴���$fQ^p�^�4������Po��t��1�� 7a��k44��W ���^G�x_��,�%����Aסg���A��	#!�M���TAra����ttt�k���,��0\�c����Ja�0�8t�8��i�Fe[��hshAL�d�)�Gb�5&%d{��y˳1V���vђe�8K��'o�e�億lH�q�a�*�2��M��ϳ��
��E�	j�ѱ�P4�\^��{Ap�N�t�η��0(R�S����U�h�^�n��N"5^�ӦR[9�dY>S��l����GF�.�F���w��/��HY�!H4��0��y҉����u����N�]G{z˯���:��Hn]��݁������h�`(z�m\ኒ��$�<�m���J�W'�Y��ܶ�	/��;V�A�)��h7ߵ�|����� ��~�%]i\�P_�����͸�CA8&��(�R�Z�q�D��u!�.�!"�����f��$��*&��q�
���6�|��5R/�C�z�%2w����1���M0+S���O����� ��I�d�� d�Iu=���%|fhqг��uj5�Nc���o�.K����Hr�Ǖ��VYC@:N���=�ݛ�.D�t���-�.NN�?�,j֑���;�մ�7����o3M�ם	����@�mkZ`�͕�>������m:iDG�p����}֭~NL�������T������.3V4�@(s��苜W���o��׈�f�������t踲��F֧�r/_�(��x�[�"�1����s�<Ҁ��cs��d�L��J�(4,��s4;�$�����,R!�AE{�E2��9�[_�&Vq'�a�h��>��;�����s_����Ů�6�D8�n�K2S�\���͖g�*P�����CBC|*vg�OoV����1�t��[>��	b����AV� �5^ǔG*OY�8�������D��_h�.�_(7$��Ӎ{�Ȕ�E�rh�/�!�z���t�s�!����(o2��B�1��l,r��<1��]4+|�L�����G������8^8;�*#�o*���i��"'�&��}�I�4�2׷.7�ұ����Ko���5��[U��ٟ�i�o����x�
s�S�t�-��U �ݭ:��'�F6�f���c��ހI��Uu��{��:�G�
/˶���ޙo�54��b-���x��:C;��<��P�{�˜�,�P���M� �)I%���NB�"v| ą�F��׵�ga�(�+�I���_O�wZ�+L:8l�����8]i1���i!	�Q�o �aPxf�ȩE�
@����u����ʩ6����{jP��R��uK�Z{�y@����|����{�ԇ<�	�Z��h�yY�Sp�ȉ�s(L /_���`A��?g����s�yH�If�|F>�j�~��gaW]t�4�Nz�23�j���]�]�(�-X�:�����x��]�z��2�]wq�93J �]T01��T�r�d.T���L��Z���/ξ0�������0Y��h�A��ȒX���(��>��O�^L7׻�
pN@.+7G%W�y��S\�x�6 !.�́ է�5T��Қ�G�ɐ�Q�&��
�`�m��Kh�r}���%j6��MX^2��	z1�-ʽ�~)�K�Ȗ��ȉ�b�qٔ������-N�_��u�ֹ��^���'��5ic��4�R�z� ����P� '��V�e~9|(�,����T���B�6�/�2K��G� BШt����Fcx�*�4�7��I�����`>C�A�r����_�ɐ8���`�ꊦׄ}s?C��|5��d�^�v�n,bҎ���Ԑ�^�	���]NX8���ف�#e	�|'��h��y��=O:K����G_�a�j��@\�R�ԼF�)��˛�r9y+�%Y���[s)�䡸l	�����`����U�Ǩ�Hw-Z�|�w~!{����ț���O+vl1^p�b� w��-[u!�B.~��\'�9��\�Ø޻�j������#v���	�J�j~2D�&��@���z�5Һ�i �6�m5��M[7�x/�ְ�%��Ԡ�F�>-��z�k�e��z��Yf�0��?ȁ]Nr����y�-�fIR�e��B�ے&)���P�����I��H%
i51��.ҳR|� Ah�0�Ό�~�Z�#�Au ��	�J��i��is������Ż#�EI�c��&ǆ?x��&��Q��˕=S��m��(��[���{� U�C{���X4_ ��=F�Y�_���+�21��~4v}�UN��Ӭ�˄6�����Ckj�����U �5�������"ќYA�bRRP�l���c#��9AL4@��ڵ��S����*�;��4 �~�8�%-���_�G�֫ ���U�62?��HJ3��-䘦ɽ�WA���36р�q����X�;U��e����Sz-drF�Tb��!�x���f�S�+J=Ԝ�,��S"%�z�5�N�pP���*jIM�?s ��=]�E�%���e�kK*]�5�:�g���%ID����2(�x�A���r�_D�P��s�9� ��đ���>�d�]up��`�Kv\����p!{��qG�DD����j�P�*�jf\�-��)��~��Y>=�k���F��>"�2.N���� RꚘ.�X�C��'��+?E�M�1��倓�G��f��Z�AU0����TdN�O���2��`��HQD�3��4�@��|��1A�$��2�Vr�Z�V�bX*�=��t�ZVfє��a����+g�O�%��`R�*^heb��0��cۼA�'N��{Z{�n������X�(�^ޥ �7H�"�/�B{b�l�}]�e􅥃�bA�q�(�d:N�B���]d'���u�P�F}�?>�o�D#p��N?���[���v|rp���s�>)]�6T����+7�8a�i�`R�	M�W�ӕ�QiJU�P#�<<����ͨ|�Т�<6�i�2i%���.l�E�=�� r����Ou]
qA+j6Y+��i�)�a�t���D7���O>S,���k�V�9�)Wq�[��(W0���ac��n�^t 2�g
/"/�W� �Փ�hȜ�-�-BE�V��N�Z��ld^ )D�	�ȅ���u�[�B��Y������ *+�B��	?��8�^A�f��(V�E���%�lxݜ��W�?��#����҇�' (��1pE�C��4G��LM���v,1Mx���}}�1Pi��7Dk�Lp��ȏ��0�bմ�|�ݩ����t�Ճ��NA�8��!���������P�~���3�k���a9���\���	�XC�z����4�G�%=��C�5e:7:1c���r�n���NYF�ج�ߴ��d:��#��H����׺� P��}���v���9$	�C{��'��E�<�H��6>�	��9�ύ�ĉԎ��D��w���;��H�D������$����^PK�)_�����W�o=l���$M|V��<��	����H��D�f��r�����$�d>�B�.�sCb���e|�ݵ���K����F����Yc�l��F�ͮ�X��0�`Ǭ�ȡ!&-�׏�%���q�lO��K�I|d����A&�UZ�B�+J4�+���:���ˉbK��F����uyT�[N#�|�]h�q��ߛ�pc)�#=_��`�8�Q����З�|9Z�oW��-�c}J����ʇ�Lѝ6��Y��Q<)�}�g��"̼�"cZ̼�g�<���-�lG�d����d&K�����&8�5����O�fvRW&�̉������׿S��~]�� ��2�޻�_l�	;�C����`H���]w8�@�).s D�>.�'�V���I�A�ABX��2f|U��P@}aXa�H��K�����j+����n��q�#3_i�+�bn�v�@]>h��e�PnՎ�o��������gM�~N'��1���a὾ʋ��;lf��8t��W>UjKV>⍮��ɟb���ۆ}��/"�qi=�o����B��U�y��Ba��E��B<���b�h�u�IA���!qpw'"�f#7	�����u�Tg}R:����k2�c��u=eY������6�PWn����N�_�]axi��*�̑�g!�#�
��yN���a1�����it\���:�bmi�A���2W����7[��U�1��1C��;�6���^g���i�VH�ջ.hlX5����c�J�����z�S��?EN���]���r�(H���{cl�V���d-��:ɚ�~.�_����o��ɐ��Oի4���1�y`����D���xx��󡶃WJi"E���f��;cBJ�`���bR�C�����"��7�@q}ϟ�P�"xP�e]��@���Ce��H�{�_k�J k�w��F]7�+%JH7�.O��6H�PQ>�/��~���g�GU��w=�r\#6�������x@4�Q �x6��P��k�'���V��z=5�+��3Ȥ���� B}�M��^!nPv�/t�Je��֞�pP��(�@���4Z���'��h,�.���.��ښ��.>r�# t��2�F۴Y�Y���g���i��2�p���5�ܒ4i?x�R�r���	%�?~]�9�W;˒��mɡ�{�i8�&M�{��{�l����P(�w�����L� �#�+���^�����ζ�f��D*޷��=>��tᨐ��<=u�^4�hlo�:���8��+;,�@�y
��>�6��4����R����<�~ei!�eze����l�p�i�#P�ii�nk;���p,P�K��H$�<�.���c�����l)UJRT��t�VKmlÁN5���5��c.K���!BC�w�ˀİ�����^w�tߦ������S:im�h�;<�%��FL~!�����e69�g��bW�gV�䌆�'��	B�f��@��}*Yt-Z+	/���������%;�=q��I��z�c��<����^�n;�(�D��S|X�d!��L/�4�{7��2��C��V����!*����쓣�goe��nXޖ�%w�8������[�� ������b����P��Q����*|=1���=���"W�=�������Ns�]�y
��5�/����Wr	ֹ>P�y+C����+N��f�-]-����e�C9��z�p��I���6-c"�Ao�L���T�36@.�)s���	�V��%O3�� ��I1�}7��IS͓�������x!lT��o9�d���QreG+�֫(��D��2��IO�5��
yR\F�mҔ���<��&er�M�|�,R��Ӷb� 3������^ۦ��;1�^�լ	b�oN�H7����0��V�O����ݟ �]������ �]�o�MoU�����g}Y���r��ZL;���h/� ����- ��&D&��dP�>s����i����Y�E�=���H�1F�jaM��%[rk��f��j~����Aa"�AY�x�!��~!Fk��Fu����K�3�����&Jan�<��Adb ]��F���&<��ИiƩ��+�:��t��\�a!���s�k��0��� QKC,Gw����Y��v�O��XW�)�q;���6�E�V0�i���M
=+H��ZVd=�\D#ЍO+v�r;!r=_rB�o��v}�Lu|��qsȚ%���x�ȏMkI�auQ*���dvӥKLn��űn��nՈ�*EȻo�?�0��z;���*;��L�tuxa;ϧ�6ꄥ٪lx�d|ژm/n[���[�'3�Gc�9)
Vfl��fk����6�)j���B=��\�V뜨�`7и1տ�v|�?�� �r�Y
{�f�����P� {��`q�7��|���}ZNM�A�;;��>��J�U鳯�'n`\������Ĺ_R��K�+��d��?�%{�'��3�%�V�A9ч�����=+/� lj��+0!�)�hkg'��׺n^��;?x�C�!t��k;�����m�� X���$_a룱s�H��Wsz�����A`�{�d�zoQ]�ȕc���:�Y���k  F�?�����|���V�?<?K�t�u�ײ؜��})����\x��l��K�f��!q�t�Oy�\y!��:E�����~�7]������sa�����[��s��X�-(���j�#Q�����9Ri���E��%�ӆBίSϬ�?����'�(�~���YtJ�c��dyo��&��	oQwq����-��>3�?��
*���/{0��tN�v`��nHh~A���V�0�����3��s�RPJ��j=�WMmpn����XD	!�lDQ�tl��b�=Ǒ>LA�W;�1��,_|�ǠbS�{����_$�y�i�k�
�Mm��i�1�¡ {��
�I�.ic�o���k��~��k@���������n�͋"�й��1����Y�o���3��#�����@�G�n���	��|�9ҫB�����[+��PѤ��� YD�3 ����A�3|�upq�\�>/R{�7Nv�	X�5����xA�+�֣}��^�Ԅy�YPu�$����5��+�������ؓ��If{Y__9W1W];s�`F�(���:�M^������Z��||�V�����L1�ZX�Mp�=V҄2�g�T��u�=���4���E��ݲHP���u��o�T����RHz/��}b2ҵ�K���Eh]�T�S:Ț��wpZ9�"��鴡����������(�E�H�2�M)�~�l��a��-V��WQF@V���t�V-@:�0c#u�>���X�l��f v¢��7#4� ޺]�1�"T��Qa�un:��=*|"�L݃)�ک�~7Z
q����&&#�"��	WVf�E#��?͂��ը�@`��继�|R�	#��y��[2�{�Z�U��m%��	�ЦN�԰{���R$:�!K���"��g�=���eG����Jy^��r׻��:�C
�E��Ħ�I�$�}�fI�E8Awe��]���FH�r�+�u��(f�\n��[�T�������[<�:"s�}c��+M(آ�3 ������ͪB�9�a���X�W8��<ײc%��3�ć�ӈ�SP>�88�8V��-G�
 Guz�yu���� �J�V�Y�<�C���/���}F����m����"@1f��*d���8B�% `i���[2AМ��3D�oJ=]@y���٩(�9׵=A%n�b���P���F����1����JJ�S=Y�����.=�_}����O���u�4@�f�v7�2]�0�(l*������p�ruJN�I
b�uaq���
O������o�]��0���0��]�{J����d��%�3�/�_������o	�����rp`V$��=w��}>ޕv嚩}\_cr��M�!����kf3���,�d���~U1��'�7
�H�-�K�%B=� ���r^� U��x1Z���D&yOb�T����:_�����eGq4�I��5�o�إ��=�\u��|#����;}*�+�����*<���N��@�khԂ-<������XۄOȮq�����.�bh ��g
"��d��)�����GB0>{H�}�JR��.19&�ZO(��J���J�𞃳�����-����h%���"�Kcm�
8k���b@��P'��nl�a�\���7d_O���qQ���vCg<8ϊ��tHhW�%�P�KӾ����m�S׭�o�@�H�+�����9�h6��ȇW��:]݁��It��(��ad	���v\�"M�\� D$rxm��]hV뭚�Z9;�N�D�Fmo��(�_�N�þ��E��VT&(��x�;�!X~k�kkc��)?�4���{���@��>��NY�B�Wjz�U7 Эy<�E�9�� $�����}�3���/a��E�KY���B �w���j�� ���Q�XI3�1�P�!ST>��1��d�^�\�w�H�y�&O����H�>)m����N��J@ ��h�"�6����0�����;W�憡;R���u�%Jy�ln��������dV��,cKE���<��I(��ގ���F�Q�ߓ�!���T�3GK�ң���/^^9�zҰ�qY�"SŖL�e	ɐ��/E9��Y����<�e��J"�I#NK� ��hz��`T�}�pp,�;i_��yR2�Yxm�b���@����^P�g|����msr���9��G�BA�f
�_��K�U�JbDa�����ugi���)Ql~%;9&Rs�m���űl��L�T)6��1*����� �|1~��+�c�.<�)K�
�X��� ���bgR�;�L}�%ٳ��#z�Oi�ߏe?r��������^ҋm?����U���'��c]'1���W�1�vpC����g	g�oIl����q�gw:�V��!�~��*��8���g�<�BU��5�лfؐ"K��<��P�l�#)_�<�p(b~l4)��H6��}�'���w�4IRO�F,2��Jf��_���Y�+\h�(���Ţ�8��Η������r>�(aȇ�X�]��<Z1}{m�����p������9��8 ��b�PcMG��4�M'���+qՔw3D|j��T�E3��P�7���0C����_��0]ߣ�{3�a�ԉ�k8 ֑�;Q��n��d�ᓯ�i>P՝��gP�{!S�>�n6 ���qy"R;�
�!\�В_���;�j7C"��G?��� ��U[W�ԘE��
�N����cהk�� �����k���]]CE	62sxr�� k�_�ޛ7O���%��|�o{��6�������A���k�n�~�)A��P�4Av: �:�fx��҅�m�O��u�Ψ��p�j��p�
w׬/8KݕA��c� �a���=�6�e�4�5c)5��f�@�����V�S�.Wؙ�Y�K�4�k�A�;=���'��h�H�F���L�q�� �YpXC+�����J{h��坱0]M9Q[t:�K��˹�]��~ @�[�tm��w,�4�c�g�E�ի�!�K�-�^�ja|P��Hs�bH�9�M����9p���!���"]������T���]֟�0�t2!�Z 0K橹�����%d���@	1Dkͪ��{%��7����ZY��,1Mo�\�����oU�i�~<�8�*'�SѶ_�^��MB,�M��շ��+��<�O�9���WhT�O�k1f�c��42���f��*J�@���8H�Iw����<�H�tz�9�E+_�6�<y���c��l8hu�;햵2|s�]�Ϧ�0�ARA���F���Y �/�t�;J�}0j�#=�2��o"W�o�}��3�ٛ����q���8���Hcunȫ�A�23�mq.��V�sW0����&�5�b�^^��*��ٙ����v�c��\��qA���t�eB����W�6(z�>"FޮQ�!�Ǌm dh��������t��n﹢0mИb%��9,������
k��U;hY�Q���~�� 8�e+Er������ՀW�Q6m&� �#6�k�T�Pz� �~G/�jzeA{�54�����T��,)����K�t#�C5}��<4��.�Lu]�K@��A	���:#�/g�(؝|�\�����!\`�.�uւN��'d؊i�-ҽ�FE�͝M��w����*�H|L��5Tֲ6r3�f�)��̸��ϒ����]G����O�fHo��9���Cx��&5��(�H_p��UOE����"E[������^�*$��?�>F��)L5�CЉ��r����@�_2a����na?֋ބ�b��`����X��GSh�<A9h���+çU�r#j������ܤ�JS����K��-C�8{�ڳ��f ZgU�+�{UO�*Y'��匫���\�B�QT�X̟@H v#�a1KT�}��h���ϊL�����oP��L�O8�T(i�XRـ�(�Fd�3Kh����^a;��J�8��.V5 �T/�ǲuM�봑��_�
<�.L���>:�G�5~q9����N%G��c[~����� x�Z�42��u~i;��؍%
P�5$"^����A���{�"�
���So��g�KŽ
Z�����(�\�ȗ����^�C+>�H�b���'ˬ6 ��4��3�_.KA����DR�ChC��Y������$ݿPY�i�����v��8���X'#���W���2q(�DN�A����S�Cg�{� �j𫃸I�x
�/��Oya���&��{!w�p�e��_��UxR{�Fx�f�����6������� _��B15� �W�L��I� E�f��P���'���CHݾ�����+r9���ҩ��N�Jm@���V&�b��9�w.ZO��&]��f}?Mvx5��W�7~aJ�&Ѹ*�}���Cy?�k���i�n=����b��Xㅅ�>=��\.N��� �H�������jy͟�k����CɓY[��E�T�T�t�i!t�tx{����xP��x���"ǷĎ8�^i
@����H�y�Z��t�\�+�\J�l��@9a�51���?5Ѩ��uJ�7�$��Rr[�]�����L�,��G[w�Y�Ea��2l��ʃ/��͌p�!��?�'d��[��vA������in�j��5\g�}�P�LM2�O�����������n_��َI�٧��."��H�Si�	j���b��%�e�.4O�`�\{�W&"Z�3�y,1}-�Շ�@.���Ѯ�a��)��UqO�g�gf�b�@rX@S�Ia.�â��������͊�w��A0���`�3W1Zu��g$��R5D��K:���w�A��;&u]p̠ͤv���]�2�9�6�G�}؜�!�(H2v2>���!�5��@��q�6�Q��+�g��ɲp
f�1Xo't<��.�z������y5Z�7�4U�u5�����C���h��C�3a�����NZ�By8��_F�Vd�� �ԲP�<�)���b����zd��F��H������|�}���5:� �yP�w�+�f�#�Q��h���g1%��b�Z�����L��J�4��h�01��SN��0�Q\�V��С�ы�`��a��Xj��`ǀF�9�Sͼquǔ �d!�(o�2X�e���kt��W��5=rw�,���|t,����X	d�����}�C;�i�J�����ܐF-�I�"tY[�__�.rx�|I�A�{6X	C�8%-1G(��H��E3�b|��+�m@w�\Z����)8����,��
������?2]��nk�N���A$6J��i=d0��*q�:.�e�s=�aY��{e������� �i";)�K%�;`��T��F��kx����Qն�!?U�G�J� 	m��^1�vC�b�d=����������
�@��k��3���F
�X0�M�̬������ܛ�Y�bi�����p*��ִY(�dd���x�H��#���B�����b%�bJ�ԋ�ˡ��$V����o2��oR[v:(�!��ۻ�%#���:!����d��:��7P�abJ�f�p���W���fQZ���*����
d�h�8����te�\���Z�Q��}Iw�����=c��؇�!��%S�3��]wC��d�!�d�5s��`��8;� ����U
<���m�1�
ج<&�6�(*�iw��D��#�bw���բm��X��Of4��*�2;�����|�����Ҡ>���68�R��]մ��-q]B��͍�؜�Q�3���^����U,�(�g��jṍ������z��������y��o�D,�|4Nzϧ�<z% -���"�n�Ҝ��6ƽ0�M:��3�v�J�:�9"ك#�{ё���N�`%�b�
䍇FGF�>���y>X���R��ŧ���kSm���}��K�\�L�����OY��K�	��6q��}�&�R�4��c�	fߴe���c%]-���𮤦rm.�����J_�i�n:3d�=�QCq׹��?�o����(�V�������F)�V�t��|��k��)�b�|#B�N�K%����^NX���R�)�.���m&��*��1wO�mʿ����!�8|��%�.��%h43BCs���&5���y���hW�r6�&��
�sWo)�(\�[6B,��a��RE�t͑�i"q�:����-�M��'q�z&��U�sg�&�M+�ӫ�>QS��.}�˴ �׸e;�$?�D�v�ҨQT�L� ��S���Ԗ�"!�䲲��:�4NN�ӳe�\�j	�'��Z�����(��T^�|�?q�-ŋ�om�ߝ���NC9W�Y�.3��������q2��n�Vk��m�zY�E��}��0 �E4��V8/� UJ�Qc�w�C�#�'`���v4�i-�P�C����?����=�yU(>�W�7΁wp����ӝ�����7
������*�VcuҶ���I�x~v�iP��g@�nB�~��o�,��˴���G�f��j,�CC��	}2��������N7��r`���0��)/�ƹ���L���d��^�HR���_�2�A �ޘ�xU��4W��{Q�tr�������r=!^�U`�4<Y�y��#�v�K��"'�)���\�����@,�p.�����?�P����Ҥ�M-��<��ۍ�|�4gL�,X�n�r7���N0^
zP��v���I'(t�&y�7P�����0t�'���gJ[���tyu�/��G��@�S����9�[_ ��r�F*��ǽ��HN��?x�v�B<A?�B������=���AgLdS&�e������O�Oa��5��͉���E�	��2�umG@`ZN���pLFU��q��>)7���K�;jV;s� �a�e+R��&%X* �P��W\]��p��J�Ȱ�u�b�s���/��U nxYo�&PTpY�)�X��"g�7�l�~�Ι�l��RN|���`�Č�ZM�K`5��}jo`�z���p�Ij�?W�)�WOԎc�����=��&�񍭏)��u�z�.�<9��_4>zfh�c O�{��CM3X��6G!M��mW�Å��`X|���ڔ�)���q�|���k�/$	N�z��Ji��D��L��ƣ[R厂^�v7/��wu
o@��Ġ�37�@��D�Ҥ�V��[ہ�>Q��W�UKP��0�v�p�˥O�Hj�;�vɻ�i���є|xƮ	6��_V- H�v���۾� �77��Wǰ�m
��}�O�`��st�ɷ�1�ůX�!�PO�����tq�L�Y2��(�]�))Ay��X���c��O�����/޼1ҰY��OA�g�(��n�k���A�-;�A������\_�,Xvt(oH������(�V����6�*4�Q`�}�Jdr`!C)�C'[�b|��"cj_ao��*�1�rʥ�+�M�N~�;�c��`x�;�PM/b����������G$|H޵��v	M1�����z�R0�;T��[;�JZ��8�L�`�A�|���5�(���?M?�_ƺ�J���S�%�)�@V�uְY+������S6��e3�0p�O �$��8/����@�YN$?!��E��5�� m�6<0dG<�tƯv,Oxm���bV�ᩌ͖z�a�u�N�SEq=�f|��;8@�����������.8�oU�9�7��6;�-�񫀨{��N�����r�C�Y�%6�9�F���[O����6�5*3K�
\?�Ս�c��,J
�.Gׁ�t2�-_h�N��.�a�&�`W5�fW� K;���IV|�RCa.T�O����O�@���^RkL���&��c��TϮ�ܔ�hA��cŕY���� ����Qc��g[������~$nL��W�O4i�������l�QY��I��[bn�U�[����{,�AZ|t� �aqj?���柲h�O�=J��/���וK��K�Zc�I�!8Mt*�m�^z��gW�楼~��FT�w�H�R���T�!j���J��_��]}�H�_����7�c�A�����;G�ƪ
QC�B�}�������=1J�&*�eqh��X�
���m?W���Ė�ݳվm���T�3��/x;�Όz=G
^�t��ٕ���iN>�8:1��4E�Eꞇ�]��(�Kf)�{�Z�Q�{�6E������n�K#�s�eփ���YLd�j���X#&����y	����"9ɖ����`�x�H'�\L{Tj�]�S�y��=���QӮ3��e���I��D�,(k������9@]�@Z�e�-�S���M��6G$K�>u�lj�����>�ltX��+�!��S�{p���f���.ș��kO�XO�y`�/jF��j��j3�k��&�̈[6� 1*�3�4QrW�%��9y����d�I]ɐ��id9F���Ʒ���C���F�K�M�E�����x��B�ɱ(���_"Mp���'�ʜk�KAA]����gƴ�zg(�O�y_�`�I�B���N�D�Š�?��$�=[�Gk��
S���-c�����yzc���V��}ݟ~�S }��ޔ�G�K�gجH�b�
����u%N��:6��"�͜R�t�q�?w�$�ܚ��6���|�/&t�́�"ž���b(��*3��<����}X>�{�N��,F%~����(>�a�/ڌu����x�[��Wl@�������WC�:<{��;�d���z"�I�FL�8�f�N3C�8,�Իh��Pi�����RD�&�۵fjx�4+�O��8%%J$��e�:�Ն�� L׾:Z����cx1/)"�D087Ht��)��~j��V̙����t\i�H��,qd�f��b�WY�Ρ,�;�^���7�y��z�e�ǩoz}<W�`*���Υ�b\�,�Qwb�zY����N����PP������#�'�M�����'���V&B���+|�fS��:�d��hw���#i��Tkԛ)�	T����$.垉w�?����:�W�:���h�a.�{q�i�GsZ�2Qi[��k�#D��݀Q��&�?� 6�g�JY��g���kӃ8^`3p.�h��t/A���>���:_��Dr�W[�N�`	Rl6=�n2�-D�8��g��$�]zΫP�Ğv5vwH&:�Rñ����~v��;;5��]W�1�pxJ��w��v�'9FBO�e!��ܮ�fL')�̚��b��*Đ��N�?�w����o0�l�L[#M��=����̆��
��W�YC��3ROGKR%�u��>�oB�DT扆Hw�MR� ) e*����t�����`Kp��� �r��,���f]e���;g�a{��8CT�Up�%Ā�-}���O��D�*���9��v8D���yl�����wKԇ9��FZ?4�U� ��fL�>�o���� �!b	uNo�$�Q7Q.�"U����O�!�C�r�s|%\Ez
|�f�V�ӄ��⥷`�ٻخ��7���I]��ݰȳ�Y�8ܮ&?��7�D�e�~�h�磩�1^�3l9�⟢��b0�OȾ� O��A��$1�<������=mFb���.#-&5BGMQ��s�)-��SJ��q�N�����e)�5v�>��������Pj7=�y6��n�xO�����4�߭��$f�<��U��Y��?,��V Ȥg'ຬQ�<����{*���,���23���*� p8�W�wT�Q��i�����pX��b�ߊ��$Etb&��L�3��4qD+�J�fɤ��SO{o��ч�w���k&� �9l�9[YA[I6�uj͍ �[�X%]?����	�8g�t$���L�j�6�c��~U`�\(��R)a]����;��!K�J���$�jP���J�������Zn� oc��MW(��c����1�v����Q�wwóڽE7��Pd�SCA,B5���y��!��"�@�S����YQ�\���o�T�$CMı��f�����r~���S����u�ʢ�;>3�$�A~���ؐ�|� �n�ʴ�~�5G�ZB�X�1�F�^7?p,
�}�-y!%J�/��*ei��x��cP�=D٥�u^�7WS� (N���z��P:�'�[�u����=�LG�<��=��0�&����2Y0j�/(��?kNk'g���P�ɂ�&n���"��с���XZ��|��`�Cw�֕���Q��*'�+���WI�5�Z��tL��D��T�:|����EE�]g���V��+Z*�>=���C�)�[��߽��o=�ע1 �!��N���>U�!M�d7=�c�����^���|)H���M%O2"���Z6ݤ�Ro��d�{PT����q6�փ������ ,-�e�?g�n��HD����I��w��|s��B��-Q҇�E���(%g͈?e�8eIxX����$2p�J!ga��c��
����7G�����y ����m @WW���F��e7|�|u7�<�'`�?�A7P�ֽ̊�����k�g��$�Q��-� M�-4���J劽�s�كn8�j2.JC�������&�h�V��]ma�j���Z��&)�_�����bJ;m>ۻ�y��C��D�N䋙�g(�V<p�����x#�(G��.ph H�K1�&+��2�F\,��t������nb��r Z��y�.�t^H}A��Hˈ����7���=!���\��ɂ?pTN��l$'];\N*t��!���~G���h���Lq0X8,�7��P�w e����x�]�<���<�#1�}����뒠�w��z�t��˻�q������b�z;��kqԐ���>^��h9�dF�����H��� ���2Q��x���Vp5�Q���NȊ �w�xyZ_diX�����f����	�@h��,����6�t<,���_�|m�'����fE�ئ��k�д�p5#V��pm���"�p�|CKCmZ�f�>�`晢�Zp�.��F�6�(0��J�B���^.�7uc��TE��8�����ez�e� ���:h?�������˝OH\\8-PmXz�&��WA��>p����u
r��=ݷ����A�<'����A�hKjHy'��6�%�J�����6�W��R��*���sc<EiW�3��?��Z8���(q�}K�`�st3�W���edNI�*g��_�m��]�<�_9�ǌT5-~����Z�v�V��:A�S�O�`K�Z���W({�ȯZi�plj�{�s_lS�e%)v�Μ�,�����pc�yMs+��5��*;�k/����+C��@fB N��Ǻβ<���ۥj����q��α~�hOz?�Yu�~NV 3V�E��C�Q���u4��㌾MD3�7D�+���I5pt����dв|x��>���
�����f��É솔��z�R� ��#X�~���7�1��^�͜c$�sl_����V9PJ^̻:�����;�$�h�?��7�$�j^�O:��~����'EI@OH�=w�Ky���47��/g���EYI΋� ��CMpQ�:����@寏G$G�o����ܓ?�o�n��/q*G(j�yO�?��sj5�U��Raׂ���=�B��@���*f aD��|�ǽ�� "*	���&_� �t$
�Bd��ަ�e��(ҷ�Ķ�t����E	Cn>���6��	Ǡ�zs���D�TO�bEE�cw;-�P���7����>Q>�^�RLGU�Ƒ���N˅X�m�'+_p%��o���ɓv���?#��qUn����Au~^��1S�_i� ���X�6#X��f�(JU��� ;ޠĠK�����3�.BH�=�e2���"{��=�ĥ5�����#�+�/�dZ�%b�{�`e��[�n}ܕ�6��w���ZI����$�A���|6�g�M�|XP
�Dg'H#U/�ӌ&����#ݖ�_�D�2H������*��S����@S�M"M ���M�h�{�0Pq��;{����� SN�_7�,�?uRS0ᮧ8������K,:��n��nĳ���:w<���A���}�)��c�p\2�[��A���Q2m��e��+ļ���IƞJ!���å��p�Q�ҞZ�C4��)���/3mR}�葬D�F^s���5L}�~i��f�+��ZJ���0d�Ԣ����i��_��zxz�&Ir0ޣq� "3���C���F������CJ!���$����$_�!�����De`	 W�z��81�0�](�)���F�!
]�O`f�i���L�^�J+ƺ6�l-�Q�f~Yf;خ�/��\�Y����w#�?�o�����|��3<�m����"#�Ë�!�hb�9,�N.�N$�&6s�����pӰ�Z4��^L�ݧ��s>�}\���?x��ҏ'�+-e�B��'����ς�q�cX?�6�ݬ�dt�T�\��2��EC^ӥI+��r��? y��I�sb���
��R6�Ѱml�d38pI��� ��#��*�<�*�8�@��vPʃ-�Xha&�p���y��'k��� >o��ܔ=���|�U����{ �x��D;`�3 �gB�	5]���/��%Vc���7������DRV�*�Ա�?M�D�x�29�VX�:a�biD����D��χk�+��Dq�`6<_��O�l�mEOJG�ҽV�\�fۆ��p1�eV��� ���o'/,�ҙY0�K��5,~�4d�:�����a��5�q����i§_KgT�C��O�T�{���e]�[a�$���?����|�pf�uzXPϣ�<o4y�V$7~(��՟����*J׿����9(��&;\(p�������Ìr_BD���GM�B�:�
QT8!<XL#͞�ݸ�>�1rp�h����S�x �%���$�K�T��a���C��5�>�uZ��Ǫj��_[o]x/+j���C�� )��I~u6\^9LcFa�8�b�5ẋ[f�d6�r�YO�5%+��g� �R1�_2O�^;-���4����J��������2��mT�u����B�U�1��R�Tg��=��w���/�omI@�߱$��s`�C�ΐLD9cI1�n���S�^����`�|]M7��U ��'�����Hc͡����10I:�&9�0�:` [�4C��3�M�I1�$$��y�H�5d
���o������������j�}�q�~��~a��sZdp"X㦗 ��+�Ē肵P�ɥ���Dd���?�ȷ1^��tn��O^v"�~Q!�kr�� KN��P�{��TD���|���F���Mɷ�J	x�8'�cF��:*�i��?�'���<�ySM����Vs�/HE�cxP\0SS޲`�����hR\���jէ���[H���"p�^<��.W(?g�o`\SvU�z�lH�ۦm��A^l-�9)P�$�;�G.�c��K()�%�O(]��k�L��P��xX�u3ܤ��: ?;LȀ����ٜX![��Hl
ĵ0ӹJ��P�\T�Z�}�5�3��`�O�#���5���n}���C���AB^�����K�ڭᐭumHK�8��ܕ��-���u����x��u���겪ގ�#c�X�Nu�o<Ʌ�V�:Le��BYVW�J�7c:C����*��:���ջLҚo3�8,cmb<sT�c�����wi�W
E}2��cW�B��Q�b�z�ۈ|���Sg]Pb�P:�Z-������䗵�j+��Ŀ�UrD'^/?2�� x����"n��)�U� _Ͼ鳾�A�T�m3��ݏ�o��A�Ѱ��MF�<�l�+8'��x��ۤ���*WhrQ�/���b�Q�8���'�{$q
�2:6R6]r(,�{r��we$�'�%�&:G�����s;��q>�_m���^ڿ�E2���R#{[!�|��@j�d�����R�c>�D�1�g�_�!K�w�hj�J���V=̿<K:�q�O?f�j�J��T������P㈊7�����	w�Y�^�r
O#��Үo�&3 T�,N�P8:���#*N���+����C^�域�����N���꼡��zP�:)"���⬄�c���^r$4e�#k�Y���za��̻6��8Z�;��[��C��+�*S=�Uʓ�ו���?J��Vˣ����_HS�uq�vO��m�;�r�b�@�b�gt�t1��N<PJ.?XiF��O�Q�l�K�DOLӇ�ڴ*̷.��Q�5F K՘˘rS|�E.���g�G%t����ʛ� r�ɤ��9
��N��rѲ� �!o�Ҙ��f�j�`� Z"@�+�a�`#0�V�mb&5Cp'�Ҡ��a�B.�Çn+��=u�̜�K`N��Q�0xChǉ@��b�=��)�"�ɉ"=f�8��+	��4� ��$�
�.�{s#8Y��q>����mOjh˹�\HD�f|B����	��x�M<��l����^{���a6rI��ȀĀ�-��
9A�l�"2m�Rd�L��
F<���V�t��6p��|�W@��~nW W/nQ���l*o�Ui7���OxxMև�m}���2B�C��|iu͘�kFrՃk�¼�n�[���}�,6��%���N		�>�c�\�E }�}?J�
wc[߯�Re*45�M���$Hr-�d�����v8=�9T����f�v�1��5�c?�� �I�J��o��qqm3{��J�=������E���-s]S���	QMV\�>Nk{���pk��N��* w������K@�܃m��?Y��V���5��x<���KRFx����ӫ�v=��xW=�F�i fy#xav{4��$*�C�tn�K~�x�>��� ����-�u�{t.�-�_� %���:����e
� ��r;TLKJß�_]>�[W���ji�z)P�[��9,���GJ��G�� �d�p`t0;�vþ_&���c`"IJ�t{.�^~ZJ9s}��Gu���r��m�.T?T؝��o�ǭsÍ�g�Y*Xb؂��Yrj
��hpo�b��yngv��2j�V��Q���Y�9�<���J֕�gY�6=q��d��o���0��^]48R��G�e *޹����P�8���C4u�9�zP��Zڢ�a[�X���%9g�<���M�/ٽ5�&j�=�eHf*��}�d����A־DH��}�� ���R:HZ�S���p��p�o��!XH��঄�Ch���J�m�ڲ�Y��ū`��IL�K���Y#h��mf�`�/i��v�_�D�\� ���<��ج�rF�l�E�$"�D:�YV;4X��E4< ����Ӓ�B�%3]���s����Ni7K�E�.��S/[����O-���IG� "�*��T#�u��@�ۡ'­�Vw������� t��	v�[x�Bo_9�]���yŴ�z��:!�[Q����S������x���� �|����9X�T���d7 EE�Ϟ�m����!���jafh�I�1d�s!O����6@�U���Ğ]��3�͔�U�={gʅ��
�T��P�����Ko�s.�����]h��_\?wD�����J��������/9���<�	��M/g�U"��ϛ��nI�x�a��k�ᗈӦ��x?�i�!CE8J��Λ��L"H�aW�'���|_�+?�o�X�jr^d�Y;�{fp"��%�<�p��֞�l��K��=j�~�D��oo1M���Y�!�����\K� r��� =8EW���W�ڒ�A�W�qð��_��6��Y�kjK�	���:3MG
���}7�+��+�b��
s�[fٟP,j;)���&}���2�f�*'1&�E��}���4���8�Z(7>5�����͸q�Y�JX����\H��Q����b�'#�셓��.��BY�G|�&���d_ݫ�F���-K�5��8<Q��/=.%|��R?�nPh��3�~j7������g��uZ��r��7�ka�E��,�[�$�����B'/�:�4B�C* ]���s�M�j.?�薐��Dk��+��TOy�cu2E��f���c��m1�(㤗�^g���vzz�FI�Π�F ����Oo��Ł%�yQ<�Fw`�T�R���4�|�N�s�^6{��dO��# �13F��BS�`��l 6y_؁�r��-�VY��\x��?G�vE�u������ʅ���d��A�0w[�^�EB��~��ڙa���^�L7]�.Z�~C�zUOz�t�۱U9j�f܎�f�*���|��"�����w{�Û�*J/�����Ѿa��^	l�Q �k�G�) Y�˳{�n���|D���1ҏ�r
&q��F�:~sI&8I��rg�{H�f97it�,�R�a.bV6S��<���ă�uNyPK���5z�RH���M�ar�<*��΄:�Ɇs�����4���EC4�1��8�C������Ktt�i/�S>�����҈3���1,�;a����*�UP�Yҭ�/@�=��OV�����j%�vtS�n�1 Q��؏�\�ħh�YЫ-?���v�Ϛ���'/^4�{J����B�������VSaM�WK�0�=�(�9[�o�kZ͠v'����=�@�����4yѕ8�y����H�jQK��������q�˪��T=��Y����� ݽ{~,��ǔ�d��!��O�j�����Ae#Lt���pv$�e\��:�����ghh�sب|45�N���$�#�8����Fa�|�Wa]����=\E�ǫN�jJl�XRr��E�8e!�Eވ9�vD���M���P�jg�j3)����±-�QJ�L�):���VpC`cs��K��"�����SR�e���C��O�D(���GY�Fp 
:_н��2%����qo�/^��vЎ^������#���Q�o]����j��c���q���K�\}���R��_��Ѳ�{{��T��bX/b�H\�*���M���A��R�.��(�c!Y�k�C��3�;>1%��)o�.��_�*���6����٪�{�떂;���a8`�[�g���u� �q�pQ�L�8j�	�t�d4O�Xy��I]�W4����L�nW���\u�B?/�e�+�¡�xX�F��G��⭟
��P�*NO��YY$gi�Z�׺��8�\a�P��-4t#}�"}n�>9�b?�$��������sᅇ��;��I}g���58�?wumy]�V���m���;7��/pB*�N�Eq��X	F�h	�s�񩃤�����.��օ�Z@��_�7��\+kv~h�u{�7,��O{͊���LdW��$��k������k~��N�]�����My�R1rg�F.��j��~��P�L�x�:Yts1r�8�hi5�p��rL�Q5�l�8Cj�c��:��T\P�Ws�o��Ӄ��T���'Hn׆#�~fs8�M��<�4-+q`v��\���	�͍܍�1�s�M��;�S�	+�Ē�:�#נ��X�r�{���i7�j6�)�khNu�PV�UA���&�0/����4Z��E�F�vo�����|��Ar���!5�n�� �B~򀎓�*�C��RS=�Y��a�!i��kt<��Y49���[��̭��xڢ��`Pw*+�9�W

�"�u���ZD79 ��o���"LeQj���%���f���~��MهE	 ��S7�*)mCv�UX-T�K	�g���G�HU0�����"Cg�dH�>�Y��mV��Fg�1x�%�et��e.�h�RTP��)e �$#�������� ���Bͬ�������@ɠh��M�і���>�;\&S}�&��)��������Yt�*y���C�(��^_���%S�����OlZˢ��]�WF/`��(��F~�-�����'^�-�x	��YFY�� ��l�UƸ��7gO"!�ӟ��<BzӞݻ�����k�rY�D��̂��2�L���yV�P�"_6{��7����.�[+�ZPf�rd��k٣z�D�b���uB�@ʆDͬ�Dg#��C�p���<����ϡ��,�Kql�M��*��Eء0qh�	��K@�+�l�op�	����[8�|����.��b�sR�0M�]�z=3&�^]=�4�o���.���kB*U��#i9n�j��������^?�7�:}�+G�ulF��g�C��s(B���#3�B���wBή�&e���6��]9e�;��]�a��u-~�rz-n����;��׏ƅ����cǭ���
z3��5��E�:[���6�N	6��e��A񑦌�z���
�P<�{_�49UF�v���XW||bt(l����;���_-���m�O����*�R�u�G>��ݱF�D%�Y���;B��k_�O��[��u<�U'H�O�5o��͋~z��ǘ�>�huk�e`φ����r���U�l�' 	`��==_�u|	������h��Q�KYP<,�W�w4k!�J�v�fv!+���*9qH���/���
�Ҭ-�iZ��>��&9bV�g	N��-�.��T{4���"�ɧ��)�):���uS�G�V�z,�A�	�h�S����j0C�J[7���oʀ�H�6��3���3�R��U�}�����77�u�UGa\N X�-���$�������8�R�Y�2Ƣ{:�)����_�ޏ��TG8)u��d�ysj$q�r<�V�O�ߥ�N��Hvr�
6����pu��XM�1�pl�;���{�6	��Zϸt�T��̺_�>[��h0^���2�t-lZ�_��.���b޳ǩ�@a�,饰4d��s�r�ٴ��ݠwsZ=��z-�Z_\�c*�}����EN�HДG߻�gاjV�No���W�Ҕ0OȾF��:L�Cp2�Z�6�6�Pr����t���-�]�{����Ζ�=��2�� [i�RP?3�U�f��uP�����G�ߨO4U�0@S�}�Kh;���s��5�V���K"aI�B��h(
Z��ܦ`	h����}]h � am��B%�"Xr�3LT�VH5Ѯ�[Qb��Z�8}�Vk�(�o`#�_�9���߮��Ĕ_�k�q)Bw¬(/��s%LP���\��s+hb�����ԳރK�T�i��&��:2�\-�C��1E�x	V(i��/˸���_������;��u>�_�2k Li���=񳧪\��
'<��Í�Q"�О^ �9a'*s��H�����yI��P����Ȍ���SX�����V��}����6Jl�y�=ɪ|�#��E�B���+G���ѻ��`���2��[����%NѴG:�K�.�5�6��a\���؎����S��}I@�:wտ��]�.�|Q:��A�e�ˊ�[�wy�p�B�����y V5����m�|��w\����_g,X�h v@��V��a.�@ǽomd^��'���r�+�':~�f�TU���%v���=|C5���M6"�Hhp�]�r�{}� ��#&��"r_b� 	@�T�l�f8br��]�,�9Mndл��NTE�~=x�GC�ʀ�f��'�^-~<�I7W��0��G�Qq��A|m\#��d��_%��U
o���A���!Ɏ�uFW�2N{���Q�̥��a�#��}�F5e@:7U4�iLu����ĭ��]��
DD��6��ͬ�-eg�GX���� ��]�b-e��;�0`�����ah���*���-4٤I�s�n�<9������F)EՓ���'����:p�AF�NT�P���x鹋j+3�[��&�{IΐC�o�tzS�ߊ��$!�ZL/=��0p����$|rAZ#��<޹��u
�a�"M�ףt�U��K��j��KO�#�x���41�Nu���Sr����~�
[��!��8�m pG�N�<Q��b�v@z �)TOٽ[)�����bh��D�}�6�:o�뽩���
�~4.G��g��Ml����'P�<��A�6���\t�,�l����X7]d�h����%yq�;,e�I73>q-h���%(6mQ���e�3h|+��� ė5ć�6E\m�{9�T�e�����'*i�ʧu���0e.~â���� �r��ؖ,��g�s����8�r�U�V09*ꍦ�{�_���(v^%�6�x�ߌ�eA)���$\K�[�BF}U���W𨝩�R}��ɐ�;sD������d��Fk�����NջA*��#S���5�{^3J�i�%��8Ēܹ*o���Gr����o9�pE����s��������T�������d}�8-$a�}���a�_���b�Ժ���!nL���# ���P9��'>��dc^%��I�V}|���L.Y��v�y0�F3��Bo�E�N$�o�T�~��PG+2p�!��%S�-1w �y.����0�؆��#	�9�)3ӗ��5,���}��%@�z|��p�\5��^Ӻ�(h��z*L���e����<��/y�g�!>�B�?��;�A Ď�i�S�z!=d�� ��6+����2h�g� �Cd�?w�v�\�kes����3Y$��r�V�x�M0$B�fd݊H���&�q�z���M`�'=Az�	c=.�Ԃ�3�2�?&X�$-��/G?�Oq��~����)�+�/MP핡h_>��2����#Ț�h�|�<��	�j��V9�G�ueP��BL�a�i��_��6xi5�wL\uY���gi0��Cʷ==�G�����/��_ �E���v�Zb����9Pz��*�a"8�oB��mE+�����V�$[Vw�T��gq:AS`�<�r�)�CBf��:A!��T�������_-s�lԟ�*��r� ����j1�Ub*�Di��r��5�U���%�@dMR��<v /Uy�"�v�;�F-��/b�?M�ֳ����7�����G<�@l��ed��#�W�V�J@V��晇g e,�O���v��q�j�M�*?��)a�iF�� �[8
\����y5��%��Iez| gl�MWb�C�,�zU��������u�9m0���-�ڃ���)/�#�<���~��n��b/b�7��9����%ޗ�_Y����Ѹ��]J%)�Y��ы��,yC��&��hhI����-�81��v*�a�����ٷU�wϧZ����w0��{����'�@Y��H�N3��@]:QL�iX��u��1.Q�͎��e�U�����<�`�����j`�~E�7{�Mk�Kko�8ш�^p(�Q���6덍Xzq<@�p�K�������K�LQ�
i�K�t��;�"h-��W��"0\�0
~ޢ���^�˟��;]�X�'A�����Qj�/�_&/amS�Jۄ���>�-�%h@�1�h��)���2j��WmA�?�8&�]&�����ff�.���K�6
�M�/a���� �vFO#R����Y��d_7��6�9peQ\����W+�4M��Um«2�=�8�+�6v�{k�!=����A��ە�m\�#�l::�ť�wue!���#��W��f�:�NJ�,sY�g%�1��ǣڶ��5����aU�TWZuFk �MtK�㼺� �\��ҩ�����k,�&sv��W��(���+����d7킖Ä�l@���d�ǰ��;��p�>3��A���#W�i�~2�n^��R4���^1��9Ո��O�;*$��Y*ttG�.� �׫�(�t��6JWp%����r�:'��sb˗�S;�qn�s�ե`Y5�[�!�c �/nP�q0�#��D����Ư��{?U�pYWK�]��v��ʫ�(>���2�����y��4��&�ԧ� 
�|�eq;|:�χ���w ��
�e�Q�N����-��T��7��={I�6aR]�:u�}��.�`q�D�i�1:.(��Ŷ�PtOt��
�O��������8��K("�S$�wMT�H�I���k��-2e
,1IX_���;�*n�=K����i!��X�;9H	Z�ǘ�t̈́�af�b�Pz	|M�p�@ǋ���=Ec>#+��@�@����|��-����"�l��9h��Ns=G�aut��V��K��6Ngu�cO��峒��� _�)�[
�'���r�_��{B�Hȸp!�= �Ӏ��}B�"2�p� �̟G�k5~�d3��0O�ڔF���=�g6��	�\3�G)�3��ha:};�����0��,;�˪��#��Pa(dVT�C �U�y'��o�z^8E�WG���^J<�0�.�K��Y�5,�D��e>�'P��u'>�mQ7i����z��"��r�I�n#�R����:���>�.��Iճ�4>��m �ze�����]��֪vڶ	_:��%UO-W�j-���I(�O��U���%��#�����z�ƥ����=m?�KȪ䰏�W��&־���)���;�n��-�H!���e�]���R}<S���d�|��X�n2�Xz�BV���tU*b�9���g�w��#���o��D�q�5E����s�1�3�.ʊ�+|�Q�m�+_{�m�kaFBס�Fkx'P<�:?w����l�KJ��)<	�FL��@�^�m��j��� Ҥ����l�0�I z��k|3����-�2�mu2�Zf��1�|0ޚfI�D _yòQ�F,u]��ER>�L���W�.�����j�OK�.�ȚH5�a{��Ь]�|o��@{�b5�p�|�v��� `�ߋy��a /�A��18����"IcCaD�Z׵�l�=9{=��a*t�m���e�L�u������4v�R�#q�4=�y�ǫ0ފb]d���u#�T��g�EHco]\���tN�%tݞ�AVg�y3u|d��(G)�f&̎�d�>� ���z=|(�|����x*������|Nn,��"R�Ga�5�2�~���5
��r�v�����*!���'S�x���m���ʪ/���Ԍ�9M� f����A`�Mk3������x	c��E���c�	5��DW^JG�)ka����������C�*��-�Ú�H|��j��f�72��cT���x��O�H��3CޡS��ڻ1���	�d8�D�����v�r ��F�@͝�����GKz�k��׫\њsUI��?ݑP�F1v�G$�q0��Q`�~I�>�B�u��j���4����93=����rٗ�W�8����a�����8�kZx�F���4p��䢝�M�|�����L��z_��'}4W��zd1G���x:���4Bzie�sPI�0Pz�{�I&�����$�����Aj��-��ǖ]:��MX�	`�*z�Z�  ��~�*�{�P�u_��:����K�)Ǔz�?�K�{LA/��	�Z%s	����ur�	�?Í���]ҩ�����{�7�Z`���c�D�)�-��Q��|'`��K�о�t�.	�G��"�*6�#~2v��s�����cf�nY��Nཝ�E�}S&�"]8�ΐLn���ac1�܍�IP�8�i�
���"�7=!S	�BI{}Hy�f��7�iPn���y9� 0b��~���y�Cx[pf�p�g}�3��>c�Q��y�g��?O��z;A���_N"�O�k���eČn-��?�L�Ui�7�}�tUϰnA�v �}	���Ն3���/H��aĚ�^�=B�sE��r;�S�u+Ӌ���N�Oi����R>%0/\P��]\m:b�	,v\̥j������O:���4�sij��ȡCdn͠���V�E�!�X.��+�U5��0���m<t��S���էIY̤�sQ�	�qo����L����R�9~��v#L��&��GmU��y)�����r�Z����s���8Q]�&��� Pi�O�F+�*>�T��#�Dh¼G*�Ã�G�������E椘��.�`�h��,0�IL��m)�����pV�)͍�{F�H�s
-���sy�qڦ޺�,K��B���>[	6hGP�|;9X�z�i�:�w����=�NڕCx�#���9ͳ}�?���T�ow��n}��N����d�7��T�@��?4��
�=�֮�	W^	�bs�\g!��ε��kn��x���Rq>�\�1����7eV"����ь�xNѣ�M��Qd|PQ5E�l3�/�9�s��L%�*���
��Z&#�BB?Į�x�a��ч�2�k��H�6DY��d���50���Ͻ��T�7ߺ��Ty��sZ�9��]bqO�B����;�� >�q,
��A��~�hE�c��A�~?E5 DXp����!�l(��7���b����A��ވ�Ê"��������$'�b�{�n�3�F�Z΂I�$OLi��h֝�X�GgF7H��wj�0�������1� ���i�߿b6�_Y�$��#� hi��j̫f'c����z��$��[���b��'�$����AX=A�fSB�Z2Y�ĵ�km*q���1>��n��+��\^�Ć}B=��,��E
'���$���
�-/ӽ@s"�m�k��x
n�(O�y��#�y�c��)8�%-�j�&X��A��l."�:��$K~\���S�:�,�g�FT4{�oN,m5�g"�EV�@��6�'�8RFs&����B~⸜��Z�wZ��d+rL�Q��;�U^N'�v��Ь��F����:��J��p,<���ι+��׻ȶ���Ǳ������` �By)0��b��$^�.��1���?#Jf X�S_���-6���kL���1�T_߯��o�8g ��1)��|���ge4���v񳝼ə̀���oe�}g�D\�5�;9�X8{^��7o<�,�ůc:�ݨx)��ɘ%P�o�'�V�l�9�����l/�nI��d�kdX�1&�R�	iBur����~bG�#����ӀY��%=�)R�.�`1 fk�L�,�^$��n������u�i:!��Do8�AF�����md�c��#c��h��oP�gr�1Qq�O3�7NoAb�ݸzu�3�H��͎�⺣�f����q��Ie�:U��R�F*Qh*7�%�JB�e��x �b��#�_�?�߈.��dw��Զ\�$��,R���Ѵ�.�uk�O󥒎��9�h4	֡
.�Ʋ�|���Cֳ�-�z��[��C0踟'�tA�CV����;WԶ�Yɭ�z	��X$%�/E�>��b*O'�t�}c�����v��2�w
��t�. l�;֩	�+�Đ�@©`z�J�8E�u��]2���l]I�c�'n�uоP�[w]O��.����o#~�c6�=��+G�l� �HxF��>�a6#W� ���.i�j�#	�rB��p�*�"K�N��yΧ�z��?-.�%�l�?"���#U�7�F�T"�"S�G[(��mp�IY���mc�@���)���_���Kڻ<�Iy�*g�Yq��}ʅ?����n���{MM�Gh��N���/%�M��=�?����!������o�I~��o�V�#�O�v��ޙ�ׇ�D}�t��q�B�V:����
��gS�����\|�hKV�N��;�nn��� �dH�su?m�z��h�hg�LBd�'�H���:�%C���>��:�/��t��p ,})Y@�x=�'��PW�g�BY���ܽ���=�P��v{� ^�J�5���}ҼZ=�W�K�gP�O��G"����FͲ���G�^���]�)H�0�恆ԱA���W�/*��#�<���D��r�
�j��3i��Nm�bA@m�+(R��$�m�9=�cz%����g 7��c�&[ پ��s�<~9�N!���b�]�$�ޏ��?��T�Ś>Jpa�m�F�����MN��9��w��s4g?�`O�Y��7c �jF�R����T�OKdv�'&�Yߘ9�+�U{dCg�\�t���"�oeIYq�{�.�y�I��T���'k_F�4�����rΫ��<��Fv_��w���4�K���[r�7����\�<�xS4�-��m<���*m>��Ǧ2�S��~/;��h�<����肻���Ѯ���Z�V�V,�b�n�p'N������/�b1P��/#ui�yՉX`�b �|o0�lKZe����sV��Qѱ����v�}�h�`ڨD�UO���eE��WC6m̿��5�a� X)臈�Η�W~�V��?C�m0��#������$&��Qg)���	�_s+s9a��cm�X&���_�C��?d�}��N.��m�T����ڎ'���;���=H���b�
�j}g��7xv-���.��ɬ�>cn�C�v��+ik�I��X3����L<��v��TW�_<�Ԕ��u�l#�49�~@_����k*�M�2�}�a�xA�H<%4�H{��Y���r�#/q�!嵷=�Li�3�5f��q�m�{��Li�f�;!�/��R/49W�fw:N��c��O?JN�V
A�I���Tف.�¾���E�:��8U��	��X�KnfP��%r����#��k�u����a����?�E�f�o��_���_��	�~G�-O�l�	� l=�� �˽���md�,�?�K�������tj�s]j>>���%/�����hU�rO�S���z����H����3��º}�s��M\����D�=�嚮��v��1wR���"i����*J�Яi\�Cj,ʀ��$�;qW����huf���!�)��d9�FO���
�q;�>��Wֽ�c̤ئ'_4�D��RK��
�Q@�Ǎ&�n��j���]�h�7B5�-�w���2�3iJj��~�-�n=���g��7�;�zU&�����eYZZ��ސ��%)ln�-F�;n�6��[:�2"L:���l�з��{J��PpZ�
\�f>���8����żD��)�;Y��tY�g!^���tDv�Ϟ�kO���k���|��4/�^�4b��j&�j ��
���L�m}��F����[g��`<�q�eI�CV�~d�IyYD�RA�H�!�/�S��{�A]o�2�3���)r�ۏ̛ٛ�=�_� �unxl��M�x�
�׎��G	�����gCƊ���|�,�*�x�{SL5-��L^^#��/Ύ� <"�~H������/�*�f��A
�&�.c���s���IdA��e-�sID,��Kp/�y���?�J��i`��_�~{^NvʌĠdZ:���Wl��I��?�~�!�V_�s�\$��y�~��4�uV�pH����Fk�k�w�M�׶J�
Җ}�,�u���C��=���%!6�\ɣ���T�|}փwZl_���!�*����:{q��vvn�M��f�5�O���Y�U���7@yH����I�hi�Ug��7
��$����I@�� �q�U��0�'\xP��i��>h{q�w,�O��a\�r�+Z��	r��f�1�Q�S,���+�Ș�<��I���\�����So6��C���y���h�$�d�h�oC}�X�h�`���=�u{����2���4oxR�=�=����[8�R�n��`���$�4f�B���^3Ap�B^[BQ&M[��Cw[�<��!@e����s��j_������K�*��_�KJuk�A���u����Kde>X���bU<&�`y.u�2����?��13_�qw¦�C�-����I��ٓLQ�������D��<~��4 n��є����|��T�6#)�Bd��$��סu�=�����wHKr�b�c*�(�����iN,�:`5{
���nFG� �,O�38�k��{hЌ���.���_��X�&b������
����9 � �t�˶�i�x,r&A+�JD8���P?-C挖;`	�����k��J��;�J=/t[�݀�z0�+4��s�6{&�p��y;�C��64MQ�jN^'+��L3%�}��ߋ�&~v���!NO��=R/�E ˘c�>m�i�ikúء�}��#G��m�[�xe�ۃB(P�+��҉j�G��m��z��T��L�Z�ధ1L���jzύ%G�jO��[�v����dѭ[�!R�*�ҳ��F�,�{���� #o����t1_v&�O�{�b�"I�m����� s�Ӗ�L�d���e>v$��ɷ���jҀ��eV�wq��8��C��6Y���j��j���F�$l`�c;ZGa��W��x�3�V3'eR�g�3	x�����s�����y���q��ۀ�ؤ��9���e�MK��bg)��턅��(�Kxu]?�����h��m��&QKiS���d#�j�vzL�DD7����Al��N>Ĉ�?��;�uR���$����%A��PK!��ዺ���氇����k��M9�,�����b 2b��?)us�u�]}�)J�{�-G��e(|}�k����IB`�8�F��w��vB�u�,fȢ�-'�]al��9Y*��_P�ʪ�_���1/�g��=/U��[�&}u���(�\C�:Ԡ�h����P?�Ȓ�g�T�'�Yo*�|E�J�)�<��O�X����?�<���3G�j$٭����-Bd�خ��Mo��h}�y�i�l2a;>�<0�/7��֯F�>i���Ά��U���;e\���]İ(�g�c����xjh�ce�.������8�|�3�ԑ>�V���8���V%�� ����6��e�l�����nֲ.W�/$�n�-�:�5����\���փ1C�~�8kZ��wV�Ҽ��N����0}�a<5�^2J���=���f4�*��؏��OR.O�:^�)L���t24@]��}��:�>��گ�A���1��d늙�t�QP�춓��Ms�.uWJ�RJylJa�9�,=��M�F�ũa�����i�&Z�^8�^D�D�YPi�G{��*h��n�[�Z���,w�����W4H��{n���:�ڪӿ�o�H�BVj�cQ]{��h�s7oҽ���V�K�"=VGe�?`i����3�[�K� �Σ�C�}5�,�),#�Y�Z���Fj������K%�y���B-��)h�+ʤ2��ۂxt(�G����Gj~³7�.���[:�>�Q ANq��������������O� ���9|o��X FS�Oi;oK�sҕB��R�Ńaȋ���#�P7����פ~�$�/3��ɕ�Y�>x��Y�R��3�g��3 ���c�Bxة0���'����	T�k6�^��n���t���*<�I"$e��풑VuzO^d.lN�OI����X�2F�L�*w���-S�����	oBG�������.!=�!z����P;H����-��D���a_d���`՞������"��m ��m�y����Ԡ����.��
�3�� �`�O |{Uߍ�;gPw��QR֫��E��#�� �t�:|]��<����1��nB�h�5�k v�[���!x�燑����2!A�G�tun�֟��{pǘ�gץ'��F�G��K'�R/ə?��|��)��Kؑ����Hr�:\�l�1ad'q�ɸZ�������P- ��QY������ǕJ��鈴ǘ.#���Pש�P��Pպ�+�k�D��͚T/���V'x[r�B�䍔�pG��9��x�:���C������5/����AKVdbtv�
�V�M�H���`������мS[�@���>Of�̛1D(�������~������Iq�]�3)}3�w+DV~SqԸ���O`���rm�%`�]�@0h=U�(a �����J�w�!0��^�En廜՞e
���ޟ��~��^��z6R�Q�D���R��ӓjs�a���K߲���6��湒�9��1�B����<2�wK7�����/[�b���8x`�P� k���%`"��>��5C��o����ac��G�aF�De����KΟIY��w{�)!]�pb*\^zo�ϑd0 �����d��7->�����?+��1lW?7��������i[�~����%�¡�p0�Y�ow�j����Џ�.J������RP-�oC�T�[(tv.���B���Z�]���@>��>l�	�A�e��J���Ð	s��ӳ l�d�2��b	?]X6���yU��D ����;dK%iȑ⎱��j�=��5���1M�I��;��'@]���������i6�;P��u*���|���=S@G��w�?�k��h�C����d%��S?s�u�a���$ӯٍZ.n����Z1ǌ����z��$�{j���D%���db�uм�F�������X+�,��ӄ�R�j�KO`p �ܑ����W{q,`AGc����c|��y�{G����dT�DK�@�^��B�5���{�Ԉ���G�H�XWxGv��(� r��c��s�Hn���d.��\41�M��/H��*S�'��/`er���^r�Q�J�L�|6�jA�R0�[qA 1{ؼ-5mýl�"t`)�d$['<��.�u�-�'y)�oNe
��! )�(��N�K�\����JI.ޚԤɧ���AU�ggi][\���8'qV�]w	���q� ��n�R�eϽ�||@�
�7ܜ����		��NW�����Ku���C,1�>�C��Х	��7��NT%|�<�x,��3��oSA��R�/Φ�e>F1&E)r��!q�>�6_��~��Y����9�~�%|wD�:�/oϚ��u�� �i����d���/�O'a�������k�\���_^�w��� wl��,���h�Z$�ל�����E�ȯ6�6�~�L���:'��٪?����ˬ},xF�G��q���/Q���YB����Mد�ev��7��0�x�s��^zDEUm�й��>�����lŲ1�{��T+�H�7'��Y�E9���[eX8(3�)���GHJ.3�U�A�&%�
�hz�<(�Gjژ�|mJt�c����څ��� <����׬`��
J���[1��D[�N�[�_���hb���9�Y ]by��쀆ñ%�^w.N4��_tc�$��N�d��l~�|�b9���~(�ͼ�a�_#�c�4��W����Ȝs�H��܊�r�92;����`������)Fֻ��8�{;������UQ#�@aZ	�w�W�z�D0O���C���ɅA���,�GDt�EH�ג,U�e%;q�Xqus�ϻ9&���Ӛx�����B�<b��/F��R����t�� n��]3S�9�E�׶��
�ĤJQ�<n�G~�KJ}b>�z�)6�3�[��eC��uK&��z��Ȏ�P�en��:�]�{������vE��>'�` �e�u�Qr2{25NKG�܃��MI��$";�J���w5P	��^t���u�ˡ�au���[B�����mL�cȇ�3Be�:	����ɫM���2��"�����V��z��%�b��@|%H͊d�?��}�a�gOh��b�y���y�����h1���o2�̇�~7]۱�KC�� ��Ӑt�� �g-ֽ�x�0gSr0R�$}��V����υ���9%��]�q1�xĖ�(^D�Z��}�
l�L�����t�,6��w�� ��Õ��Y�/7���w�2]����^8b����mޕ�m�ò�JZ�@��[��ev��$ (���w���),��H^��1���� �SN�qݣR�U�h�}T�햣h^J��g,Y�6W�$��4ZO���HH����,�G[A�e)��
`b#���g���6�#R.1�R�OQj�9?���� �L�3���_ޢ���:�o��~���J�_�,��*��^�`�Z&'���_�پ�EX��JV$���K���d@��6?��ʥp��o�B#�����5
%�J���wt[��8�� �V���> ��q�����^�ߕ�}Qi!�Yhg$n^�?�e� �{�C�DZpl?M{}�������-JG�0���pε.���0�*��4�	K��$�K��L��~L�+���IS3��WJFx��لP|]��9�`)�AR`*A��)��N�7�x���+�KHV�,��8�L����<���$�����KIV��?�p+�����'c˾�H�)�n��GRD؋�1]Te���.�tn֝�ϸ��R��-���4�+m�5w���B� �5�B�r�FU59:���~��2���M��E~��]�����Bϓs�ĕ���������>�W��ymԞAS����G��o�{qp��.!��~{��,"��rE�p�0]�p��,h��Bp/6k@۲Eμ:�Q���^���8�!p�DU��XL1�*�'<���f�X:�'^��;V�ʁ���Z�Ka���˳9�Q���|��T�)�������2�Pw.����$K�C�s_	�P��ay��;�h�Yʎ�����(!��)��z���g �˄s����W�V���g$h�6�v�-N,h��<?ٺ6S,yE����9�{�t�FB}��îP���+3+B��LDl�m��ӵ�~�9r�wH8�ř*g�e��Ԏس���ޒ��6/��� "�~�YT�&vu������L��W�M���$a��>�}�G'���{-����j��/ �1=91=��BV�\�H���\m����G�EZ�>�ZE��B�r���.'?�
��L����3J4�pNA��>!�fc¢;�Zr�Ѷ���]�����`<��۰5��k�m�U����Wr�Ke�����(JI��h��VZ�T�Kϒg��3����&�.L ����厹�A	��w�<bنΚq1�@C�$ޫ�Tһ�)}n��T-���@+�ꧥX��)�a��Yj�̵����Wp�/N�������wD��=ܭ�(�$��тS��^��w��8)�o�걥Wu�ͫGF#Ġx�B�W_SmT��ar�"Ǆ�����|�BW[�UF쁛�Ҩ���J#���`����*�`��ޣ�[���|k�g7�!�����Rǉ���qᑦ�L�U�4��7��^��}����1:�����s鍏�E�Ϻ�9��������Ǟ��6�j��m�  �����Gs�6�V�!8�쮇�%&�o���������[�@LRDY��C����Lol����Q��xzw�I%׫D�#xd[��Ї���F{'`~q><��Ʊ#c&�t��s�+��'=r���`���"��P@��0�l�{�+M�)Ko1� 82�h�����Mkw��+Q����rC�_����X0�6cv
B%)�����!��:N�
�3|��7F}g�o(�X�H��r(mz�(���/g�7t�{��9g�ss!��=��ZDjVR�������G��E���=��a�a���B��M�Y�4�����o�֌��/�	ͅ�B�ߏ��k��"՘9Shc ��)�� �z�d8$��Z�(G�x��BD�wR�F�����<"��q��p3����d w	E�kU݈c�L�$������1:#u�5���H��'�{;DP2��&>qYǫ�M��(���2+�bEdi���X���4�w�7+~�g�=w)3��!*/�-�Xy7��-Y��iYHg�{��F+�+�8H��EW��L�؆��X�J�D"��N���/�^�V�0�����0`���_��G�rh}��G9Ŋ�&$�|�pk��ſ'��;3	"�-�%,/c��	���7$�O�x��;I�t����J˔��W0�#P�jne1���p��Q����d$?m�{�Q�(��$�XC�,���"3��k���EJ�>uy�D�BBT��\��-� ��QF����c�W��r�س������4m�vtU��J)�Z;�!E��y�����*tFxxR"�F��=�n�t���o}/�>���s��b���������i6&A�AD\`���[��)xCC��!�e���l�m�{:��@I y�'� F��~~ѼA��(+ޗ�D�?��ٝ��z�٧2���@��Ѷ���:b)�#d&N7���=y@�=,��EG�r���UɊ	���(��&��L�2L���RC�R��xP���wƣ4��{�(oD��M�J��j�p��2��KW�d��6�]g��%��Ep���G��u��7������fzy5{��N�%v4)�$>Q�c���\��,N��ŗk�@��*лc�W{�9���5�IK~O������(@ТqFGЋ/���o}x����/a����B�/9W��x��9�"Y+`f��<Q�HׇԴ�/�5<��>s�ҫ:)�����d�Ѩ�2�{�3�s��B� {j�kkQ:p@r&����8��[�i��!ۚmzх���Hd�#���L���:7xиw����ި�L_�q���x�:�)���<,�	��L�����P
�9�9iY�H��o�+ވΠ�R)j�#�>�OklS!>���rE�~�2�E�� ������QC��g���zV���8����g���k�Ë���^��cѝO�Ӆ�*��w�<�!�=aOO��j�cO�+��Ig���:��l L?�i����ȝ
��Xa����#@}c�R����>.<w7�Hz���z����2v��N�L��3���l���z���T�pE��T|��r	#�?*H�_��⭾��������jP� >POc~A�dp����4i�gV����]����,W���S��G�7#��eރB�Å(b"+�'@6�=bg���;��w�xǵ��d��/k4�CJ隱"A��-� <�sD.EB�P;s���U�h���:8˒���AEcȹ���n;م��uJ�jM�tJĀ�?
�,�ht�çFR�͖��i��ƾ��\�|�x��h�CpH���g�#6b�c&�-WM�&���O0y���3���`1�@z-:A�'�3�����-�-꠶i҆��=Ham�q�<�\6Iwv�^����H���#"s���]h��w�>M9ރ�mϫ0M��7"���!D�U���8��
 DHsyE�2n�@S/�1��X�RD�չ�﷘+G0��v�Q]72d`�m��ƞ;��N���53Nh^�wV4��d��Hzȑ�2%@c�G�C����K >qtF��A�(f+�N��[|PF+�B�Z�qՕ�P����%�A��_�ߏ���4��e�0B:I�(�m��Y9%��2���JJҿ=�O/���o����f�39*����ƾMk�C��f��_��'!��qCf}~�������f��v��i(����'-�P������b��N��k҇��s�{(KP
W�lC P�n.˅�'5'����[.i���R:�����&�Y�p��t0�)���ݮ*�I�A�T|����켶��(Ոt(7v�� ����j���l����i$����(o'aY�3?*`�n�tM--��i�`!a�E�B�J��:���>k 8#�� 
P�F^�e�4 16/zUW
�'Ro5o���H���C�ˢznAe�O������KdG��О���[]�ٵ;�=+Oi�GO=l�D�ƴ�)#[,TA��Y}���:TQ��IR�J���bOb�B�����?��ÔE����U���tLԮ;�/T;�/u�/M��7�m��PU+�C�6���0����
� S}�a,Ӳ�XW�AU'H}�v�-�è=����>5 �|
����\}�I{萼N���7��!<��4�Td,7Ck^���o_�a+-X4d�|}�H�H��A�S��V�L�5��ͨ,��kß
NCY]�=n�[v������o�����l?.@��Ѐ�BйR���nn'%�_�X�Ʊ�L�bԛ���	���-g7m�b�Z��
��b�u��BZO�y�S�
��`4��Ä�fm�(w;B�j�"����b���[V�����K�4�#�-�o���a!�9
���_�Ů�i T!�J�6��7R�'����P��~Jί�\���.A��|�� 0�Vj���L��u�UV�����w��������}���I�g��b�B�|~�' �����=d%�X�-��j$�--��t�*';�Ro�e�Ĭ��n[�n�Lm�o��K�x�e��Ws��wLv�ȿ��xE���5����{V�m��eH�������MK��ҩ�����
��C8ʧhR��:�!��!���U��;�=m��P˧�F��lxOh7�t�F�C4ڶ�<�*����[���޶bVGՔ��oZ����D�ϾC���}cQ���U�J�g��ݸ�/#���m\�u�<p:�ĢǍ�k ���k�n��k����:&���u�j��wq�s�~�@.qxx�V�O��)�ƹ{��B}��!u�ࡈp�t\ǘP�U/��ޮ�5gtl�zx�N�Q���y?�|e־2�3��,�?h4 i�P�l9�]��+�9�`��wE���9�f��B��˫#[�!'M^c�(#�%T��m�!�mk�J� *Om�Pa�i��JЖp�C@,P��KȊ\��,H��X�# <�0�zrӳ;8�Q�z�$n��׺�tO��|8�����Uyp2oفP�h 
�M��b߭��Ek;����DJ���V���Y��$�G%*z��X�f�?�V�m�{eɷ�j.�a���W�q�6J��7�/�Xunf'�� ����_��*x���ި����moT�w�����4�����B&t�E�l��vupxc-=����쥃B�]�����8���}�,����@��V
�9��6�m aj~6bPȈ�8���z_�.��o�!�I3��q�C�'��VU2U�����	��N�X�l�Mss͗�_�n��ܡ��#@�����_�E��P6d@�M��ӛ��a��o<�.��d�G�gq�W%(�q��<�W�P�wk� 3X�a��.����߲r���vk;�V�~�f��Wd6�X�'�0��i����ޜ��}=�v�z�����R�U��O^/
J�>��*�����@��zZ���y�@(����'�Z�CJ�
+��HvG�mpk|�w��W��7=�!�����Sn����n��?g�B)�*G*7Ly�������T�������C�U� ���k�RQ�>��B{c�w��8�F���_��g�'3��g��S�g�]��%+]�o�ºH�,��ZD�Y������=���\�ſ���mR�"+�xД;�� �դ^V�H[�Bmak¸����,/gz�`��ա�4Vm>���	d���k�l=覤Kr���J���B(�rޱ�H12��{x�ԉ�猨_����)#�-�kk���aJ�ı�ë��I���v�);�j��UosQ�(t�H�&^p���P��=vC1�;������,ۺO�0��@�7��V�uv�j�K�0��?JU<��@�g.�%>胊�=�Ŵ�[���ly��9��8 �������w�c���n�8 �p�s*�u�0xj��D��cGU��ޣn.�g+ޔ�@6_`{l��,���'�l����3bȶ��f�������W�gn�4G��ψ#f0�r/�h�_Q	�1�u�phF)\�t'+q���M"������$��7��U7�
u�N>_'=�9hOL�$P�b�4z"�Ź��z��#�o
�����O���$��y������G�Y�s���)-)����PTϬI;J�q�2�;�b?F�9�7����#���-U�����ò�PC�a��\�4��.�l�kw�%3_�"h0S������)��W��u�#W}�εέ�x��R/�n}/�+�aF�'4��ad�V8�YO�x�di!�F	_��/=��Bbel
aP���;5�0�����L�չRI�껌uT�+r��7y����k�)B*L^��ZN�
�{%!N�V�)���=PY���(?м��"w6�h���4'���|׏�m�����ևX�, ���W��%$&�4eg�뜥�
XH�N�\��aRG	�.W�^z�7�\�^M�r`�e|���)48Vt��vG�2U���WYH�φ�:U��BXjj ����@��x����|6�*�q��7iM9�0��JzٟY`���¬�������m������O���U_
�v<V���U�½.`la�-����̚��i2�wN���z���l�u�-#���hՕ���̺��H�ސ�����M��HD��ȼ��P6-_«y�
B��0�ԥ� ����m�@�^�Y�#zA�_N7����Ba�+<9����}�7T��&��σ�v�'.�2���5����g9Clr�ٶ�w�~GeۀCUt�a�7#%Y5f�����p}�jA1���V͛��Xm�|�t�����"s���%�q"Ox���8���D,�v�$[�����[w.sY��vK�h>�����)�4S�Hp�F�a�Z���vrh��%f���$U$%���g[�39հ��ώ*��CR�LZO�5ױA���%�;�bs8q����5K�!Kѷ��g���Q�-�T���tcI\�g��$8�.NF���[��>���z�������$�C���z9;Ax�c�A�,��P۸X33�~��ZP��,�A�e�8x�]K?��;�3c�l����wMlm�8%m�
��T)���L��$R�Ƕ��<�ߐ��B��ꆁ�r���2��>��M�� ����&R�؀}���Չ���y��U��}MBuM�Z:%� �M��'� �lRTX����bO͘+��m�+�k��p�VD�a���>��"p9X���p��3��;)^�����8��(�Y�1��W��[���Z3��^E<�W��A�����Psp���b�s��Po\SHf	�^8�MaJ�@�D�m��x�͙�6C܇Bk����g��0m���@N�.÷��.b���Y�-�'�^N�ص�+M�;C06����.��Y�^p�������0�����p�һ�X]�ܬ�K��^el%�µ���.o�w��˶���JZ���т|�D'������h�d@l"tf�i��Itu��]eL�y�6�j1RC��r�M��y~H����'�E�X2�.U=�>�� �_1�����fjx�\l�	�Kns���)�dDG ��3�i�1��^F��Z�OV��) 䞐�^���r��M ��}�lPN�=��3 P�B�'�*��e,O���ɧ$#�|W�X�/%:���ܸ9�Go�+�V�}�:��l����b����ǟ���MF8��+^}���O��gy��A[�O���=B�\������mh
-�h�u-�xYlH�\���	ec�B��Ƙ�mRR��2ziq�)�p/����C3J�<�?�J�Y��CB�z��n��>(!���m�O ���`v.0���U��w	=b>֘~p��Kq7�|��'7���:����q���,<!$�	1�6]���&F�Y��3�t8y������}����I��m��3��Lp�$5��r4;�b^;�`�W\������l���g���u���q��4���f�K4��z���77��967v���"�F�~�WM� 	���63�-�4'PiNrq�ݤ_0׃dY�f!�0J��m"x 5
�M0t��?��L�3R�7﵇��f+�-&�#v �7�3Hy�y��[*Wݢ%AjW�m��"��s����_.��`��)e.^ymC9<E�S���"�[?�I]���hBБ�ܱQdĤ�8�����Z'G� 3�C���DA���i:Sp@�����+o���e�Ϲ��Je�CI�s�,MƄ��ݦT_/��mr�MR�
�2[T9BA�L PB^i*�����h�X�����D ��V��qS��wbC*�@��-���hE���+��Sk� g����0��l���\ʍ�,I]�����u�9�w���H���]�,p,�w�� 3�c���?hCǚɘ�;����29�D �`=�HZ�<ܿ�A�#�A�>�W_���=y��Ѿ���� �d�;�A�jz��wgeU4��Е�e!(���-���\$�r��z��7!�u�}9������~^���_��P��J�"����h����9AI�ħ�	O��醖�xJ�Y���%���^CL5��[8��t�o���5=dK�z ���m�97�A���~�t�cm4�e�n� E#���_�7k]`gfo~?e��>�
�X-+@nE`�`)ד�æjQ~]J'������K�,=J~����9�$�Y�[�� /�������0Ny��(e�g��K��e�S��O��E��2�VM�������B&��F P�tD�S�;�qIU��o���j�]�l�Ka���w�
0Cs�M�jJF�0V�=І��׮{=J�4q�Q�R�>C�9��:�gir�lxk��EB�%.����A���,DL!��\)����~v�����ww�K����z-�@U�"�]�~�	.��&!Ԋ^lO��h��2&
i��WH� �w�o��6�oUr��y�f��Ib��k/���#������j�3�[�V���)Q��|��� �5$�,Lm�=�3O�H#���	-]ʎ����}�V��́y��;���@L�SS�y�m"A��`0��������#eja��|<�V5�!�����4Bw���W��K�=���tY?ɞ������G5�;x��c$��?��Ń@3u�jt��Z�.h:�3E���M��42$�t ug�������L{.��66��}:|��SE��ae��a,���4�~ �c��ݯ���7�f���n�"1��2.%ς��KU�q�cT�v5�9���2H4K���� �+���1�����+>�k%b�]E�S������A����}r��7��Ek��Pm�����l0ǲ�Z�Z;�b�p��K��Ț�tSC�v��j<Jܵ�!���L�\��B`��]@���.�v�\n&�-�8��e� ��%���]���Dupx���R�Л�i,��&�)w���0Z��g��E�h����Y��;�M�RX�J�-Μ`��*�}�^(ak�b!�UlsG�Q��,d3$�d���>���D��0J��N������s�#���>���,�VЎ�>��h?��.�����w����� ���s�LA��.�J����۵F���`@/�11��*�aT������ ���/�m��I^mN>�lۏ)�r���3�h���Ƥ욶\f�(J8���K���.'X�D��A�e��ğ�NA�TV�̈���*b)�Z��D�Lǒ&���T1�wARd��|\���֘��iH�xѷ09��EÃ�%򉁛Ԁ��W��']�{��f"3���nΦ�nTu(���cn+�栶1y+D��
�O��4�\Mzc�I����FVb�j9Ď�p�(��*��by��^����jۣ6�ؚm7�v.ABt��q�o:�����Zѥ� ��,>4i)]���"L,p�S�.�A�n�*���+�����;䛰}�ÄM�kWQ�С����Ć7$��Dj3�?j�dR�F,� |6����0:��c<a^���.� Pd���&��OW+f�����y��K���ל�]4$E1~m�j�/��"`���)���m��1�N��7����13s���Z���*����ë�e�8�yo�&~�+q'���-�L�78�l�8�����0���>u�%fI���Gs�@G�j<K���5>f��SJ�rt8|����JpF�n����"@Y�1ȫ���q�[�r(_��3oE�iZ���Z9�1hR�8�l1�2� �܊�BiR�5r�z�z&��4������-��E���6Ո�I)	u#�[��j2�s�9��s��VZ����{����Q9��[��ta#��BR�Xt)p�X��J;fL�ͼ%���0 �[�e�R=�S�7�������JO���ꙆlǢ���	u]���"�i�{��
���n-�|����΍&��QU�%���ͦg�Q��γ��@�W"O��]����wU�_��_�|~ȷ�Ș�	�}��I���|���a"8�����	���]�ׅ>]���������WP���^C�@���T���e��tg�1���lP�r��z�آ��w��89XoH�(��C�K��J�2��65&��ņ�|#�v.��]�I�=�%ϵ�Pa�W�]>�F��õ���Q��IY�I��O�+��ށs�IEb�縴Q�����G,�E?�e{�ߚ�'�Ą���f�H'�ˎ�0��5�]��\7�ɖ`I�5G��`%;�j��V1,W����9Ijhqk�[~uV� <`W`ugMG�|󉣕��:��I41[9141�=�����%�h>넟��m�N����[V�-���h���j6�ܾ�(��/~�=������$f�y4�/���LɃ����ny�q(�JQ�s�����B��(F3�H͐�[�Ѡ*#E\�MU�J�f�1c����4��l��?�i�%�F~�2����f���a�Mx�.-x?��KM5 �4�>� ?ݖ�Z7�s�B�Z��<x��Pe����4������*P���W�.R�e{�xl�K]������댾�g@�ieNj���ouw�Y!�E���+m���J4H�J�y���W^��ؠ~]��( �s2J��-��/_��U� S]��h;�I���`zA�="���%5*��n��V���w���ib��i+��E��.7C^a�HS�_��}h�����b�#3���2ء�n�$Qa�{v>��E�̼ɮ���_/]��B�?�����S��X��@ �=��B���q�O�)ɝƷ]
��� 2�bZf�l�\4�{9�Lk^e��͙� �b59�(�4*ds�Q�W'����EEc��KYNG��upǲ�P�o&!Q�$'*�8t)M�A��H6O�d�T��)�	��Si�l0�)���K�+%�|�7ʹ�Xz�Kx�î�4�Ta)%6�Yq�`���.c�p[O?8GR����n��3�*��t'٩X/9�p}��'p�1�Y܏L��gH�J��0)�{�3�!F!���w��a�,���k������^zj'�{���j�Pxs�SDG���J�N'&'��<�bv	���d�?��G��S���Lʣ�F��݂��AM�d҈�:�*�1�#)?8���ݝ�.��&���$h|�7N�=2 ������>�-?t8O\���u0�����`S<�a�k���j��LZ��0ђ(���뇚Qe \�vd�瀉�:�A*}�C�W�����ɥ�7+�Sȱ�CT$cf��*�"~])}��#�s.%zT�?�Y2�� o�_f�l\Z���Jd��E�U��l�$W���y@Xo֜iX�W��vy0��fb�eN�3H�g�c`p��F,�x�x�ɷH��J}��웴0f�P�}�~`�!Vn�ا���:�ex���},V�<���=%`"½!Y>����"�7`�E��?nb!�˗��,ߝ���딻��7���f�"ė<����h
d����ˍ�>/�J!��I��M����֍n��$[uо���j^�T��5Zv��i��OV$���镞��v�a=c�4T%���3�@�C�n�ϔ,6��.���?>}� ƞ7IVВ��A�|�����/q���̪y
�m.!n:eY{��d<�2���Ε�%�ZU3�;��K�mz7⥎*���܇He�Ȫ���4lb�xc�m�7�����0��=��:��`�����O�Ԑ�H܍�Ɣ$hq骳{>�x�c�"�p������=`-
M��@1l��i�U�̪#���W��ʅI�(D

h�\~o�Zr-Gá)u��0�c=MƲiH
�XQ���E�99�֠����a���� N��|^YBB�p��m2�Э�?G��w���vBW#�0zƄ� �����z���Dv��_S��녖��1�(�6��f0�,� 2���`;�~�n�g�֧>�bJUR��:hAB�4�Z	���,|��b.fl�ܗ��ꊪ���,�l;��z(�eF�}7lH�XBI��W�^n�s�>l��ʨy9E��QO ���mI���6��g@�J��:���{ٗ^��=��d���l���IFb�9z�!�14:�>�Z�n��V���s��].�/D�P�]�x= �0؟s.�A�+l��|� b�1|Ծ��T�0t "T�xH̔�������	��i��e�g�Z�
��)%)M �N0S��C	].T2��.�2�M�& 8�)�8��ٰ��;����9�w��!��r3�<S#N�ױV������^ /h~(�ȝ��];	Q�&���ǜ�V���wI�n�60{����iY�JtIO�wK��e�oV٢xE�\���e,ǧ��&B���'m�V��ѶS��`A�dӬ^�si���~�[!�;§��i��(�6k�������� �J`�k�8��	�-�jaha^���(J�:n��Q��ʔ�T0orb��$|b\�[���ʰ�%q���d��/F�ݾ��ۙ��saB�>iX]�'gȊ=���+����y�$K��'A�j߅�����%��m�Xql��3�/��}M��YQ�lХBR�M?$ۯAm��1�%~�U�{�~�Q8%Șs�g`��	zW�hg魜"R7a�#���dY��U�� �3
A<�Y�ɺ�9��K�����hINϥ���=+*�J��V2H��׽�v4�Ǖq6MlsN�Ȑz��va�&[S�>��%<ctc?w��9��@�b���7���p�b+g)��FO7 �g5�i��2I���h"hxJ��ܡ�h
Uf!��g��7?��a'��u�<>[}�J^�ݨ}��A
~��X
6h�>���?��o����x�n��e]|��n<���lޟ�U����ǜ>���Zܨ~@#jG>��!ļ��}�����r��ϼ��m���1ϼ�����'m�RD���/W|��TJ)}�:\3O��\j���/�I9������Yh���c�O�O8 sE,�0̸t� �3f}���;)fWu��4Q{�I�}��U�#�橲���FLQ�z��^?�<� a��C�Ɗ���7҃Y|�B<�����Lڛ�v)�Z7�P��'74�6�-2�hqǞٳ	�Lِ�(ɠ`N̈�H���z"������%�R-��/��h��d|�Z���J�ݻeM��O�����l����ޮ^�u��44�F�.ڐ}o}����a��K%��z ��	�1<�zs���D������)"{��R����^�$)�J�!�\ӧ���&�X`lz"c/sC���ū<GS�3���������[��<����(|�8M����u@؂j�j�JZ=��mG뎉e �X^�R3��G�`m���5둰O��h3��P �ɉ6���A�M}	�M���9"	������q�!l���*>s~p�\�����~�^����l�s������Ͳ����%�;�]��ƾ��p)t��͉D�u�����'���]�/<|��q�֥"�<�3�ɥ����F��\�a�%�@n3���.��#��r_��/m��n�|Y`�p��m$B;
W"����I��LH,�v�i�(> 9�,8*�Ľ��ha���o�~��i��o�Q���M��5�,e�*��l��v�z\+g7�g���N
���pQ�^ XV�	�b�E�9Pv:�;M�˴Dh��~�-�﷝!�a�hΘ���Nz�n�r\OF+Ľk��cucr�8zhsnߠ�C�sm�g@ ���,��#������X���
4�7m��g8)צP2:�)� 0�g���	�D{�8ra���>-���+Q�?&A.��3���k��'�VMǇ�U^5B��-ax���1��{8�j��o5����1�y/���F�A
zbO(��x�*Zf���4o����ttbW�s�!A���jM�h�&xxG�@8��Mi`'���x������O�Ԭ�_5Ah���+�3�:K� �;�Jp��=	U7�+�O<�w
��@j8yܱ�v�w3�w�j��H�Ǉ��+�Jy��鮈��-�{�*�vph�H��$�*>V����#���u=�B�1�;Q�@GK�@(���a�R�o�V>��9Y�o��,~[�`�b��.\h gC�iH:���k��$3�`A�� �/p��Eu���b�L�J�x+���,EN|�i$3�v=9"�L�ib=Q�$��s��<D�0O����H���6N&�<�o�2lR�b�~x�x{s��v��m;9�C@����t��8����N/2�}�������Aj��z���k?<��J�-�u�	������p�/J��+O
[d@��A{E��'<���ʞ��3J�tsrV�-����{c%@@�yg�^n=��Ѡ��'O�Ry�w�4��+���qD��$���t";�����r�W�~����p�oт�����[*Ak|#pM�6OUL������W��Y�,�h��NZ��>������G��6����w5����F	�
�M��J�&�'��^���Q<��_o��WJ�� rX�Ru�� 2[��umۂ�8oW~tw�efY�С�)�n���D�FPס��CD[�S������#=�]��1"f�a&A�R���K��`e�����9?ʴ�a׊�UF��;�,/1�Wh�� ��Y;r$��F@�g�*�����PΛ��[���J:ꭶ4ZzϦ�U\�]��/?�7�2�Zd�o�:��dur����!g}d�F��R3bd#9L���!�j�~��9K�D���L�Ț�!��nUS�ފ�=:̎Μ�qR��u�vHb��!���ڥ#[e<U�׎!Ο��臣q^b
ݦM]Ϡڸ��ʺ�R�'��Mۇ��R�?J����_��~W=w�St������wa��.���!|���~u�����U�6���)d���T��>z-;1�d��/]jC��2X�"��+n<���Y���"V�2��e�1��(i�����>A,w)q�}�.T�F\1��g�xtT\��Mf�7 ��вH��?�|ʡj
u����ا	����S_
?��!9�"�~9�����k�z�]�\ �Ul�m>� �r|�d�*�Y,�h��9��^����>kQ�aV�|��o�c���I�y��3���+���S%��v��6*�CW�S����b�G6IDH��na�
A�B��Öϝ!������a�
���z�s"�\�[$��,5��R��p��[�Q]��F|Y����Q�*::2h2�/�_�p���o�T� �/�%LFQ�k�nW!At6S�v*� ���D�4���=��I?�
Ű|�4�F��WD�#;���3��5Hj�A�w�R����.�H��l�pTؼm��Վ����P�`�K����x3��������t�ݶ��8�>�m�SF�R����@�؝z������s�;�^띇؊%��"�ޢ[v�n*��e%�R�)����KiAj㝈]	�*���IE��������+		}��4A�8�p�#]Ħ��W���.������HG~��'��R�-|�GsN�U��A�n���v���20�1I5��T/3���Z{o��S�D�KP�[��>ʧc�����������ć¬k����+�|B�"�r�x�ܳ팘��vh�3����Z�g�fCs��Cݚ�u������x��ieC�Y@]uX���E�c깲����4^'�mxK���3�a��ld=#��N=�!=���6�����{Ay���zt)�x�` c�W�����a��53B%�\�f#��W2��Q�����a4�{"`���^x���4!m�FaAf�Ê��1�T3"�����~B|�u��~���r�ǒ<�!��[�t:��|�-u�鐔�ޱ�ē[����ᾜ�;{l��<�"|�e�yT�ΦM�e�+�i�⒏�Ѕs�n����f����v�4���?�`�k^*qʨ��)��	��I,^�k��Ih��8Q���i��C�=͐����W������8����T�"``fn��;$���R�ƑC��!�l���RU����qs���`� �E��UC�X����sǚ�t|�/m�='lcA`�����?_���(�&�Y�R,'�yA��T5���pӔ]�m`L܌�.�	o�[ٍ���	�9Kk����Y�OZd�^�1?h{#�>�tP�+g�<�H6�>w
��<G��Kd@@�D9���(�3Տ5'7Bu��$���Xmup�x]?w��R:iG��f���輷�>j�������9�#�&��Fn(�eO%A AN���_�I�Q����-�@��ory}k`m1V��t�o���L`؜��v��/7r��FCp�����'�{[rw'�����xrOg�U@P4L@��c1Z' 8(�=���0�I�n��=�|N�1��]��p�nY��~r7���I3����[���`�}�yuu�LN�x&��ſ|k�Q�G���Y��1Am3ҭ��O3��}ɜl�ܣIQH|���$��HR�k�Od���э����v8��!Q��V�?J�l����0�ؚE�v*���>7t��Be�6��:�P���nA�1��)�������||*��?c�O�x�s|W�\C���*@G�_%~|[�uX8iw����<!5�����}�H���,,V$6�5L��R"^����h��;zِ�5��x���@h5�K6��N�_3{zmB�$�[��9��}�g�S>:�Jxqy��\�b�˔;ȳ�xOܣ�[��k�Ѡ�5 ���Rl�fV��<��7%26l�֢ 	�'O��dM���p5k����NLMw��E�����24�j{�uͲ���v�Gͷ�[r܂�<�n��P����m͗�y���hI���;�&���2to.��siӉ5����վe�o�k͐C�k��O���)���L�hכ! ��v��:��ʈζ��#\�C�Xa�Z>�S�0�+��R��X=��!��w���$�w�@b�FA�7n��UD�N���3��Ny����
����-�r��wsޠ�^B�~SL��b�5���B|ə�`�<*�.���o�~��T6�>!M2F�7M5#���	s���B�K��������/��_��m��;�Q�
��x|���|׭��q��3�"_��X(8'Z����ݦ�`'ٿ���p\Y��`���,�-�����6`8Xz�n�KǕ+�;�M���eͳ[�0�,NNd<��Z�%ϒB���?�3&
�����)��ݣi���R�>��e$��n%�pE���%���j�X!��vJ��R7!�r{����mR��CJ�2_�v|�v�0b	.�*�|�M��aM����J|�}���Z��c��H|<���o������r��
�oې���B�3S[���$TF������G�%͝N�:�W�}Z�G@�3�dטY�i�W:f���� k��U�Ƭ<����JH��� ��+�;8�*��F@�U�s��R���4g����������L��2�y���#�1�PC���p��[�	ޫ��"��$_<e��ؓ�i�xg�k��c"�uHM�Pu?�W�P�GM���V�>�\sd�PI
���R�RO`��"΃�L�>�����H�$��$��k��#��{$�E~+������"
z��a������1k���+��T����ƪ���=�3fzY���+�N,�JV�Xd|���u�q���s�j�E����* �}n�o�F��x0[0�����4T�1��B�cn��mL!�����(c� W1�F�a�8�w�8@�Js�I�>�0g�M�l�!4�]K�6=����p��� ~"��m�DNt���Ew������\���=.���R& �Ӿ�SY�޸��dA�ZSWL�¹@�C|G�D[ݜ����d�FwX�ϸ��m���g�^h����dQ��S*�- 8E�&�o$x�v�i~9���K�BUQ)�ԐM%8sùl쒏{%��Q~=[#k�{Pʶw��K:�E'`j�Ԟ�/m��� �r+� ���4������*��U�h���%2z���x��c�X�g��3b0�� �������n�!���=D0P�݌��UBW_ڳ�kr,xw���d���^�}�	�� 9pn"?M�8Yp���:����<rB�����&�1�iJ �Cq���ox�@�yB��=b�9�j��|AW����g5�����;�j��`TJTt�o�����~���`.6�d=���R	�����r�2���O���m,�`�	��جl���NJ�Q�uWUF��XT��Gx2pz�7�֙<��[�P���v���aD5hZ�[�R�����`yN��c5�)z�:m�Ф�*Ry"i<B��?TTK�i~�Z`0�~A&�C��i��f[m5%y�����j�.U��b香�y�e����b��F/�V���r�ǐE���w SQ',��c�e�-� ѝ��zB\ܸk\��aa���9.��oĕ��怒��M*)�J~�j��8t��t=��ɓ�K�J�h������H���RY��lz�V?a�%�jk�x!Zخո�+����
���؋�\4���0����$g�����˵l��5��[l��,w��(�h[�y-�.w���g�p]���ut��yy0[1�^�/���h`ݕ[?���p��؝_��;ᾯ�
ϲC�l�y����X8k�_�H��*�9^���q�?�0tC/�2\��ٶ�	lA8�ɇ3A�8ڼ%�dC ���׮����2]���8�
��3
��v�CX��\�f�P�JgF;��J3CPU|��UC�$6�'�O�Ho��#�m�ns{{v0&r#�Q,�e�+lW+J�?G�^���A�7{���T$�Fjo:-���Pf�Ԩ�- ��D��������}<vJ|�.q����F� bw�1�-��g$�;��kTX��V��{#�/B�w����N��c� ��+�J��v�}]o�RG�o��즥��i�<���T���4�@�1Qqt���].)��B�\��U:�~��o�z��`���uS+���iw��4����y��l�JX���{[�K�`k�e�\�ˡ횮����k�t�������E��7E��-������#bG\�Үel����u�,u�U���̠�ǒo%R	��n0��}ʅ��/���˝7M����~��tRO�zF}����2�	~��8٪)�D%�����q,�������Uો�<l��ݵܺu�&�9V9� �uD!m�f�����q�Fqѩ�7,���}x�o��#f'3q�A-�,�ćX���!�o���c�J��WzȊMFH����\$q%B3]�,�s��K�a�.�7����.��HW	[ʩ�h�`�5T�-����謕1h�Z�_uwx5=��E�� ��(��y���i��m��#HWPao�(����U~vz(�����^�(7�ӗճ�/��R�5zu9��`/�N<�K��O �+,�>,�_��Kkos��Y
'�Sǥ����!�x@a����
@c�3��urJɝO-�
$B*��#� �X�i6��!w�����m��i�� �������r��D�7�J�����~IH�`lO۟&�Y
��<�'�)�W����yr�E� E��پp���K������(2�9/����K ��f�;8$�kM/k\ �l������/�E����3r-y�G �1ě~>�I�� �!��A>Vd���"w�-⧿���Y�0#�x��w����X^���4����Jb�ȷК�{��m�	B����
u�,��<�m�Ĺ\�J+���ʴHs�Ӹ.^�x���Q�{.5wsN�6�5���,]ށ@!i�1�̡S0��/	�6f����� A	���(3aԦ��XqbҌ�B���_!���ƙ�L�f�^���N�NB�_An&�&~O�h���ݱ��h..v3�	�g�#�/(e�&�p�j�Ѹ;�g����@{	W ��� 1^�t�߉��X�$�ګ_���_j���������%�N�	��:����8��a����$ͪ��&�d������n�)��w�'�a�b�x����=@I�R���@��٩���F�Y�~�C�q��y]ȵ6�Gg�d���1���: ��3�o ��辤��y
�UQ��*y$��p+w9K�iÙ�������I
6�P  刕Wq�9�OY�ᠭ��q$Y�z�D��-��,d7���_�G��Ҷ���C�Ͽ�����N�)za� [�J��K$N�O���/A��e#��En��\U�jsTx@�k&V�.p%y.��|���Z!�;pS�TXd���qͫk-fH����C�����NO�ڙTY�u�*
�i�r��c��L���9���*���^�G;\�m��?��Q��8UX�W��(�/Q�r@U�Ps�RY��B�[��ݹU�-�I�Ѝ�B+�Ӱ������(
�I2�=�K��o�-Hr�m���~N!���g�w�Abko�M�I�̳��~�Ǻ=V:=� �&t./��%]���J���1@���Q���$@���Ǻ�R���F�qu���]R�.�3�}�s���.�jrL�0>֥�*��R�4�o�𶩞wG7�e�HD1`O�&��ܗw�tC����Bq�j8V���{�D�4�jM��4��U���0A���a�rG�g��~ڠ�i�X/��[��u3i�m�=G��M)����ZM�-�2-�Ě(���7���Ͻ���:de�Z����^C�R� ��B2�A�Y�]�TC�{��V�.����D4��B���4d'Y+L!Ftg�
q���Ҥ,^��u�%��N��J��{$W�yΤ��d?�ں[@((��L����^x�,D}P��H@�j18[�C�3]^�v��R�J�?�J��Q��nv��6կe�>l�1z�r��CNm��%�㟕JE������Hb�{XnS�Bj��=s2[�}Z���1�����p�x�	iO~}���B��N��S�`�Q`-ϮC�׾���]��p�o%Ru�{�]���"b%�OkQ?�IXN��Dp�9�v�Bl�=ì3pߊ��h�	�k�ͦ!(TS�C��"1��Ӌ�j�pw�"#m���S<!4����Uaꩧ�=���v(2ˤ�FzEE�g�$ޱ���_��	�N�cŁ|�l#6�f���r��	a����^т�!��p�W0��y�j�i@'  ϳ���0�FD���:�����A=K� ö:c3�ج���œ�5��2���<����l�&9�&$CzI���J!{ 5�x$�G��۳k�^��( S��յFD`�����s�g���i�#��^7��oZ�����b�D=�U}�♳�����0�W�L]�CǢz��.�.�.������KQ1j��� #W��gx����ٖ���N����1������s��T�V��Б!�S��� EV`C��>_�8����}]$�M4��%�%#���.D��чс��m6/�Iu������ .<�Q��ɔ��C��f����ǴS��	���]ᒠՉ�����cδ������Ѥ�ŝĨwn>��fY��"#�A�V����Gr2}����"���	OJ�x�� ���<��s�r�]~V�:nk"�'�D[��7�O�N�R�������Y�S(�^d�$��L/���y}�:�e)Ln1�^f^�X��^$�`��&7�;�p�ׂV�$ bG�w���Qs�t��:UA�5�� Z������ɿ�2*N�G���j����@ch� t����-QƝk�k7eP]��@�$E�^'�c��w�Ixl��I���Ď0�B�������At���/�mߛ�z��bc3gz.5n;o���#������k�3�콹�t&������Bc ����U�����ٶ�����}�P
��0jc�M�Ӷ"e>ªsb3�l#w��IT!���z���|\�/�����e�\�t�7r��P���0e�F'����C�^��X��	n[��v�of��9��z�ۤ�bh`S���L�]Q9l����չ�̤�&�_H)"��ٷö�,K>��p|4��)@�z� ��""sE����Y�C�f�n�Y��:���%H��RIPӊ"���=i��|�}D�⋡��U6�;����)cSvg�&���C�O*Co�p����#�����}��x�?�/��ZxI������#��x�/{�����X����i?Ê+M�T�����9\��!��/���'R��<�A����sP�>E��n�P����ݺ�߷��gO����m}؁��=��^�k�߼)���&~n�#�q�l�Zb[/0H�w��z�� ���m�|X�t�!|v���~iu�s:��)go�;1VD�ԋui��Q6��HS{�;�F;*
�\������n���ղ�S���E�Т��~b�I�Ifm	�|�.��(:�#X��1����0�1����ܼÙ^˯8��jU�^�W�ؙ&F�5G=r3�i��u�3v�Oĥ�_�oUr��8)�0-Db��?�M#��r�8	I�Q����R�~��`��虿�dK>�|�!�\Ǽ�����m�g'^m����´�2	lv{��X�L�Oq���ۃg��L�Hι��vL !m$=���9a(�UK�+�����T���K�����,�nσ��N�`g�h�5Bf�'���s�����{T���ʜ{9v�i�7B8�_UK�a�6�\7,m�F�oC��Q�8r�n·���ز��כ=�M-V��[��=�}��"���E��,a)t)�Cog>�|kd	'4��t�X�gk>��4_!�����6��CK��VX�idY��28Z)bd;�v݅��t�ń�	-t9S�PՓ;I7���~��U�����m债�^D�,p��j-�l�����3Nu�i��B�"SM.���Z�-T��}m
�鄹d��kܺ2V�u�%�ߗ��a���p���V>[����Og��X��s�\K�����]Lx�E�ZR�������������˥�,.��5k��$D��v�N�g/)adOl-`G�.5�G̉F����)��37+�fH�f�*���C[qK����{u"IIƽ?Bm��fx^��K-L���#�[y�r�S�3j��ꐏ���R�ŵf�9	��z��k�m(�	&
�����Q1����;$���K�	H���adp��>�sG�oN��A�σ+V�x�)�i��񍐑,�LB+���[nͯ���6�w�i��C�]�.c~� Q3�����Vj%�tk�d�YaG�q��c �=��N�кcQ�箔K��{1ހ{��m��$3�2��j� jI�F]x0Z�e��>���1 ��Y0C1��H��;� 6�]�5�pT��,9���XA�o`a)�9ۋ5}�r�i�j��v���??�7�3�;�1F_[+��n(`�6�w
q��b�q\0n�R��3_H%��a.�����}MQ�9��Fw�G(r�@��-W-E����x�)�Z��)��~m��� �%���fB��cË��5�B���M�N��D��=ms�Q?&A�Җ�~��z+��0O"����{�W���֣���ތ�Y3U�K�T��C.?�r�Ii�f�-@ `�^�w��/�=��.*RMWB/S��Kw����Z�~#��(|�a�p4QUZ��#�N�zNSt`<�I�y�u���Z�#w? $v:ME��|���B�#��M`]�M;��Վo��;��wvC0�TE�6ZG��] �<1^Ə�z����t��H��|��u���GSU���>�T��I��xp.�b]QmS`�H��¤�\V���#v�Oy2S? �=,P�>�jf��e��Wrt��y�c��A��U5x�zK��p���x�k���^"�7o\��E�`�s�&$9�|��Q���To٧;��dz	َ;í������S�ĳ1��ׇ���j�xGH����`|Vf�H0W�N|��s���]#[N`���-�ԅu/A��;b�:�XU�%`���BCWx�9j���1�#G[4F�
��k�t���fk	c�wE�R�K��'���p
)�S�g.��WЭ����dS9,?va��fp������H`͒�~
̓���o�u@Y#N��k6�*��ȳ����#ju�Md�ٓ��@����Q��#���3Nho�^T6C�H	��i��@�C���٨��q����e`�xޒ��-���5�����P�0���"�_���MP��)�O~@�R5)�w"i�ي�n�I�(��ԁ`�w��މby�M�d��"ձ�JW;�_���Z�N�P��r���h��;���u�|6��ߐv|3Xf8_3�u��*���n�S��v��6\��LQ�����7eFp�OVIto�9iȘoei���֋�o��N�Zx�@�-n	f�2�V��ޔ���0����}�i{%����n��u�R�c�$�d��p)<�_�'Sm����&.j�J���{M����MsV!ɝ+������ �x@�!���K��6Ԗk
�0�БJ�Q��P�8���_�o�G�f��H��R��@��,iOP�u>�.�XL�3���u��A���Tj9���R9�'�m%Ӝ3�5H�>o��Y��T��D�=�Y��i&:�x�[ت܉�J��4���ss(�~����r�y��0���������,)В���]걗��c�zg�XlB�$��sd�Z*�.P՛&�iU��0#r y#+܇�T��d��v�/�u�$OM��y="S�C��%�ncR�;���l2x^�"(+�T*�Mn��(S� �a4[#�+k��]�V��1u�E�b=Z�bP�ܲ3��M�ۥ�W6�T\���6�d���ɛA�[�W*����{j������b�d���}������n],��S����Wm����$�8'�Uh�� [���K�Ԅ�97G��@��&.�Q����	0��,Z�{�9��p�B2C$ y�����62�Gm;�����@"͐�nD���Te�P>U�#��j��""k�B��*��%/�a����N8��/ڇ��j��(��w\��t 5�%�O�<cl�۔R��v���<���`�6�d��3���|0���w���f��.:�]E(C���S ��Q�#G��X�MA��a��r��<)�?��-ƵݿIg�
GPjΦ_֑���{U�-@~ gi�	�r���������^�|�Qsn��E��"��Am����Fhᓢ,5��8t@���牄�l0��შ�Ա[f�o^Py�"�E�|5���2�
��eb�{e�̾������v��Py�'D8n��2|�B
����)�+�~XN5�w�Mpm���hĐ��u��G�"�AVF���7��i�-��ɯ��*ؒK@w�#�pA��N��S�G�A_M'6�5܄��N���pI�r�C��d����]�G���<�V�UZ���r���h�ڥ�
M��	��Bڲiϋ�J�3�ǔV r�k�Ww9��AuU^A*&D�L0U��_�^� ]ҙ�`�ݣ�0�x���D�E;�d�إ��b4�I��Ҋ���,K� b��;�5�	��ǒ��0��gJ�6+�la�����"2e�n]�s�F��t�M)�� I8��Aw@�u��U�Wը�sϴy��l���!�p`H�-w������$f[j�{��"<�VdF��|U$ɘ� G��ܞ@��d(Uu.Rt`5'��0�����pMg9�=uu=�x�	��0��`�.ڲz�OC�~fQ$Ө����-����p�>H��4�5B���(4���v�.R4!e�ƒ24%3�]Qhf&�L}�TMl�N�謓눾�F�秢qѝ;�t��2 ���/%&�dW��Eȯ���&r����:�]��䇀���п�����~��{�j�M�@����;�mVD,?&������XdG�w���_l�`]P���mJk�[h&��v#b�֥ȼ���+�܉�-�H���nu�q���T��0Ĩ�%�׍��:*��G�����O����hB1���(�THkq��Q�N���[�ٞ�'�g�߮�ZZ8�UE�\c�V�ݵ�<������-<-ɱ��k˶,�ik/C5[�k�>�$-��죀�P�ο<8�����F���±+��#ǼZ����g��Ƕ���z{M�di9.��M�_�m��*�5k"�c��]�
,_��M�F�Uq&��7H�n��G��>Yd�m+�>�;�K�̄�	�@ا���,L����'�na}K���sP*�_����C84Y}qU[5�V�J>��r�����>�-�\�C=t�@��!��V�݉\��߆�e�t�|Y� ��xjϛ��P�G�قL��k��5�t�tW�C�Jja�յ�QLg���aZ!�����"�U�(�0 ����^�q��g��_�w�́�vT��4�'�3�~���r�PP!���-�!�1ȵ`���j�n��7-�J�����Fa�w�X��ȇ��K��	��jV@�S�*۠���i�-?�P ��9��.���0��{��u�m��R�����zߧ���@�Q�4tݵO��ǵ�{�6����8,"�0�Yp�}��Iv̕h�-��������O�G��k�3:ㆥr����i�.��#>[ ���Ϊ����F�K?m,�G5�g&7l)&���JㇻFk�<D�%�B���千!�:�FƾNk�{���1�`�ڣ��S#���=+��̷&¬��*�˂�Ь�{���!���n�>��LDZ6K�����g�/6�6 �3+R���$i�<q?͌v�O;|༃�A�O��	�+�n��e�N AK���=��2�Ӓ�\	ϰ�:��(@[9�M����M���C�V�\�)q-���5Z1����<%��
pZ�G.���q�W�x�[�$�d�A~������M>��0��	m�akg$���ɬ�U�������}��[cì��s�!�4b�%�N��&�����d49���գb���q���ud��f�9@� �N_D�'����zw�_qIFʠ)	!-��5�ѣ�Q��T�Q6l��W�\ʨ����y-��Ub��Q��#�6]bi/�E	
����N�"��k�$c)���G��@�H���=)�%�ī@�jy�œ	ʎ��kDL�����$F�������?\�W����LF�6�mv�l\P��B$��m��8�sgH�	���V��W�s�3��*��B��4a�S��f�6�AwN^d�N$L��]Y�(E���1�)�m��JRp�xx��@�:-�gSA[�J�&CWί�WN��F��U<A鵴��L���8k[���Z������:=C.��㣪
�}u0z����k�練��g�Ax�o���2����@CY$\z8?25��$����'q����U��$O�O�w��uA�5�~��0��s`��o��-������i�UU"�To���ў���{��Z#�9Q�������Fjc\׎+a9و�2yR�>[�r*���Fl��!�M	�=�)�+�|Y� �Zw�}�i͢���4�'uS�*A��.�@ɿ��"ww��"�>��O;� Q���\���>$�Z|c1�?�ԃ���W-Qp�(XL�`������'uO
N��=Pz-Nާ�|���00}��ld]{�i馣l�pgmǨ�gЖ�h�,m��`Wz1��o���N��i���=^�8k��D��B�9��A�`0�7��j�������yv�WT����Ō�nF��5q�Btj�祂lRP$
�W�D��Ln��q2tS�o�8r��y�<	ѡ�[Hd��a3:�8��JLU�-�{3�2�����;���R�͌�u��4�1ۏ9 �?cN��i���t�:�ZH�
gu�A�/m�B��518�g�aZd���!<��89���� �nV7�	���=�g���)��r�tN��PI����w��u����J�b3��TW�ܩZ��F�T��$����K���eDi�z��躘=�L<�j�5	�w
�ω��x�#�s|v�/dQ�u�E�i�@�־ȩ �7�=p½!�fj���X�'��}�T�kZ$c����X$,��T7�4�=���閹&{�d���H�����R��2q<'���=�"�<��T�4�*5�-<>e%��%����y5T��[�wn]\
��O~XY�a���T*���@���Qf@4��t�H�8 }DV(7a�B������N�/QO���c���E0����|���R^�q�f���6� ̪��ŝ6�v�L�{e������#^/��<�tU��O�x�V�c/b~����"m�-�|�aR��"R!a��Eh��6�'���P���1�'O�"���
|h�0�������r]�L�h�t1�ts�"v;��,�3�xX��a6q9��� ��kKl|Ҋ�#�J��eW�!4���o�i�g�ց��:lҏr��H�� Y?ɕ�#5`ȇ�.9U/5��*���-)��z�AUd�e�a��M�zIUh}��bN`�/"7�����
;���Ll�H6��`��i�FǺ�h�,����dL� ��^)�J���C�!�z�1�ڣ%rc��q�V9kgȰ+�;t�[�`�a!�8���k�O��~�X�B����;�<<�c�#�������Q:���Cx۞�^@��1��� r_MN<��o
ޓ�[�^��`���;���ʶǄ)��|�sz��4�[�@P,�"���U�zN�x�U|�ÎҜK�����&��;�vw��/TCi���Nu�Ծ�s�j�l���j�y��rU4R���^����0z҉�R}���>�>y& &@Y�:<,�R�h���{��&S<���@�?��:�M94�v��]�)Fyi9{U+	�q�/㱋�P%%c[e�"�z�>|�>2_��:/[�0�6�o�T�+svid�1��l��N��\q�ކO���ת�|d�no/������m�v��MC�A`�­������K�=ds����X���	�8Ї3��bD#���JL��QPpx؊��$�&��BL� \��>*)�\ڒkñE׃{�A��7�޼��*Q4v�'O�녜<��+��[��U}�~�B*Β�����7Y����K�L=�[p ���Q4j<�z��Ffgu�0�1���b�+��əT����A���܌����{�tl���� �5�����`�oF�����67�V�:��W�UJ�v�G�_��S|IČ�'�/"�R�m�Z�F8����1�=u� �v,lu,�;�_��
�묲�]�������&|�!�C�G�/DeE�M
GT������x��X��X�h��������G�`HS#��I&�ݦ�M�s��?�s�>ݠҋ�E&�˲�2��*��QB��"�R���P]_�<"�JX��g�*C��FnǼ4�]H?ar����IL�� pl���O���g� ��>ctb���ʷ��ѾJ0�������on�AtjE�`uevg޷�l�v��s��%S�	X�#�2Z�5\�M.u�joLS?��aQ�d���vC��0;EB�#�H���Y;R�� �K �?nT�ȼ���f�wu��p۱ߤ�sC����b�<$���A�<8���h5|�/��`󜮮��vxڧ��������f��	��W�S�s�v�zM��IA+I�kL8�������)&��4���&��d��|x������k�ձ�V���!�I������=�˥��gm����#"�W��Ձi�8KY�[�^rZ�7����68����@�E��A��	Gg����!��f�J-u�?��n��M�,�~�?�U��I �Y��f�N\|�w�ćJ�$�a�Q`t��9�:e ��/#p�geЫλ���锥�4%�k��NF'�@5��ۆ_+o��`���B�D��c�;��B����o���^��҅}jx/i��',Me�aJ�� \4e�w�Ca�� :Nn����b��%QQr�c�����ß���b�)/�H�̼�Z��3��\��qk�Gb����EZpm��(��kX���EY�N2�ڨ�� ��~ܨ�!�0�H�+�C��x�	��{�/|6
ă9�A�u�h�ol%���i�A��b���,��!=X_�>|�
s��ˢ���D6��s����/�f�WpM���	��re
��śe��	L�H�$���S��J��<�JH^(�9P�5{�@�\�~F����wC��Ȕ&2!N:���x~�8�N>Т��J(�5�,$����<�aF�ϳ^��~y���"v���4wc�b�5�b���Q$J��SO��$�2��<�t�z2�j�kY�"c|��c�X8o�En2��w�E8uC���\ 8�R��e��z�R�v�H[��LOK*PN1jҤ��V
����!5 �!�BL��_���j^w�������ğs�J�]}�H����I�ѓ�'j�"���l��U_�'}�f#�UQpD͝l>o8�u�����[�[�y�3���-����O1i�9���0�dc{�u*d�4o�~`�x�4�w��,���M������_f�M9��B#s�,~��>��L�O�{�XdJ��cˤ�(e��,�Rp>u�;�VaL�����'f��=`��/iQ��7��#�����~d��sˬTYNG��w�s�"{��[$B�N��;�O"��=��~��;�y���4���)s��nZ ��$Ӫ����-�9������E�9����Q"M�<���EO�(8� x5�F@�����;�tJ�y�C���W��h�}(\��a���
��y�i��=FP��d������ˢn�t�L�e/�������U�h�̘��yyE�C1jՄ��B�'����c� ��|��l�6LE]��� B��~�L��b#v���D�m��t?;�K����ٌ�N��t��a9����Rz��T�IA8_�$�L�#�ʛ�G���3>�����]��,,�M b�s��'F�maU�Jhk���ʠ�% �B��?��z-�EMᬞ;d����RX�Yԝ����BL�FkW�p�>����Ҫ�[���.�]b�	��JK�/��ܱ����u2���RQ$�����>M�tr�E�Uծm/�=� � R����Ջf��q�P�Zbsm�a�d�b����O��9~��h��l� �6m/ߌT�-Y� h�aeU^v��q�c4��k��I��ʆ��F?D
�sa� MSS�WHة@�x/�u;�-�H^-|�j��Ž��q�9vף�*���&��É�\p��C`5�3�hH�+ߢe�P � ��0�;��ZB�S�UX����) ͟i�w�[<QԌ��D�#����)��1�>�9V�K��5�A�p�7@�rs����gr"02�i�j[]�'M��U[F�v��RNJD��L���*�&�A�*�{c�c��z�ۤ�!��gi�]���*�x�o$H��-ٜ����8a'T�c/k��8H�w
�� 1Qh���f�K-�[X}�4��S��D��%t<�u��E�t�P2;��[y�l���ϩ
e�:\�r�����)��F���݇p�u�G/9��3�b����\qK}w8���`�(-�r�?>��:�_�u�2>����W�t,��T _��Yюt�
��Ä/ `z�L;ر��s�c�Bl�s"Ù8玡�20��/�ŲHИLr�?�A���t�� ԥB�|�eJ�U�Ma�r9����(;:�F�MQM%������鷛���_�m��7u��D�&Q�9��A�	�+�K�uR���x)2(�'_ëx����#H���0�G�[��kLb,~����8�_��y�������WB����F?�Cd�xB�qF4s�Yk�B1����j;�,|?��a�����6Ն��){�,�ݜa�C��;1�|+�t�?����E� �����YR��4 �˥W��D�˚��4qv�� �W�l�.s ��d�(������)i�����c>�NT��7�Lς�6"������x�%�z@���_�^k�C�TN0\$y%x���R�����1;��v����DWx�gIWZY��&z��q����`V�u�]k�������n���p��Ҡ�l8?>LK�W���*Q�	��{*�9������Z��b�%�M��AA]��îb��i�^7�"T��ցm�@�A���T�P��1���κ=,(l����C�Fq��%�qioĻ&!��	ݼ9mߍI�����;p�_,�s���D���W�K��ùi�I�^�i�'S��D�l+.��!Ρ�C9��Ϻ���`N���sD�o(`o��48�#o��:3�;��Q�7�l@<�����II^Why���߮�?5~?P��ר��6��p��M��r:4!-i�F�.x��(�lgǈ�u��n��c���~��..��d��}:����Pc�al{�|�s1��	�J��F-0��
�[J��B�{�5���#�����&��n]I*��n*`�#��s��� ��*���>�K�X~�2��L���׹�C�[�uޚe+E>?�\�BcIz2R�#�8���찭mw�ˤ�����=5����:�+��
P��n�\7չ`�O�h��Ư7�b�*#�8uiS	�=����:	�1��s�)SP�#+�Xc<��$��ePh�S��:{%<]I���ݹLU1Uܷ���m!R����ڢ,OA^�3"����ډ��hr��%�M���{G��:�FD�k0�ʫb[Hl!��dR�ƢҦ�U"b�r���5w�����I1�b.���K6����X~j�u��%A������f��%�� $06�3�4]���ɸu���1��4Q���~?=؂���E��0�鉶��B�����Q�O��'�d���'L�����+ǀ�e��շ����i�9��㚆��>�x%���W��.g	g{�]�/�e�I�F�X�� V��Z�/�ʑ��GG愥q�P)O��	��{"=N��S����n���u���JGb�b���c{� wΉ��'^�d"J2~�?E�_��bƴK�lIWbVu9�>�m;0�5�!/��r��Y�֖n+��Bh�nh�|����AC�v��/����ϙ�t㤨RBJe�|Y~K]6��<
�K� ��U�wm�]K��/c�FZg��ޜ�C�}6�^��:����?)���RȘ��i��ʋ�����=K�X�����u�)�/'��G��Ѣ �A䒲9+�/(�۔sC���,~]R�����Rq�:9���6{M4���o��^�s��b\�F#�ꭽ�����0�:�$���bU��wX���s圑�TW�3x[~)�{����}�����x,�2�Wk��B,z��J�l�[�^�ta�Y�[�_g����x-v >8蹊e@�^�צ%�s���Q��4�XQ�pV� �~7A�҆ ��P�q�y �g��0��K�ю��m4>=	p�d�����¨�Z��&���ְ��}�e{t�7Ni?d�8�t�O+Ia��2i�U{�W�����s�����`^��i���5n&�1��Rqc�]gОf�����M��aCq'�cS�׋��X��,v�F��A��(z��ܴ_Ķq�>5��t���L4�#s�_�Ϫ�+V�{�G�z2i��&��mG#���Z\^�=M�c������
��!b0���R��q�I�4B�9 I1^����	C�r��?�jZ���E�C��8¡�Z����*ᓐrOk
���d�u����.��:&ݭ��A�W�[�
���T�f��p;�11I��6��8٫֓��v��!|%��G�+�mZ~"�hE��^7X�7r�i�}�rYpWY
v�k��z�+}�����CW��5XuĴ�1S�ϗTw,���e��n����T�j�y���K`_���R��m�a��� ��n�3��d7}9��a�af;e�C�n���R����Ѱ׬1���3~[���4*�|\:�ކ�^6*m�g\��4��ɨ?����C�!�WT�Fv��pN�U�ol��D@�~сʱŽ^@�A�2#��+e�$���$x�A+���&�Q�I���w�^vB�E�aC;�'������RR#3�x񢙒��D(��Ӵ����XV~��V�J��z�z�����R�����%��($z�o.�t�]��-�n'�����ɛ^�a##��͆���B�Y��'���j�Ov�Y�=��O��7�h-ˍ(�tX-�g.�.��"\�t�
�'�xx�7�Q�#@W��ջ��a)MS���~zU'�+ZϷ>�Τ�t$AC�ɢ�/zxF��JAPg�j�w8��S@Q%!�P�Dx�NZ;��AB�'ԧ�#�U��, �)A���;��@��7�9���/$z㻉3�so�OH��t��E�
��}̋��.�o����C��Q��U2 jq�Y�<[!V��z{���d7��9[���MOd�
��i�N�U"�m�* 9��+ �#���Z\�Tr �&�]����ȡq��U�)�C�m/�)
g.�z!��1�U��30Y4Uh)f'��TU@=`���"�n����}����I���_ϭ���ʠcG���h�Rj,�F2�;��[�7k{����I��]�uf����'��t�1њ�$�ZΑb3�G��fH�9�m)}?F[�.&��yИ��J����|�i�ݓ|�(ai怶(;`�$�L���6��*��-B(S12n�l�`�=.o� �c�@��zU�ي�6�\.�&�Qk\�G!nG+�[��6���q�CR5�Q:��3,1��S������>���nd��ԯu)�������]�����Q�����ě���
��P1�����]X���W�ੇ���craDv�����0�TY�"B�9(��Jw �����jt�-Z$��X`�Sq�������R^s�<�Q
x�T�*��^���;�ۋւ��Hs*Izp�=J-�M>dy���5�~��<�w#�O�9 ���.��u�Z�qDY=y���KK����ߓ#Q�b�~'��!���N���ȍ֬�EӘ|���Lk��!xS��
;�D$��0Է�cE�0�&KQ�؅�hRr�Y8���%�:�IG�a��v#�}10��(Q��h��1g�F�99"[��)5Pб��! yʸ��E�Tq1�Z����%�u��l"��wb7����v�I=������I�����d��jrm	j��?o���yf���A��IR�3?��?��1��ljИ�TԞ�5U���qxfS��HEi�n�J�V���ɗ�]�[�d_����j���G�:d��{F���6Z	����Ĉ�fT�IH �&�kJ4���9�{~�m��Wf�⻶&�O[ϕ\��#B����,`��2ʿ(���[T�´��7Q���$c�B��n���*�7�Ux��7�+��L�1T�>ԙ��Ias+"�}4��f�5���:�A��"!��wD/_lW�&�;�	��u�H`t���1�jd��ak-�`�H+(u;�	�$���\��I�z���=���F�q�W�$��l�7�ğ�IA�H�K��4��y������C^9����]��S�]4��9pZ��jZdAӼ?�"�+�a��P��x�6�Q�o|����@)c�����>�]'�m�/� 	�I�8 @�(��|�ZI�Rε����({������p�E�t�e�u��Zm=�X��4���<�V���Ӡ;P�K��3�8�{�Mx�����kO�#�8�I��R���ȸ����!�|T�kR �m�G����ه�w.��o�g[z Y�[��z�*@��|b{���n���um�>WH�����Z�[e����n_L�p`���:LI��+f;&H�}���
�Z=8ФZ��T�J��K1�-W��+����u��	�&�eWx��+��g�D�5},�$��~���q"�ٷ�&�z�%v����B�sD�hÔ�a�܉8����q�(�?��-������ �[|�
����X4�$È���I��W�/d7��FjO쨩�U8�D^�$=?:��b29���Q�j���0�8;����L)�������V]^lg�j{C��<���S�����^��;�x�̫�b>{���ĳpL�$/?��܊�QXJ�NL��|bx�]�XI*<�����#��сuho��k�1��^�����s_9����9a3���F��R�H5�Q,�綷�
`m��k�tQ���"`t\��F��}����6PuN�'��M�f����z�4�U+���	��N�"���<r�'����5=c�S�V�,��wW�H�u�&�Y���;Z̷��8�rc5{z�,��/Lt����F�q���GJ�W���� +�_˪�;_ѿ�h�o
�gg��K��.�Q�A�*W4���æ�oZɹ�:���MG :�8�!��u���J�W�ֱ���Y����|�w�Ȼ����.*�՚�-��s��ozT�k��b��<6����I��b	6%wU��S_��_Ћ���z����[E4��fZ/]1�0U��v�2;�O&�n���}�R{�*$D��_�)\�t� P��̺"˻�|��	"���d4`2���c����q8i�#�/����x/8��./�н]v�V�V�."E�t�-�1���(�i]��*�5Jˑ�R���>/�T��2�9�ݩ*ٻA�k���3L���[BCŏ�(��Z���Jy�G�X�6�r�s<�1d7�9O���FJc�Dx���@�咥O������S���+?����&�ߠ}�]'Rο$��H�uq7����Py�hnBpw-��I�gax��A�֋9��e ��� �6
�:�d -ܣ��>;�At�"^���9ɟIїN��N��Fw�m�mk�#K��p�b4���%TW9Ł����u�0�_��|ل�շ�SxOa]z��-��neBxm����ko�����r�<J�D� ĶK��/�ᨶ���e���H`{���qm��8J���M�ߊ1��a�����bط#5z�/�R̠��똷�M	�c_��]���b׮�}�v�0�Ӊ@v���jd���ֶ#���#���@��K���>�.�N�����ڐ�4�έ��>��M��O=�eh$c4��Ryڳ�M9�
~?{*U��1��O��ќz�|p�c�:U����yY�zT��%q	�5oi�v0���/3ȟs��R�C�}�ipIK�=	?pk)H��r�Ƿ�i�o�E<}�0)��pm�$X�Y��~�0L������.S�M��7H�kO��CBXH�d�b5�p�\{���ם ������� Rmio�K���6Y|���$�Ċ�\:��	��54�J�-[��4�_+��"wp"���	a�饠Y:?t���_2wާt�����U���s�W�>z�rVV?�[Ȟk��l�'���1���LD��B�oL��=�ZI��^i�+��Ú�9��ɹ4�����촠���ZO��pS���9��i�h��)z��G�'b�|�ކ�L��řki�I���':S���qUڈ�4�q�÷���vLs�+��#�ҿl����q�xm���h��B��!��q�+�Y�%q�H���r�2PX�3�f��B_����/��U�a9s�5�� 0`����| H�<n�u߄�?T[-*�'Y�l� w���ke�˯����.�<��~oFY�y*=CpDs���MC^�ĭ~g�}e�ö�ŬC��
T�(������d?N+�v��H����h������S��WJ���*@��QZb�s������z�����Y�Qj���k!�jbg�y��nC̑���
9��{$�L7vVC�����:��ۛ�C1�v����UJ�0EP=G�����k4(^��8��;����T�;���@�2/k����`?>&�3!3'��\iڐYI�h�b����=�S��C���N�L��6w��b%�ߊw���뀱ӑc�Q�u��kx�� 礱P1K��%����u?F�Zo�J��fVW�
o�P������~��me�c�p���/�#o�>�p�������F�}����NA�0ɛ�C&�h�%���;t��̳l1Щ�k#���x�"����nv�W�z���K8\�X�I.�`10U4����B�	3�e�r�o�����1�
"��KuB[P�7���S��|Ԝ(i���D�ˢ$"�-�J>�X� (,�0A|S�<�� �JT�Q�j�����cD�%�?{w�`-�{�iڬzs/����w/iػ%ԭ�k����|E�����}�1�lM+�s ��H����O̥����<ޅC�W��q�V3� Xp���]x�{�m"�I. !���ޓ��J��eQ�"���7�������=��2��D�7���#��,x�Y������	~��CSoEƌt��u�."��>�{c�8x���*�o��&3��t���~��'��� &WB~t��o���T��H@��V]]%�޿I' ��ETkH�Ցs�i&҉����os��7p6��m���
�wL@���G�I�'�S�� �7�0���0,T%H={{*�G\7H�{__�Ep�f�����)��u�X��}ě]��������u?��4�B.��\o:� �c�/�^�C�K,-`?�}e�G=�r<A�V���չ�2/@��ovO�c�A����}�a}J):��l�%�t%�CF� k��#��f�R�Vn?ӥ�����w����0���#�l�:�M������R,U���h ��kBm��R]������ZH�Q%x���z�Ú�_H����:��q�<��1��H�}_؅�:�9V~+�<$z��i�{HPu _:r�T��p�=�n�	��+7YV����1_�QrK�8�nq�U��.*��*8�KА��D4�:DU���I��Rlj7$�[g_��x�b�bR%	C�s|Eh�h9�r�=�,���
�� �-��B�N=��+OYd� 0�n����^����fq��,��~���1Z=�.mr�T�|jƬԑ�NË�钄�p�K����"E
��y`���o]�7Ty{���j�W?�#��w4971	_��-����3+�^]�9�K(����ZP��iZ�>u]���0�����7/����xM^���9�Y��0<;H���qud���hO�1��u�E#a��=�����͏Qu��f�n��kTt1�/}b0+��i��2aO�*��k�m+\�A�G�9�65��g1sul��z��q�#�U�>��3&p��_�A�=��G0��/s�"�H�.�=DķK5-���`p�ax���d�Eᩢ:�2'��,_he$@A#�k��ڧ�_���F��si6�2z�Vn�]�{�����#j��֏n�˾�iݛ���V��������r�K����.n�"Ip�dk�l�āuH5�9�jTQ]z�_�K�8�4۵��R��X�Ir�#A�A��jYDE_8쫠\��'¹$j�d�Go&L\�e�2�i�x��SQD�D]�HU�k�����4��uw)�S�Q�o�����
����+o�����&�#��Uz�ڳ��ԗs5�����ɟŋ��xi��lL��Sˤ�T&4�jHcE9RZ1}�'�%t)��(�VW���S?�BP��c�b
t��9+��/"�����m(Gy[�'/��4<8�
C��¢ ��ٚ�X�K^'�e���55��j��e�G5�w�0�$ �;��%�	�@����$�7tp��>U�Q%.��Qm�~h�yK����m'�i}NI��,� C1(@�9�c[3��-�>w�X9p*D0��8-#f^00y�aL�N���_
e�/\��x��<� N���j�ꓐ�X,�;_l2�6�e�LG� %���y��)�zW�O���RZ�:�S���Z��-%�9�9�G��w�I�ÂO���
����ے�J�|%��׹
���vq�s�*�@Ys��%��S�U@�7M��(�P� ��[�����t���|�:]˟�D[���<�������Q�c����&��]"�ݬ]~rH>Z��$rp�']���a�C5�z�w�̾�`Z�~;!ħ��cfOi��+N�;�W�jCw��>�и�Zfr�	#2T�	i�l.��|t�S��(��g��3�mQ�]Ʉ)W�����, l �kd��>
<)0��u qj��uY��	��o��Aqc��[�"��!U��y<�@[�6b�?+
Qj4��
�S�Ϫ<R�˾{�NĀ�@f� �a ~�l؜x�Xw��=�,@�Ռ|��N/���ٗӐɋޯ\�ަ����Π�����h�W�	�	*���ܾ(�`SVѡ�R_��,	0��K?�W�\���R8���@�5��m��-×���� ��L���V}�5K����T���i��7�,�kg0z�r�+�q�F�vWL�x�'7C��C�"��������BZ�O,���R[�`{�ܩ��˜�2-K��M�&��s{ೡ�I!(b�~L$�j��zSe��b����)��D�OJ�/K�DG��|s1A��yq����Xeb��V#).�_id��9mm�.���'MЮ���Keü�-X��b��\y,�Gb�L~�2\f1�[�t[�q��5���dA���ׇ��/1q��Du<m�Zź+R�~�8�����	f�J[xP�v��(���":1��8#�������3��6:Y

�d�B"}�����%ʝi��~]j��#��a�K��?�i�� �����?���QK�w��b|i@�� �R.�;9�0�RXȬo�����O��+�q��c�*�v��*��b{D=,��ԃ8/҅��r8H��>�G�dB"��/E6�k��rͽ��Q�q~qH��V����j(���l�y" P��Lq��_�s��Q�?-L�wC�=��3p��w0������\�N!�Gi�X-W(�P�Ć����k0b'�!T�7z ��e&X`��ex����E-���hˤ��t�?荞����W���'���A�c3L$B�X����ٍl<P`�����x��R�^u$l���\�W ���@
B;�<.�I��Oe�z~�'�k.,����ɥ��;�ID�O1�
~�y�{��a`v\�P�۫��k`q>@�C4Ɖ��ɟؑ��,��w6�o����O� ��̇���`�l����S�v�^�ˣTq��Q�O���(�C���Oȳ;���m<��
���nGY7������ޠ��\U菚-�~�׽���E�vK��{{�7�B_�t��2���8�M��;$�=snW�)��}/���z�ۜajU�cT'��G��,���O[�H�^nJ�6�fn]6�}4�������@	҃*2IK��[	�!D6��6G��/hXB(f��G�D+ɕ�����-�����f�	���B\�7��9_��U���x1Ѱ�ԥ���`�	�{��8�!G��-��V݂�P�.�g��ɑ�
f"+�4���/�/z�����3�uN���ľ<')���Eg\�#	Ѳ"�&z�����UʗV���$صZ���+���	x%�e���A%A�e�k���������=(b"�d���[�S�y���Ĩ�Q�Pw������$A$�V>u`�ю=yר&�1��_�n'�DYU�5��pD!�,�9�u$���5A�r�呭�4`p礥�^y������!�bπ�]'����H?�u '+�g�_ ���V�ċ ڒ��3�J4��"��\�>��b8R��y�~~�p-w�L�8xj���qCπ�[1�!Я�Ja%����У�7aq�ߎנ^��&�yI�^��bD�t���>H�Ʒ�H���}Qr�߈��j��tB���{^y��1Ȧ�����M:�euH���#����R̮�Aڦa�P��t�R"8����U�p������-g�2��'��e F����?|H@�� 󅲻.�m�Z��7��͘�O���;���D��P�8)���d~,x���.�\B�{љ��*���"nV.�$}Xk�9��VwZH�P�*}��4��*�h͸v^Nl�L���2���M��m�NB�\ș*U�{��(�8i:�"����ss~a��#�"UӼ��Ԇ��D�.�߼�[G�8�y\����g�ۓm����:`|_K ���ר.�ץ��=�"hH�n��#�~�}�Fcxf���Yg�p�)3�-�a콿�7���,uy$�#��X�U�}�g�Y���{�C���H�`c��3C�y8�|���Z"��E=��s'���=nv�&����X8�1j��>205���'Y�\�SnhZ1�:Y�E�����a�me'���MJ,%'lb)��Zws���6	��J�{����v���a����f���m�M�����j2���~HE�ⲅZ�[�G ��i�X���\2�X��]E�!44:h�"�ƻ���*�$qn�|����#����3���iո�L�zMFtC�'F("a^|��}N�5�Y��ߑL��?��/��\�_�{��R��Ow�ՌE��{�tF~&zYz����g�|M�>��0/˖lɚ�[JG]�(�N����E1����>��۝?̻D40��<�L*��b�"uk�& �`��'�n1��Y6b�m^�0%vS�t��R�|oE��|�
Ì7�VbX��M��z;z�eL�6*�f�I�y�0XN�-(�� ������5.~�������w_�"0�ס�(�����	�P��B{ӛFٱ�U^�Y|��h�&�!6����,�7Eԛ���ҭ���iL��o��B+xб�]���vS��O��>������4��)�n=us�����2ﾦ��e�'��6�DXUݙE��_B�	�(Q���O�����9z�D�y����jġ�م��]�.Y���>5��'������?�D���m3������lh��eG�#zJX��hԣ{��o���C|=�:&�`�(��̊	S+W���E�7���!8���(9�^��_O�{0����K�Q���S��R�z!��m��`_�aڒ񏎥X�>���i-���
)�C*ߕ�e2�k�!�Z�C9&4}q�|��� ��4krYAHV�f�lDgV����G60�i�,�]�y��D�e�2� �p`��αm\H��P�hu�.ݟ�y�O��/*�:�����>���4�����N�fj���3Ф�Z���8U���Mt�ئS�b��ҝ}U����:�h*���8Z�i�B7`������>8��C�#�|��$���[�@`�����B�g(?W�>qd_I?����4��&��O��{�\��M�\����5�F��bk7L�� e�-�2������Ђt
:�_�S�%����)��S5~{0��k�ױP�p�AKr?3Д�����U	09�����n�o�W�Ǧ2�?w-�/A�"������թ��&�I�S9�D��4��✚�X����l6�=%f�&rr�S�v3�u5��
fzNe%���-f<ٻx�"nMI�?�m�y�'(��?�H��4cҀsr�ۋfu��!�2��@I�}�V�?����^W�����N�7�gF��3r����z �FI��2(��A���d�����Ğ֊�Dc 퓇�c�M��t����ԝZ����ݙ��������bY�Cd:I�7� �С�#bo�dE��]8��#W�[ϯ�y�׭�"F��.�H�Q�x��@,'wE���Ɩ,��>CV)�@j��Κ��^�Y�'䀘�o��-�R��+멼���"������8	xN��n�FNQ?�s!�ҩ4nv�9r��XrD�v�C�t������͏���16>��^2+�&H����|����;CM����$G!h��n�F�T��Dޫ�<��B��iç?I,�;>2;���5���X�(N���^���4|s�v7��D$�C �i0��%�"���|6�J�j�l"�lNZ��,�&��	�y�I1��"�#�:t%��H���yN+�[В�O���eq�k�������c��V>S������g�Bb�[��<��'���F�+b((�zE�c Sq��aw9NNچ;�4~M�]��k79����)"�O�^��nty�֪MJ���7����txG��I��_ӎ� 0��������:�� �f/-޲��͜�j.9��_�Fr��}S,�f�?�o�%�g�[�FF0�M�^)�O6����UB������ I�_���-�7�R�e��9�!x��ؘ�t���EQsk,��ԲQ�5i�X�aQzވ5��Y���BW�

�Z��`�yW7�~�xr����fiZcӂ��L�b����/������Z��.Č0�.>�Q�Yɶ��^S�:�i��q�7�~��H�Ç8��*�z�&o�+M(D9,���u��gֻQ����	@yGqGTE@!6�e�p�7ly��8��tűfx$���h3>S½C���������6o�wb����=��^/���b{��n�f_�6� 3���py�S��7��*�o��I��7�|(�Z +����
S��n��C�ܔ�,g�d�k0I��oV�(D/�~"!3���ӟ�)�8}6�` ��k�@|����]�
(��������҃����|#�o��	�i�+��hY\�m��݀1}03�>i9��;�r(Ji����>I��6���q'�wR����������eC��f6nb3��Sk<��"�Dh�HGm��RX�_�e|'ʫ%��{�
|�u���ł��
�0�NF��:�\�<~��1��OE]y���-�#��s�`�0S�F�:�/Zj��.L�[���;�A�]=��xm�9з�gjϻ/����K�b�s���	T�9��/����S��~-���H*�����_ꦡ@_�J��%gCQ�W�2Փ���^	$��q*���?�VnZX�O���`�1W�ϖ2W�YwkɊ�E=�@n[ �!�-u'HT5*����Y�MX�܇SU�1'�@,{����<��P�sY�1r8˥����U�S�mO0��B)�T vPtT��M��{:>w{md��<s��̋�a5��1���Nd �B����L%���{�Z���\�Ym�x��_�/�&p�%��:J(U
�4����>�\��=�u��T	J����S��Q_��T�� ��\$���Qk
��jPK�WY5ry7U'@Ig4���2��fGK ����~��w;������tT�5�z�W���.���b�����{�'��E��/��H��-B�;U�nX�f�eG|���_d�6�?�O�3���B��h]?��r�OH`�g�(�n��
{1�{�
��A2:[��DtXX�Q�И�Oí���>
���-�g�鉋�!����UwݩDExv��ҋj����Y! *�oG{�p�pA^�u�ķ&n�����en�x�-�Ӎ2Fꅙ�(��������Χf]�w�-�|����ㅺ����m��H����8��ף�qy=��)}�AP��"`�7�A����0�OZ��a�5�{��/պ(�B+M	�X�;R���"
\h��E%L�l�'�����%��%E���<�y�(��'D�+cB�˝"����݄�"��w����;6?Gn�X��6�`>���s_�j�4b��c/�q�+��8��?)��t��pmq�c
,��bg��,�ٔu��/�P������>�~H���|��}�5�u�<�vd�X��Dz#0U�q����YqhP=��7�3�mbh�Df�İk(C����3�p�3�M"F��=m�~C�J�|Ş���Z��c�^j�D~`���m��>G������"~�tc�CGV\Km�4�#6 ���RM�.�.݌��/N;�����I=s��Ps��o�3�Y�:�{���Iɱ�� Ǖ�{uEQ��b'�G`�(���m��X0ڙWLϮ �f���^�HJ'%��"�(Ý&�L��D�Hs�� ��������6�e�J�|M���� �6/6��O0�9��"d�W1� -�Fp�t��As��^��`����u�A�л��VG����d��[����Z����;�V��M��p==V�twB���FzJ}{�!c�����Vu75�Wn��A�y��G���k�̞�c�����<���z��ML����ķdc:6��vV`�pS�~���,�sv�lb4`�$қ}Oے�{�*�HbRۄ��0ۊǦ%l�g%	�V�J��2��I��R"�����u���`8D >Gn%R���h#X�O��]�=�`d�ز].Q�@`N����\9K�������q�ˤIU���7e�0��TY_������2�b`do��⩃%�e����ш�y��E:u�h��)Q��/�S��,�X#26:��Gg$~��mp]��d����Xvk�qx��\4wd�c��H�B��2�% XXl����w#]q��
=��Rh[�V�e>JJ��i�H��%�-8H�[YG�z�#2X���;�$c4��������{K��	��,��ؼ��;�y�x�cu+��a&��iFL +q ��՘��Q8A^ƶ�"
t��C��|'��;i����CZ8��~�RW"���J;6;�7~�I�	|�g+�;�6sN�t:�ċ��h@��\�˟����|1��t����I��:LǤC�C�Y�cZ�!�w|2惼�\�F�q9�O�8>\5�TSe�I�4�Z1XA��m�`4c	�^@}*"|�W�@�-w K�L�_J25���
Gu�����}�5I�2@Zq�*5�~��Å�}�1$�� ���T�jfG�?�_7�Df�U�y5ۗ���� '�[hrt���lbB��]���w� ��0�X"�	��YW�C>��s�=)��Q冮��5���M7���Ք�Ug(J���+h�wP [ڰd�k�\o=,�L����.C�p�8�i8���W�5����h��^�xHE:���B���P�y�v��)ŎE�y��YH��t�vϵ�sN��*�Σ�����u��K&��x���+�ɫ� UC�I�V!��q7�Z� N��O����!��|�* �����˿��`-zӴ>�/�&�����R/+輖{�O�kq~6�6���B��&��1Gc�o�־c LGm5~Ѝ�j7K�_p3�:	��C�/i�.y`�0��S�m�c㓣B��
�>-1��X�Q�S{k;:�Ĕ�I����
�����G��^�����3�����Ӎ(�N��yÜK���T��$�;,ZMȉ�jG���(�.� ��'��םN���PCi�/H��I���h�/����H����lS�_ʴ���2�~�&"�X��c-Z����\����tp�l0e�}�r'B�=K��y�I����3�S(����z�dX;����d���1�����M����)hp1��^��,FW	>�	�K"�~z\C�2�F�T8�'V������lp��Wk6����T%״��!r��M�,@�����gǔ�v����y_�}�s�}��?+t|Ҕ���rf���V3��	7�S��w��%v/��a^;eӿ+����c%SG(0���q1��"ɏ���x{*�>�a1ꦟ�n[A�n�^P�2eW��Zk{)�Z�O�y��8M�8�����ȭț��i>��f�ѢY?�u��_C�1�#���j�;ϺG���d����fʴF��rE|��ok_�L�-S�bIͦ�>��?^9DG3�a�xdIh�#���	AD۔�轜_��0b�y*M��.�~g�2���.ԟmם�*As��QY�@.l X_,8T�����liď�@SYv?9�j��$��u/�0$�R����ठ�5��=���e�9�?��Ug_�Ip�d���.�|[�������&��@~�T�g^�~vp�!J?��0���:�[�Wu�&�ۍ7�=���O~9��}qz�e�oV����c׈�0&Ȱ45�6� *LWÅ�I�Y�7~����0:NɆ�	A�M{z�OA������%b�0"��8鷍��j|��Q�/���D�2��H�x,<��!w����0���0.��OdNF ����i���B�,~���-�'*�������JK���e-���A�˄_�+z�1��h%��sH�,3`����4�P�	�eH������NW�~&i-�l�zK�����S[�5ET������R���c8��b��6?�U��D�ĵ��!�W�R�:D�i�s?�ӭ���,�[�_=+)�j:D�DК���D1��&:�(�� �X ��w	��C�$���`̶!h��|,{"'��JT�,2�bs5�{�(�������'�;bdIoOvGns�gK�d;�F�-0����>4�ɥff�V9�}ICR �{ۚ<�<<i¿R6R�������[2�_	�S|�&�_���B�#��w[�Ay��� ���V{��|�VNj�,^��í��"E-C���S��L��:@>�'�qh�A�R)��֮��޻^ؑdj����{Tz��X��O.N%[�R�zp��ӟ�w$�v$	E����(��HE�K�����2[�����X�ÝN~�G����j)>��^0���l���G'��5�)���Y2�;{�H��o�;Y�-;o��>��n�����������2�D���:�Qb�n�1�U�f�vB/1�2Y�aS\�!c^����{��E�W3'\*'D�buE��w����lE�(C�6��=�[��� ��>4���W����0�Gs�ߑk*�_qȺ���xp��*��0ͭ�zM�L���d� �8��jG��`�2[�� �eu'�MDrN��ǣ������Q���5�g��+w��H�1W��8�~IW��/��Ҩsm�.�����Κ��UQ��<Q���OV�	wF�+�KҖxr�(0I[K�ab�:�"�,�>pB���r<ǭ�?��4Y���<�>�����^ /��,�����
F��[�$��G^t�z?es�Z]<����L@LL�5^�A�ʢ	�O���hD�:ȶ�������*��*�f�V��Ȃn^0� cBoHAjK�_��y[$�r̪�S�>.R�h[�;��<|�z�Z���� ������_��Ly��|[��j�|�a�@^���g��ƞ%���.VHO�/A������\;䕼��u�J��dD�n"7,��b1�p���#4yQ�C� �7�����C�,�|۶�65p+��f��a#���zX�ѐ�(x��C�6�!?b��/=<�r�U�J2e����N(h%�j��S#D�{ ��M(�?����&_�7*uH���s�U�v;]�~��=��Az���&��K|��R����c>�y���>��m�yD�c� P7ږ��ҵ,:�:�����
�pjm��F-,X-����6��B=�l?��q|�Iі����aA�R��3pRy%J�l8��7)���t/��@�;��ER�t�7��Us�ܫ|T�D�ӫs{ލ ]�7�&����~�<5�������	�d�Ann�wH1�.�%�
_-u�Ղ�#�n��b�Xd���,��Ћi;*C�n��c����swFI C���^H��2]�ˍ��:������/��e�����_X�h�StKM>��e��t�*9�UH������f ̸Қ:/��hd�Z�Xd��_|h4�6���	�#��,=��b�/6]q�G\�H#�ۡ�_�����,o�I/�UFP!G���9�P���$�;�b���>���-��	�dJsIxK�F.�!�=�����s!o�{W�.T�
��N���8��.��qN(C��UV<���-��-��^���W>��PE����� �\�k/ϝ+�,�
���Q�!ʇ9�#�(/��no�l�5<�\"*�CY�w�!.���$�8�m�N,2默UȢ9@��'��y��_@��O(��ߺ`{b��֞ly�eY�?o����e�S�0�p�E&�:�x��׏j�ˡ���ȃ��I�&t����N?�����j6�~h!J!hN���^�O-ϲ�ȵ�Th^��~R�NT�
/Ly������C�iH��_B�Q:�*��L"yR[#nd�>���nd�����1H�����]6��J|�/���M靸m���c]�/�7��T�6_�_Y2�'�_���B8^ǹ���@�	6��$�g#�4T�!�����w�>w���%�Rf p�U0�Q`֜�^Xi����O��Ax]��m��R�b��
���	pŠ0����W�� q���'1]c
������r3���C�Y�������==�<�"�&���CZF�IQiR��퐣��12�,;���(�j���dK�+�ToX�l��E1�1t��M�����m?�zW6�s��k!�WWh�ᯏ�91����y��Aʉ4����J,o���|	^���<��1/�1��E֒�i����T�{G/��]����ؚ�=8�=�w��k���)j`]
K�E�`oz���`���Z��YI����l��&�&Y
�����VJY�*���C�|��2��� �Eu�����m��UwҮ�L�2ٙ��9��G0����F�ɋn ��+洧�� f���g)�<���-�OD�	B����G�f.s���3�z�؏(H�˚@��Zۯ���.X�����K�g����&��Ҥ�b|��IH_XG&���l1��z��Y�JM��:N��L�����;=�*%�	)V��|҇��4�E���s��4��wDeA5o�{b,��(�]d�є��lG�l��עH��5߮�I�"�$ﺖQ8�?�I�S���@p���׫]���c�D[�+S�W���-���S�	ܨ�v7r���y��k��s+ve�1%[;�����=j�-����QU��T���p_�ZnT~Pn��wo���I��(HM��tש��¸J�Q<eH���&����������!r`�ڎ"�A��nt����e�ݕ��r���d��|�?o���{46�T�&�L��$at�="sѫ�vke�IY�,m\Kvg���z��6'9�û]�_c��[D���a�)3-���Cy��-M�/�q�^*��8�=G�����p?�~�2�� �ࡩ(�Mu��,O�� }�9r�rq��[i)���V ��"�Ů�wR�iW[�G�y�%`�,���y��I��3�ću���e����#~�B�ja��z!��z�~�m�l�m��J��o��B��|׆z{H��h#H�L��;]2���j�J�����uj�\0��XͶ�0ju0&��y�����rg�X����J�{�ӆ�(`��a���N! ��Ėqeɾ2�n������*P�_��^׋x�H�n��D>��'�}��L�B%���E��v��0���9���u��\�2�8h<�`+�E�����w���r%]9�x�xl"Ǿ�_h[	�ͺ���,�s��Q)�t�U}�*���|��r�,�C)b��a~QP��U�tM;�a�?|)��FYN8Yu/c�*�9��:��)F�'>�Da�R��Ձ�Eq���ΐ�Ύě^����P3�o�4.�h �M�	D'����+8���<��,0���;B/V�<�?�
�gn���EU�j�"�t;^�$ӷƨF�k��@V�m�C��E���k�	����sN�mE�q	IM�ZZw� ꐼ�5��D�d.^�6���
��E�z�k��7�)���rΕ���B�}!�8���6�֮P*����طP��B�����{[1Y�F��(����NᝪP�?�>���e7�}����Jв!i��a�o�+	��*���0��RE�<|Zٯ������0Hv���U}A�T
�yb�Qȕ� �H��ؙZpV��
b�O��Yg	_�*)���P��l*�GJ65����U���N�ƻ���?r4��,,��h6q) ;�������!�B�����&���)��f�o'`eR'&Ū����n��7�?%���r��
R�GJ��.F!�:���%�5M������E*��y"ՍPa��"�N���2��GHtk;q͍N�<�������@c��)5�Q�Y~�{��p�'j')LX\&���낰��6�h��$QD�W�|��ts��
�«���]2\�Mq���O���h@ri����0����5<���NA�~z�iBu���\��jrq���ޟ���\kv�a@�<�4��Yq��!`Xb��K����rǬ�h�F���P���biקH��[sg�]U�����m�d.�U�;y-DC�~*�И��3e�c&����
u�Q�!���)�XL��$:Zy���wg7�
����x.x(Ɔf%G�u5 5ɱ�qk	��G����e�xl�4^�꫞Ê/�g���W��Q�D���}C��>�i��� w��弚��̶���z�œn*�;�\�]�9��
�p��l�NS1y7(>���$@g kl&b�S�z�%.���
�!Y=�l��)(AK֔�F����PE}3IZn�@cL;��P��xxud�@�~g��z�\-�J��:�g?&����׼�/���n�ԭ'Q�B~8>CZX�� 
�d�-�5C�O�ߝU�Q��>���I��r��vDU�A�0G����iH�.&2c�F��1q�uaD�ĝ�9_E۽��렮r�C� /�j^=�t�����2,!�kn]t�j���P�}z3�\�@�u�d����/��:l�S(js�`0�=ϳ��Y9KS���Kk۽`�|�̃/ȫ��2;��f��"�j�EX�o�k������](>��p��"�`��5ڸcTL m=+��D��^gS�/�4����>J?N;���@YX�A�G�^6�.���2k娷�<�B+����r�j.��<�JJ����s�j0�L��$c�tq����H�E1��Ǻ�$�ѪV�U���(�3��p�v�O$?��6X���Y�K�u���4)\�P���㇧s_��@`n�L������sp��#�Ѵ{���PZLN��S�f���8%�|�.�H0��HSg�a �h�%"�=��:�a
���^Ʉ��\�Ɣ�AE��#���/A� �p��$�w'�
P�jb���{�a����q�]�;�/OPM*g��%b�W�0���}Zi\�����B�x���Y��-m���E"s��좌+�<x��8��g�ߦ�a<�m�eFA�H_ɐ�Oŷ�	|�$�l��_�zO���[ l�u�����BԨբ�WWC$o,#W��0���yLt!��E�lݩ��\kY���T�^���g���:�D� ��֮7��X��
�mb���Oo�`�,��Gyp	G�\�K���fز�Pbdꋷ������N��� $p�.�|<�$�cN}l�Po#Z��f�i�Xz�Z�ζ�|�q͟�-`z3���ʟ&y��c��J�l���ֲ���d��m���7a�?��:���Zh�SS>�#"J�:�����n�O1�me�޵}RA���-Mw)<9�*�O��u1	����k���3."���}����8��y����y&2Cb-�,��/�̱-�� ���˹��f�>���a��a �V����s��o��G&z�^?pI�o\��<�r����夈��ݪ���J�㈚����)�^���l!��Q�Q7�,B�&Ϝ81"�j�:ٸ�Ӷ����{Sȝ�6���߷ECc����7����AF�+�wH-��V�ܵI�����j�l�`'��~h:�V)H���hhLP��@�dT9��.��/��K�cc��F��8Ij��U���X�L*p�(�Лd������]ۨ����z�ͤzPg��S�������B�/�;�E��=�<��80��Z�^%5y�R��g�Q���'
�O�y'���ǩ-C�W�?�KV���#tF]�E���2RIu�X|�Ӛ+wʆ�<���]�Tt��մá�n��W!�hB��׊t�s�j?��>qP��V�@�@Bߖ��{3�C�ǔ	|G�BJ�nsf���!�T��A�;��U-�p_�}����#�[q��g\��������;a�hz�M<�_'��S��ճ�{�K���8ؗ�^A]��ðS��g-�5w�����QYV��qM�H;DO��L(S���%��U˪���._�>d(q��*0���@�W��-�׋���Cs)��Y@��V��6E��AΏ�p-��� p�<~k7����'�DC��R$ �ӡq����\d���e�&P�@@=H�fpk*�`�:5��Z��|pU��'�\\!����¡�(�[�?��)	\�z��!K���Og��( 6Q�EA�)���.��E�b^��`�|����x��1m{�4��5d�,���4A��y�y(֑���=:|�!�AZ���R~݃�{�8�5���y}�۠.ۢ`�B^��%��� J���I�`|�D)�?�u�\��i���m�'����	�f/���J���gr�����c訅�*I�-4��e�O�� ��2��e���q�|������N:���&���l�*�a�cJ����@ߢR���|�2�{�A,6�L`45>K�����$g�׿t\*�J�*S$�n}�(^n�r9���?'^~և7��#e���7Y�_���q8����n5˕٤oc��1y
���#�XB�k�
  k��~$l�%z���g$��y<$���#̉��V������m�g�|��n殯� ����"��%Λy����U!;��^��1���܋NO�3qqq̠z�lC�b�T�ڙ  7&��k*yDS)�.�E^͞P)��T�g��,��~Cw���\�����ɛ'�ۉ�hR2_�Ws��+SmutZ�*�r�o��Drs=�ɿ*�Z	�Yne`�Y g�c�M�ά9[U�!����q��ū[��� �@Z�<
i	�d�4��|�-�MOLg�{����ʌߍ�F�5�e��S����v3�������e�+��LON ���!����&Hc� '�fk΋9�S:s%�s��`��ݯę���<p�" ��d��<6D���B�《��wj��_B�	g�ҕ.3��$�ɐz�V�Rh�����q'�e���_���(�9� >��E�(�Rj�<��U���QCtT�GR�s5����<xS&�����&O(L⻰)�m�tr�r EY*5o!$�Q���2���쌒�(4�:i�WtD]�p�C4�r���T���Nl����W����� ߃F��as�����h10&�O��l�u��`�K	Ȱ[�|*�-��iP��H�����8Ij)��i�%�h��o�ͨN7�u�6��s�V=At?h�᷻��W��m�1x}xݕ�͹��^����!�C���s����g�I
EY�1�%Ӳj��L b��_���Z��vy8�Y��xy�ΗCw���~8�PW7{�<R��O>��2A��/*F~~�}�'��#�IR#��VW�]��)`> �*�����^mJ��"�^�^(P��2���j��O1x�~�Kh
����s��7LU��I����>_N�v��)<���c�[��;� ����@xtx�4�d������zJ퀭|2~��H�.�y-l���9�� /��#�{�? l`=����_�Ao,�Hu�R'�l�_��'��xg������TOLХ1�*e1%{x�>�e�N���raRIŐd�̥�NA�Rh�a����V�Mk�������㲞�Ej�X8�1 B������Iz��*AZ��N�f�{�%�'��i@[�E}(AF�#&z:�Y�Ф���,SX�q<�SQT���>ZJH��ꪙ_���[��諙Oum���ǠZN*_~��-̕(��i�b���ٶ�#�s��@#H$Ѷ���+�
������g�w����ה�<��݂Y��*�٧�3���ZMT(��*2h3J�eu\�)�)"��0�ľ��	����LQ�F��ڢg4B�E��q_�(��zBC��U���Ut*�p?�MHV������o��GU�h��c�IlL�I����h�rM�V�޺V[`�jp⛶�OEȈ���/ixQ�g�dٜ\M�NV�(� US+�,�C��~�m
dXm���ruzn�錺����*�x�k����wW���Þ�c�n?,4(����>'%!��^Ѹ�/Ս�VSY��J��F`eEz�a�C�Z��4��N���=J�G5&��ٰg��ر�Ț2�;~M⪔Q�x�e_/�/��Y������E���~5���
iⵙ�C"���5%@��cs��k��)b\#��n&/��r>[=6lR�i���xC @�NΪ����&���Gt��n�;#
��>,�lK$��,`��zܟM
oBT5pݚ�9Fa�S�`_y.��G�f����J�W�+Ԅ�%K�
�x��b����fr�{R83�&V~[��i� ������R,&v0�Y�� +SdO&M0���{.�89qM�2X�,�p��߂u��No��d\�����.�3!M��4��Z�`����M7 H�y�e��ki�'�_l���3�*��/�%��<!����eё2�㯡��/Ҳ�aO���]�Գ�K��&�"��2's���ͭ9\Y�y� �Ǐ�lX*Sl���g������YbU��#F�^Xu�����'�j�ؘ�Ԥ3F0
�Y\�JI8���af5��Ν���d��BF���y���2�)�=���At���ω�N$Ĝ�E����˫���S����*�+���m�(����q\Ř�	�ּ��?R�g��J�t"��yy�f#��A:�PƊ�ɂ�O�h���]ށ�Ⱦ�@X��\p��K�@�1����v�H%���UL�[��#��rz~�H�SQ3��g�KWJ�T5����j7'����x���I��p>@�(�eG��W��~����Lz#�ܵ��Uڌ��`�=Բh̤?[HW�%f��؁Se�@�q�x��J���<�d\��9�ޙ�?��%Πn� Q񵉍�a򍤐̗�ht�e�q�d+c�y�ZPd ���vu���;�����P���1~fc�#P<�%�E����U���W��`Q1$P*��$+|�,��vV�r�&KioVy�&���j���]Dݿl�k�|�N�����.c��b��<��M�e"IP�ãdo*X�J��+�.�T�w���ˤ�@�i�ب�mfzM�fq�j,����6�1##���`R
��T�mE�'���B~2V-f��#7��ҏ��Q�K��KՀgv�����ߤ�h�Dt�r���(Ĭ��0K��D��1�9�\��uޘ'*�ތA�)���W�v
skF���/5� �
�	�~��.�� �jb3� (Y���)1ſ��/����2�TI��K�z������x�NpE�Ӥ!���pf��*��[�C�}��#q?���6�]H�1�eH�׋��X;AƖ�o�a0,�J��z��Sc`2�P�J��^�4v8���Y|=�%���;���QM�;��E�ݿB��ϵ���^�',�UT�4Y�N=�'��K�
��S�bE.���b�X�<�M�Ƅ�&�z�m����p����P���!	O�g�P�]\b���0wx; ��V�屄�pi�}��>��@���Mε���H�ଉ*\7�>����}41���?%4�|K) o���yH��iJ��3,����U0�Bs�Y�2J��\����9i�i�̬4p8W-�(<����5��
���{�+�X�m���6͹���X�V2Qm��(�����"8F�G*�Q <�p�݁%P�=h��t�����[G�P�M�����kA�j�S�9V��Of�8(fї
�L��.���!x\�׎��׻W�,��߼A�����G��&޺�}%����I���ҷ�@Y��\�>�<�ҁT�nT[��}�ؗ)��I��ǒ���?c�8�������e�F���f�]�hBM�2Pmq�1Xm��Ѥ�>N�m Zbń
�y�.+:�(�8����O�K�CX΢!nM��?KtS�kr�3>�P9�K$���(��5�����t�9$�f*2&��m�tU�B��%��5�[�-aՐ���u��>�J��c$/�D9��%�"Dl��J*k<�M�ĩ���*�G;y����yC^����5噅�]xIRw`��9��\:����(MF�nF��L�3_=P�y܎{ 軥�v����O�C������I�B��`O�.6�	��s�P+�Ě�	=A��7���
x�����,�Mp����K��5�=��^*W�\�4����K��T��tL��K@���	�K�:����9@���}���=D$�t�p���@��H�����P�H����m�PB����T� 7[vΒ�����Uh��f����9�ľ�w��)Ji�4�/0%�#\��d�����h�!�&�;Kc%��J�SĔ��i�O��:/8��ZHD0�I���pґ��6���g{���b5C͛#~�*و�ph�2��-�VJ��s�A%O��*�#� �ߚ��Q;�':�����s��]���.��R�Pj��Q+��� N��CX{hp�<S�<'p*�&1��`_N�����*�*\;�G(�q��=L��> Lz)3�o�q�S!��t��ly���|4�q��{�,NR��9�n��6!ƚ�I�e�K��4�ˉft��_1:ʽ�R���O4m'R}?6���YM3� t"G����ޚw��v���P4��RaS4�T�]V�r�@�b�
 ��T6uf�:��3��rp�����ٙ��A�s�L��飴o:�6A(R*���e�V,��SV��@�0U�־�@]Y��Nd�����Dnh�{~�T�r�'��9s��so8�Gc��!�u�^U|�z�J��R�[���gҹ�
kro������ڎ����K����r�/�R�2 �Ĵw���O��|S����ZRo�|h�<X����5i��5����ʕ�\:��6�*�w�����x�;������@1�u�N��0Wc�mT�҈�?�g!.w��/�#�m��Re�*�m�`3���sC���8�I�t�5���Y��LJs�oŠ��u�PHx�;�W�2O#��8E�{�����Ea�	F��Ǥd&�?��d��u[��hٗ�#c�; n��t&���-�3��6[7���b]�,?:)�l~���� �H��+�l0U���
v'�t�
D�΂�'����V��in�2�Ed�����Lހ|�������SFa0X�l��#��m�'��\��g^]Ô��#���{��������x��������#�C��2[L-���l\��E�]��I[��\��(_`�i>����-���5���uBEF�:�"�:�߱u�F3~K�z݂�����"�|��g�|�4���2jwI��.�J0B"<����]�^y}fz��Sv�FXD#�OȦ���� þ �d棂u�թ���haS��d sjKI��[��$ТlO)�&�	m� T',�6��`d��R�B�K�pH q�-$���}�db�)��?do�X�����h,cVY��23"��\�i<o��`J@m�Q�̕Q�+;1�O����J�M����+¢�)]YL��ͬ��eA��b$9^��fR��1�+����u�UJ$�e�ܨ#�lT�%�L��8��B=n���?�H��:(aDы�����{ ֡?�˒Z�o�*���1�58F�6lI0iqsys�/�tx�Z;��
�V�*�oґ�͇�������o,��|v�Y�Q�ę�v��_��V�@随*�����|6y�8��'/�������"���[��B�q(�*�Y����Ÿ����vc	�۸#�Z4r�Otڽ�7����}Չs�H".Zw9�n�����#����H�ff��3~�"
^s�*��xr��6��y��6�{�$�q��v�ѹ^��Q���[�7�����%g+&t*@׬9�jc!	R��]t;^ Z���?q^o��K�������Y0�t7�w��|Q�YW���2���1J3�R�k޵��i�����K·���=�����E�U�`��g2Z�5%����PyJ�R�q��q�����/
M�nl-�f �������g������@���Ȯ�$���7[���OAr���X��b�.{-X1���jE��ڹn��B8n9�h��,��<�A�'�v��n���=�v��zș�+e'��UK�Y�U���q�����Ԣ44�f����p��d?���*G�	>�����ш4��{���YІ�A�"O��i\�P���cn��u3�������{d1�*O���k�T���)�JWk��t_�a�Ū��|-�&�_�|�wk��7����=6;Z���g7���>IU�6��Y�jh�zk��;��n=aCX0�5�6nQOL4��$�!��3 ��!4:�ha�YAO�ě}6_�<��e���zOO�R3���{��z�Яs��pE	\w�Ȝ<�=�<�	�'�ZJ����7y�5�ⱌ�:�~���Q���3���5�#PL�2���N�dڒ�~�BI2x����O����u�(�Sʊ��HؖH?sU����%�b� ��A��Dܴ<�*���Њk��`���`9��<A ����Q���I��yėcm�M����&��c����1��=���	Ő-�N*���}��4|U�SE��U��ݽ�W�-3*��B�i�-_k�!��#��:��.ETN*@9˷�@��uO�-a�.�F���"B��*��1]�'W+��vl@oo*����;��?-� ��@������|L��g`�=�x�]�9�)Y�hq����5��|S�B�ެ	NEf���V��us5��a�B|���a=��UT�����;�h����,ӎ� v'Q-�2_I��CN����O�H�-*�4�:�B��'3s܅i̍ҷV��C�7�ZP�ڳ��6�1��쿔)շ�%�!DG�ߐ&��0�%���~iJ!�8X��}��#	e�fvP:=\���VK����0C��(�u٢�e�c��ϟ88�ܶ��~W$�R�Os��m>';���>�[ h�W	Q�!����Ta,��ƛ���'���iB�ڻ�:qA	e<�A� �$a�z���Z���>f����&o�:���26�sN�4o�:7[�b�i���8qW6���S{�^�p$w*���f��~v2�n	2��"�~���3���~F�������C�W�(p=�oL][��gM!F�+� ����6���I}b���Sn�������C/��e��=\L�HPVѰ�a8FS/���S\4�H8�D�i5X�`�º������k��y����گٯ1������S�}��=d�h���M��3HJ~0����ך����U"��>������Z�:�z2z���Z'���&˩�iQ�5��؅$�!�i,���Y��3H� �n�ȴCk�L�H9����V�E�Xf��U?rC5�6<)��
B�g�8�w�>Xz�i�5w�"g�yB�ˎR�A��A�WD��9�3�z9|����v���n�f��ˋ�w�]�r�)?eV}� �+��00%�E��c�����5\J�-C𔿀���}B rm�bBt9�pcW ��Y��%���R�}��r�5Ƭ�}�s�[��)�h/�}��f3���-^��!AaHB����[=|]���t|[zjC/2�� Ocr}��N�"@��� 40�rH--���2�������0-�󞤼�Pi9q�)�}e���hN$R5G�����C6�Jp�k���db�թa�r8�Ei�����;O繡��B��s4!�&f�J�����Mm�&�Ar�6^#CZ���,���Uu��$��`j\�OV�^m���Q("~�=ݑ����GC�$V��J�4��?0�{��[]�����)6�mo��f�`�ek����������������I�Q����z�|��ur�KH�%��W"�]�q�;���#�c�Et�v��C�a};q'��n+�����#HSQ;�?ڧCd6�G�������-��}@|5������!����t�)ZfO�R��]�������,�{Bj�� ᭯/W/�>�(L�2_��ð����Y�K@W�=�2���ߒi�tZ�����WGn|�.m��K�������i�D��(��V�I���9q��]"H.kF�@sk/�,5a���%��%/�.�p���EpUBX?mni��*z�d�ە���j�<0�^{Hz��H��}Q��_�6���Kr�eB\!�|ٷ�H"Y�� �{"�D(*ft���\
�@�D]u����1�'�~p]����}�)8}�.��(��e�l�X6����j�}! Y���_��.Cn�4<��h �U4�"�G��5�X�����Z,����
J��*i�8,h҇&bTty`�� D[	��T�����)	Y�̃��A>� ���U�/c
�ZG΃�ry}R�5W/ yt�eÝM~���ɚ�
�v�@֙9o�7F�	7JW���2�?��3U�б��F_���o�U-VY����o�MUζz���H�<ٻ%��nD��Y��{_�Y��(�����]�H�Y�L��	�8���|�/F��#���:WY�= ��6�kK �¼;�%��6&�5��zb�K�4'�aeR���vE5����:��w��%쌈����n�	ۡ"��]�@�K��I*ȇ��m�92O���Q|Z'��O��� �YHU�]o�S��Ƣ-#�wm�3	Ep�!g�����2�?	�>����bkf5��*����~�����$�����Px�	�9���.�����\���"��\��3yDqſ����v�Xh�XU�+6޳�::����h�zvA�5Ee`>��qz������w������1��KC�u\�(�#=e���ZK�ok]���XB�l�Bkҍ��[{|0���m/�T����"k�/2Cݽ�R{��5D�8�>� ���� �ͥ�� B��R����'�xgU�l�m�H��B�N�ﺾ��ԭ^/[m�on����޷w f̙�Zų�钡�WƞV�7?Tr+��og�]�B[&�1��!x��\mlt��r�Zw�uK��CZ$ ҕ$	�((,I�l�\�M�a��U�3�����-��l:dЉ�ޒ ~�!�~�)�{^Dŭ�	�o��!�Ў��?"�Q-�I��6c��y2�*��DT���v��FK��zC2:qmP��I0�i���(;�T�+��ٜH��d�*��F>0�~��,�x�������V���rBJ�a\M�}Lj������/��U�����K-U�Y�JH�x�;�y. M��Ѐ��6M ��*eeT�Ƥ+����@�N-},�y4�ajA��e[�!=�n�F���p��&��8��j�+������j�����z2r�?{zݑ�v���+U�m��o$��Fz,rK�O`1��$S��z*B���i�0��rx��j4e@K�:Hg��][����u���q$�Wy�P�K�-��rv�y�g�c|�%�-q^S�f~��Y�_'(G�����
1�W����%e��XPjTy���i�&�x\���b�����#9�-l�Hf.d�؂z�0�2(��b�8p}+�!K��Ψ/!|~�����A�t�:;�P�_������C�,���H񁍗�K��j���UqDP+�κ�/�����*
uf���S��/פ����ƇO���G1yE��Y�j.�Ϛ\� � �����H����I��P���Cv���F�q��x/�d;c�������d�a��x�I=A�(Sgz��zk��Z��j��7�j��%�ϓ[�P-�V�n0v_��rZ<rS�b`R�'�oq�㽽� �$��C�WdX<�d��A�v��_�a�nV
p�y�c��㞟��"�@Vu8(˱�6�NI��b�-'�ew��*�ː� �Ϡbx,(�Vr��<��'Hq2/�Ə"H����VL/��||/7^�%�%��5|~t������Ep�) �qI�4��*����wkxQ��i�a�6�&���x�d���v��E<�s�^^�U�yʸ���R~Fx��Z�';\��|HŌA���e-�L4�Ci �<"w�mI��.�SH��9l5�5���g�1k�R���"����?�P�'�d�T����IG[��~�K:.��63�X�85:}��I6dg�m���?h��c�0���(M�%��`�JM���f��f�*y�� ���Q��w8�H�3C�wz8�v�j
uOj5Q6� �QK�ה�ʌ}�P	�[��ag�N��[%���93BV�;����b�^�x<G���ω�R�M<�II�u���͗�U�t>���{`�@�F��K'-�I�Jĕ�/�o�(�Ƃ^��vD���C�������Q�~����Nc7�k�B�j��Kp/cw־��[�q���H�T��QC�&6C5�۳�xX�]=���Ϡ��&66_�C���	�8i�����D���g<՛��$��^��[7yR���*U(/S�,��K�Syz������<M�_�t���!˒6��6=�]���
�0`p�����?��G9ggh6�H�">��Jn�+٦[bAL|ɉ�T�CL�:K����롾�%��+xg��%���n��3�7�F�D߉�1���'�Gzft-�����6�,R-^�����}ݺ߮@�+��3r*'���X�Wq"J��h�Zג���F���/�ۑ�"^����Hw��>����& ����'������G�΍�n���wuj�|[�ҕ]������K���"٠��Õ��@G����M C�G��<�C��lY�S���S�x]�x�/�W?���'t%ۤ?U#��)�*q��o�M��'�`zЏ��R�v:��N?E��	�:�f�jK��3��ל}��-�}	���.ڇ����y����5^��7eF�9)��`yr��ZJ��c�qB�ӣA�$�a�Szk^��͔sG23x�9��y�B���T���}�
���Yä�&X�V�*�`�H��Z��Nl٧�"$���͇A����s)�q�@a@�����K��yG%�&�W��!��Y����8><��Z��͂D/x�<��\9=��o̭�L���TPo���x�1a��G��FSz�.W��D�7zbE�sՔo[E��u$-�k�<�B��/�²�ߠ��i�;�5A���σ~�����āQ'R:����avw�>�T>Q���Ø�<�=�١b�!J^����.|B.M׍w�ld]b��҈$���]��%O�I}�ٓK�]d���Y^(�8�q�~f���.#�ٷ}���_�'܊9l��s�g9tMω�, 2�4��8��L{��r�d����h�4u�b�J�?�7��7�+��1����j��q-�գ�F:�.>3A�[t��A}�3{/��P\����ϑ�
g���q��ʣd)�?�w��s�V<������m˥��m�3Zn�!��5V<��u#��y��B-[KY�O��T����q5,�\�}�%�4����$��%��N��l�'���v�]����1Nrj�è��2��רB�����B<�0�8z	�L�X����೪���C�Z���Q5S��&2�S�D���\`�Kbd�HY��赸�^3�������
�_TNs�YAA�r��%0����?���� T#��l�^�?�sӫ?��;&��7g:!fსѽ�T��\he��
}�R(��n� �k᤽�B��h�tc��0�\4�~�H �
U�Q4-|���Fv�;�%%Z)�X�;S�n��t3I��wg-�7����^�n:�g�̲��٭��cC�&?WPq+n��	����)(Ԕ�
��-�6K�P�kщ*0y���m�GP���� Zc�S�%|��0���k����������ȵc�L�W,ub���4��ځ��/	�Wfm#��+V�[�M`��W4�}1�ؒ~)�!G�U-��M� /�`�0�Q�%�M��r�p0q*��eޑˑo�#�ʜ+��SZo������C��	�E�x�#~�:�C�������}��l��j�(�Qja,I�����M��K3��A4ue��^>F�N1���T��V����+�5��+��&�F`�@���g�V��m$;��0�}mJ�<��v?���/E�Ch%�v;�^�lK�Y�Y�;�3p!Q���]:�Τ�j����E�T� qV6�$M�R�Ѷx�;��]���Uz<�xQי�1KX��g��<"��
V���.�M��#̼�3�������Ҍ��يu���Cjt�G�)��� ��L̋D�#�qד�r��jǙׁ�o�h^m��I��;�{�?uR!'�/ƣ��y.�k������ nO?�ď�Y��K���������B֢�`:Nq��a�&�D�cr3�~�SL%�9�J�N�U��S�ط2���DIĜ=I9���p3&7m�hp�p܁OB�x�u���;,������_.�I�D�R�e,)K�;Z�1���{���'w����?_GEF��¼y�q�nʮ,�P��m��/mR=}\W���A��{'���&�g�o�-�E�d>�&����*c�K��$(H��v�hz����h;�Պ��pv4��iͨ�b���`~#�4��^�;�h]�P�������J�q��F{Z�A���s���18P�/{��HM���%����0I���q#����H��Iٽ�<�' ��!^N͛P��}{&�R��A	�=ɯ2&(�S?�>��&W��V�f���3��<,�Z�-�i�lY��ը�y�f��ED��	8I��r��\�*�[f�_fT�{��[k���}%j�U�_�-3���L2؛�G�]�F�ĺ�-.�mh�jIlūe��&�|��?yx���0j5t�_�c���G/����"�[�;%\
����N3=��|������"x��/#�H�EI�c��/j�%��g�����1M�l�#M�R��7Ծ��w�����=���T�����a��l`Y��͈�d�f �{�]��]��T% �4h3���rt<E'��7��("�@���./�v���'l�+��O�3����|�>MwJ��A
��)��ke�b�|�H️�S���K�ueB ���W��N$3�޲����l�<���h���9b`�(��Sa�@[
�j9s�7�m�R~���W�" �9�p
�0�++�����/�|��|lX���ı����k�� ��9��e�x�N*��` И�����}w���,R��:���Yݫ�wC^z[��dfBV��Ȑs�p�2�h��:2����D�U�����yp�|���4�i�p��4��|߀ֵ�4���o8�����>+��eJ��XQ�ǒ���zM��Y
l56D=�H�X|�]:��3��&�ۚ��t'C��d��bݾ蛏�J0�vM+C��aư�-4�NU�`;��ޛ��w\W�� �����&�f��Gt�~ԚÐ��LB�Q�PW2Kr{M=�P�5s�(��(�8H@��}���pN��d4���H�*�|E�Ǎp�rUH:�_	A�<r��!����+$@(��,���"���㒗f�`��P��;�{^ԕD�
x��}K9J��[2}���k �
�mg�%�z~YW��w�_�&o��R��h�1��=�8p`�~��3(q���ذ�;��^��й�܀Č-���}a؉c�h�[��0��V�N[T5p?6rڭJ{�S�~
���v�B"��c���p%A��k���J;�}��L�PI�_�s�J�5J�N`o��!���[>�&�z@���tq�Q&�x��EVh���M蔧�Wi_,i9�^(��G*U�^��ئ��������a3�sX{_�M�ÖY�m���"�Ԟ�DCG	���`h1T_XNݓC��	�ȁ�P�AI@>3��э�/�z�t��k>Uu�������DL���6��eXHK��:�g�3.������oqWn�i���N��(u���ɹ�:�y��u�}����Lg!}<�LQL�G��.�5F����B�C���O&[�x�jd��U����!e�rc�V�N�����b����M�z�ӆ�u����nHpl�d�(�xiUyo��ݬRh���ŀ������߹�R~�쨷/��o��D�>�M�7J<�A��?CIȍ%��Q�=JM���y�^o�������#�Ub�#�������=-�e�VA �4QPA.���o0�H-Fx��X�+�-!�����C1�ۖ�mL�m���f|iS���`�Z�z��X�n}W��ْ����I���H��r+G�K�EkQ=�/�R��y)�;�_?���}!�u����b��r֒c/ȏ�W��
���B��8�EiC���3c=x��5����������1��W�L�@i�R�k!�rb9��|�l�׷��%��ր=�Ԏ� �UT���ж��U��X��PHI2UF��V>D&�"����K*��e�	��	�~��X��Z��_;.x\rKQZN��ǂ6����k�����6�&�Ida�[�T)}��sװ|@vI�d*ʟk��G(8����'�
d!snlz�F�M�(I�RIS0���LN�Z�� �Ҕ�Z���k��μ�?H�
����;!��x��E>i� $�QlD�Hb~C�]�i4WA>���E���KY�R����"�:�?`�&�VF�h-~�B��0��v�X��k�/5��=Jԟ�q�R��t�;��N'R��ORv��3�G4���������	��vßs�7v@B�Hu���>���a.mʗr5�kҙO�n5�:�{��A�����jb7��$v�Ŧ�����{s])�;g���ٯ�>��NB$�S<����s��l� x�g�/\:�d�E��ބ�w�Nތ
G���I��p�U��{,��ct�ۑ�C���߳�����JV^ �.v�i��,������ǎ��Z�ܥ�'���(ްM�b�Hʬ�h5!�������c����yG4.�����y�׾�8B���o�!�O^�]�z�f?f�����4�K����hԕ�衮I��t�윹x+g�6�*����$N�2N�01J V�`ɨ��V� 8����xؐи�v�]����J���G�Bw�}=�!�F�L�b�߰J����%�\N�"��g��ej�Y�C��1tq�q���m�����xc�3O8jq'����=$6��WwSS����yS��V�D�nu�{(�����{�01^֙Q�nY�''���';�'*75�9��W�[�60�w\N7�1�U�ޔ��v׈������`ƺ�'}��� �t&)Y��[�y��p�VGdKc���.y��(2��y,��
��i�����,�/d��{���'Fh���&̥��'34��É����(.�x����[p�QV�ƪL���&����ɉ�d؎�Rj�g�^�����^ŅTTE�/77��yZ,$̺G�X�>�BO���?�p���ED�ߧ�2N��vvf��ƄwT�)UvBG����+p9ܓ7�v�}G�����_n�
hL$O������yƊ!���:�"�ΞtJ#E΍Ĳ������OV���aԷ�I�"v�jhKQ pW�>)$"��$��-�8�:��R�d��77���\���.>����a3�>�K��9V�ka��A�_;����5˯f97��'"۔�J_r)��	@[:���5���l|�=r��>���c��Dl��lu�]:�9o#�~�g+�)G�w���Z�L�;�0ݭ����K	���t�$�n,��j'<������=1�rzW��ŢS"4~{������s�Z7^.����B`ěg�O���hA N/�@H�mu��ڰ�A�o;Qz	�qE��i�\J���$~���
w� ���3yX辅�9�bv0�BNE^��R8�U�HB��� �X'861�@*Z����%id�wg-S�ș��)2z�/�q�Focw\�zƩ:��'يz���G��}%g���֘����PI���gA��K�% &��#�H=��] T�v`�q��w���,f	C+d$��Mrē9�f�;�3-��V�T�(�'�)�o?nD�����ۤ��H ��}�Y���4��|z@\�qZ�f���;NF6D#�c7�5��y`�͔X`->�͓zN�c���s��G���RB��mC%�Z���b�\�O���δڅx�a��Be�9�����}M(��,������������gc�-��ߠ���t�?.�)����|ע7{lNJ����|gX�����O9�K�j����9�e@_:F��l��ѝ�5���O�h�W]�Q��
�ċ��wV1��H��9�3�=�	�۷��MA]��G@�֊��p�:Z�$	2�\����'"LLhe��r)�\�}��\P,gI!�H1h�sR�z�{/��59p�~��P֊ؘ������t,��
_�e�΁P��(�6;γ����q�Jq�j!�{��۶H�>'�h��z��u9-Ț��8:�`�� *�Έ����z0����<��Q0�Q���BXC�$���r�w͈�uTa���mf�k��V�h������sv6�Q�U!)����c�[�-Dj��͓��J�^�Cđ�����M����3Y�p4\)qܭ�,\��R ��>�(�K5<��td�b+�U`�^���c��f ��NwWWv��R�Y��VЌ���nZ��s�0c`�-�޼�k1C��I�I�YH��s�܆WKSv�+z���&	�47��s��ŭWM�]��<F�!��;�ȦbC��R�!QcDQ�Gq�[���-f����P[}�g���Y˚d�
�2�,�uj������jmc���k����� 4pu(�`�� a��U�YB�	ŝ"*۫���R���
���^�z�T��я�y$JE��F�v��%�8�)��Ǆr�Y���_��6��h5FeA;O���eEC���i��a�McXKށ���:"#� YS���ݢ�P�4E�iO�;o�L��w�4�TT�M�~�(m�6�T�� ��gr^Y��J�-���E�#��[�.���|ߗq��ks�����SK���V�L��S�ߞ���d���������I>�0;Yd<m��Tl���n��FNS��\��U��K�i�a){��=���Dkۨr��I��@/ރXٙ��� ��,#�!(�#)�1qO��Fu֕b�|goO\�V*�K����إ�$�]�r����3tdнӰ)��Ơ$��m	��YK|a''u|�K�m�__^��YcZ#��7B?�`�5�p�o���1��sXG���/�@�1�4̬�	���1[2��Pc>(�K}a�~m ��ł�mTȗ��;�}x�+��6��A��Ai���&�\�QK�Ȗ��8M��/����P �"�^'� �~�Ҧ�Zٯ5qW��?�jGk�AA܆�=Uzv�^�kN����=^�pͤ�lN�TO�z��e7yxf�=�����x���m���n�7@H��џipZ�u&�7/�
�]/K�p8�v+��3���yV��ŵ�h�@T�9�\�3��Ҋ�V�߹��/O]�Ef��>:a�7���0J�� ���t����]���(�nW�늰�q��oT�rR�W�)p �|jf4��jZ�Y�je
=f_�R�2G�Īf1)�/R��|�F�Z��g�l���D2�O;;IE��-��ޒ�e�_V��i��fħ�A?�c���D��"����3��O7�,���S*`l]���J�K����lȮ��蘃?�Y\��t����}��Y�bY�ގ0�
Z��*��I���'�S�"8�늝�!��N�K�n6�k������I;9	����r>��O�d���"�"�A�WO8eL��Gr}�H��TOY�� P.1�+�k7�#R�z�3���q�Q�DQ:��M�pB��o7�y�D8&Ҷ�:�8/Vր�g��&�1{ΰ�`���������.�v�d:����})�E�cIn�'�Ê�C�7�uң��b�}n/�.��Ǽ$}�Bys�����3�L[!i8Jz����-��x^~fP���6Hr����Wk�"9�銃U��Yڏ���gT���G���p#��:��8 �WI��{f 4�|L��<of��
2l�[��汴���"*5G�v7Ѥ�M���YC�r��C��q��Ҷe7��
�W���v;���&���~�u_�x��H�v�'�f��w���Uڪ 0��,��'��oN{>w�#+���'�_s��[�\G]�.���&�m�z�"�� >7}���)o�M��p�]�����}^��J Z�=?�&�bj�<C:9@o��I�	/�o+�|�6FA�B3J��C��O�Ҵ�=K�/6+�Řg�$Y$J����0�)<�5���l�&��Ht1�Q���)lh��������K��:��:dл/>1~�lm��Sw�Nj�u������ҹM��^�ᠭL��/���,������NYt��Y�V���ô%�Z����A[T}x�'�1��;б�œ�����>W16�{�G�^0�d��u�Á%������w�x[9a�z�#��0�`�0�I�ʣ�l����l�KdI���w����Q�씅�_!�_�{Z���qO��|�M=��?�]���kك�uM1�OF�Ge�A�p�r+c�QK����a�Xh����	�-7�ai"}.�JtYR%���mh���f ~���yn2�������EL��f�wX~%D�a+],��#Ih�AT��qg���.-�;���~!PCRsn��(h���eMv���8�D9���0�!Z� ��F�rff{ӊ������j��֛6�����W�q����v�x���������Y��fb���.��V�\�4��)Ü�v��r�ٗ
��!,�)%5�4B�O���(�(*��Ӽ������	ƭ�>%L�u��>|�B���\(�,�tr[aF���o66� �d�0XhD@Ѿu>����Bk-V�����4x���v��S� ��ѽ+���58G�>�S׀�+yBHü����]�[��[�|��!�n��Z�q2����v�n�W@�ͪ��_�E�S�n�c-���j�g���J�Ѧ�P�)��ޑ�wbZ��l�铇�K<t��k{�j��k�V��nB��5�hچ�ul�!������O��o�	A�!����.[�u;�r�h6� ��b4��G��ߡ�A�@Ę�",�X\
iV͸��#�$?o�ȑ���Y�Q�n��B'lPEiq��6�7������	�٫�=Fc�K,��.�&[�d��b ԯ�2������ͩs˙����H�O� ���,�k��J�����oȥ������l{ks�g_��i,���m�����0�K��X�&y�u��"�Nl�y�2�o�p&؆j�@d��C[2P�Sj���E���[�;��B-�,����J�E�Jy��X_]�$�����c{������?�-R�Vq';�f�,��z������O��#a��j!�Q���7Κ��*����&�s`L��.�j��_~���?�_��n�N����J�����U�ht��y2�O1[�=㚿��2zI�����p!�3���h�}��2'������CAwZ�={��t���� r��S��`�%j���sA�t�(��r�U����sDg�+G��+'��%�Cq<�!@Dǭ�q�Z-����oӤ��,�DQ'��h�MB��i�Th�A�.+���wrDx����o��k�_%ӕ/��� \��@ Y���[�$��������v%���12�Z��O�#:z��f�G�^�yφ]�����T�گ�E3�� 	V�g()3�T?_�����e�{�a����CEM����@��`�=di��h�(��>��ȥ}��V{Y���}�͖?�"v��E�:��Jg��l�����6SB���X�ski);�L���=����@�(q+��ϛ(��>��Y/����=��d�V�*v���%N&k�� �S�c�6!����^{Ӹ`2Б�t�1�$��!���x��i���+����9�\�I1�-����T��Q��#?�uo��r�V��4(ERS�y%�7N��o/g'�ϕN-!��)���xc��9���3O���KM0���������s�۳���M�9��v��� jM��2�� z�O*�lQ 4��>��&������3���:�
�[�/���W�O��]�������
u|aNM@<i��h��s��@"B���e)�x)���7�Y
�"i`���Χ[�ȸͩ ����!�@�"�
!����5�		�{oC�\~ڧ�ĉ|��S��[3�^��0O�K��
i��kG���T��L�{=ˇ���	���K�N��9���Iz���Z]0��/��ťs�4�����'R�+j����sla���B+B�U%����H�����3��'6+9Ý��� ������.�W�������
��y1 ���^<�y�cnLV��Y�&��u00�
����l�����W�(&pm&Ŋ�"�� $|������'O�i'�ܿ�	�L�6��K�'�[�#��u(���u3�[a,CH��4ʳ��	s	�O��^o,���\�`Ƒ�W�%����%5��_ye�l[�z��_(��u�E)�ۄ2��jt��߇Q����m���b��6v�_���䞣��>kؐQ�l�H:����^&Y�.R�{�����l <���}Mq��/H�i��m��s���1l����b��eNP��/adW|n�b�@2C����r���6�J�3IS"P_��HG�E�4�}��j��Į���K��C
!&ỂH��hT��>Nc��Ǹ�gi�
��p��M���_��!���%�
ƴD� A�[l�T��^a�m��p�R��K���ʼ�b�{hMJ��Mc:�7��ɄA����sp;�ݲ����Ȟ.J���z�/�2��oo�-�Q
��0�MH@�x	��y�7j���ׄ��(�M����z�� �K��~R��Z/�O	1�`��|��a�3�W�xC칱Q�+$����oz��\BO%A+3�¢X���k5��F�ׂͨ�	QԞ֍�D��?g_XzM�_�<���@L��lƤVq�*�����o��_��KD����.t�m:����9	�t�c��t��u4�Tɺ#���Z~�|9���Z:�����Q�&��X+%&w�mc�����ї��������渖�lRI���h^���f�ɿIڷ$:M@U3����h�@��2�"�����[E"ddc��]�7K8�u�pJC�DE�u�I��!|ٟ�j?��1��!"*g8������A����GN!crx�J}�W�<|�<Y��]��d#�V
&W5m���g/���_Kr�T�%�͊�{>y��`*?6"Ϡ�+Z'T�뢦vtV���~H��AS�p�7����\X�m
�������,���e/���+\Tڣ8aFA�3�6���-���U%;��t����g��!�$�nG����|����r>��4������'�L��eP52�XDc�����e�WT{�:�Y#y�	��J�N6����m��ulT���T$gܝyR�V؆#�����\aF� h�{ �H۠�V�� ����m�'����I����n�����AC	$�!�{���,�m���v�I����;�hD���F�N���5��f
��X��P޸�K)��)�����9[{�L�å2�1m�[k�D�/� A���W�n�ͳ�L��+�yr�0��E A$���YX�*w���zf.�����w>����X�%Hm�`��-2�I�G��I_�0?
��j�N�A�\El�Z�3�8�[�V�u���0]�X�����!v�{�F�w����"6��|P[���u�U��mu�	�/~�)�� %Ӿ�8�$zalә�J��,�o�������	�|ן�}��:T3!���!�A�Qv��p��z�n��?|�|�N6���wIuu���e<
���b�+r;���]U�i�N^��q|�q�F�^�/z-+2o~��O�2���i-�^[	�|H��8�9< �TsS�����v��J��������
oӮ�g�/����fvP��l �w9Vi9��� L$�%�K�iF�>OH���`�pVz�t�:���b���I�Vh�������	*�`����k�c��U`L2�� �M�K�ጫ*��-7�TȠ������{~�W��	�ȅ��ɖ�S���I�#�,+���e���
��ek`:=��i2��Nh=��T�L_sз�����+ݸ�1�-�%���A��>$�e�0MiW�'��c|��aa!y㽝	ݕEg׼�zX₢||o\Y#�8�nOZ������U�W��o�Ŋ!.3���	,�a#⩇�a���)��,;���]�8�z�w����6˓f�Z�S�t��TOy��J��f�ҏ=����Ǐ�+^A]}���LdA|��� ������!9�ܦ��#����#:hz��Q�yNc:?�Ϫ�D (,�g؉6���Y_m�W��91��/�@&��.�LRp��4�:A����<�ao׉���H����i�|r��-Z��p�w�럛��w�S��1���M���QJ�p��Հ�İe�U�>�H��Ey
V	zk�k/�XX�	~a1[p=�h�&�g��`��.96����E��v���3Z��f)��bR�[�Qq,�at�ͼ��1�׺� MG��B{+!9N0��͂Ŕ��ck�7_���U��m��g)�YC�iOH��D���a��DLć^�_�m<y�~�^m~iJ��<�5��� �p�"+^s��v�.�QB���F����ѝo��7��B��4�%?xM�NP�3��V�a2/�������Zt��U�FcD�xFĥ��;�f�	�v� ���ްU��������D���䦸5;�V�
NgJ�\�:�Y��0\�fixo��r��ڸ��`[���F�eX}�����:��
`���b?�}��M��F��]f�SO��cÜ6{��b)��s_�cV**S����P�;��2�_9~�.���h��Ћ@۟fɓ�B|4����4�2�l��+�T�<DM�r��&�p�)���Fμ�qt)��f��k1����i8���o�5�_�L�G	{"���dY5�w��q�'�1S�K�TZ�J�kh�J�r�qӫ���,����b7�8!I�Dɮ:���:[ ����!ˈ��n9�:3��T��3v�E�g`e�j��&e�BZ�ʀi-E��T��#�m�JX�w�$�fgm0�m�y�7���CO{�=��g�E���Lwp|�^��'���cv�Q;,%�Y��>xZ��ȵw} ת��6�� 5
>��dۊ�>,��:h�f;���G>W􂠮��'�[9�<�'H�>Ƶ��u���q���9w]�&Ä�_����!��j��}�8�҈�.�pX=pc�~���o�$�%���<S���ȅ{��������hl�hr��m�Pr0^�DL�O�(~����uJ�':p2_Y@�BR�g�B�B]� L8�� }����+(��}�@I{Nb1y��%�����Z��-�E��юݑqu�}��q"r"�������afe���V���{�X���J��1�]��G���r���Y��k.S�)k�B�T���`aΉԙ[ᅬD��"�L��=U��W=�H"��7(��l���cDKkK��8v�� ��_�5=���*�.�1�N�ዩ�MHl�5���g���Z�S ��O��o�͙�5�d;���`�y���Y+zS�`�|m�i��p6 w���NI,Jz��v�� ��y������x�0!UNF�%>��ʢ��E|���~�ʅ��>F�TpƋ���=� �cm�\R\s��J��k(�X�c`���ukp:';�a`@������7v��wC��B�Cb�g�Q�z83%�ԕW�O��K�g�:,�8��Õ�r �x86�,y�Tr(k�UU^-�
ԭG��'.7��#Km�~�Ē��k)�^��B@�6Ta�h������TS.,S4U<i�C�i�<�#?@�ž��� `Q�{7��>��>��}j� 4�9.�"a���&��!p��=��ye@��%�^Vs R��Á�ȴ�S�$~_va�HM��5.�q���췮��'=���ё��v�1�I�:kq-�&��uʁ�fՉH���%���w��{wZ��q
W��;!���]ސ�e/?��@��3�����rN�%��X���yf�B�Q|��J���[ѹ0ۺ��9YO��6��l�e|ס��2���9�����c�=�Ar'T�Re2�������#p��!T�PF�kz>`�w�BM���T�\�Rh(gG�Þ�#K!��"�%O˕�1�@¦��Y��S��큒��{����L����s���7�ΰ��f�;M�1q�$�0���+�W�`�!��V�p�M���&s�,�:20��^��*����-1i�B�j%-� ǽ��R^X�c޹8�m��]��>�2���,�g�VXb�4)��9��*��R�(���4a�+�m�m��wO�F��7I����`�e@��]/Oi;��A�I���`�h��?D�A�t_�̺���v���
?���//�64��[�Z|�NM0�U�m�z��SZ�!�2?@@�p��:\�}d�ţ\�z�=ɟ�g��=�x'�VbI������h�Mv��b��l�5�,b����s��|,����/�۵R	�ø��.�*s9���k��%de�nN���QIm��g6�`&[��ƃ%��K�'��T��>�mE翅��X���VZZ 4c�hW�#��pyn�R�ڲX�*DyL1�UQ'��wx�0�K�W��'mvT������D�!!�U8q�<��y���m��t�3ACj?<������0�_���3ZZ�5����������X��%/_I�R�^{�C���Z�=�I$��i��^�г&��+J���1�g'�7q�>����ou�y�M�H�g�<뷉�+�;���n�5�@�D`to��pڭ��hR�5D�|E*if`����lv �=0����J'��@��݄�Xd�w�K��Ķ'b����ȴ:Jq�r$)�*�_�h)o�k(�5�f�F'u��e�KZNS����hs)�M��ĸ7|P؃�Չ�xݵ�M�o� ^�����E��G�����A��#h>�*�,�w|�8��8�L��#���'LY"��C����:ڞv� "��(y�~���wI��9��ZX�Y�J� 2+i��Zm?�`�֞�tɩ�������I�v-�;sѧ�y�<
��8kY�Y*ۍ���~�FƎb�i�$�Cs�w���!�,e%B4<�(A������ ̀��0� �|#�k�%��ή��r���"����J�B��WƜ�!Ŧl3"v�b?H��^���mc�
��٤��(=m�A��L_My��f,�[}��-By�c}X�����0yUTaD爍�*j���� ��}��ss ��í���Q!^~h�c:�X��v�|/�Q/c�]ky>0M7���J>\v4J�O�
�>�*\��U��/��i4���� d|��~�z�_���u ��,g�~۶L��F��NGl)6�i!Ք}����r�ܗ�_���j{��#I���|��&M)艟��%s\7{����c�f4�4�
�����_�1�ߦ�e&(&$��^]'	�f��Z� �V���_�ȧ�����ZU3,ո���_��s=�Y��������7|��+�q4<��%� j��#�ېl��Z6�fǟ��}�_�-9c����h�/_��G0�F��+J!�y��;6 �����Kc6��ɩ�_OU���ݶs(���@lӽ �	#��Ȣ�ɾ��T�j���ߴ,��r|v��O��Z}Lb)�>��W�Wv8m$�P��F��!�*��٧-)_2���s��Ң�f�!�c���a �9�1�c�
3xP�>��������9t&n�U�\��i��XN�cb����@[؀�ה\�.��91�Wnn�9���1�d�~:�zK���o�#�s�T��(�K�)�M6�����p��H�	���
�6i�U��\I����׻܋���k���f����*!���S[�O�ʹ��/���P�nM��f��bF�l�͙�ظ�'=,,������.4�Xʒ͙����<'�>�vZ�W��45�l39��~c�]��L6�����2Ǎ
�f�iX�]2��^�=�;�GF���@��]��R�*m6geu�;�Go�o�L�<�����QM@k^~��R�� "�}p�����Vs,��_5a&5�a�Iϙž���W�Ⱦ�<�լ/
UNk�7'O����[����H�BՇ�2�W�\�� f��Ԫ�L09�W�UgV	7�k����]�!r�@	C`�%��[�l=����*j,\�Q�ʵ ���mr8���Uan&4[YDE�?컴���d2��+���2"�R>b�Q�o�j� �u\{�OY�]���|���ͭ)T��cx�Қ���G�?NC�� ��ۻ;�9D}H�֬�[j��*�"������M��v+�&K,�=��f�~���� ������6W�K&����_@��hX�>���j�F �!S�%,ص1;�Q��[���"������mx����z=�dUR�f������P�aje���*X ��K�ؘ�s5rb�����k}�E�|�v�;�
���x�&P���1���I@��˼b�I����'`�ɼ�bS��,U*!'2!���R��f|�����d7J����i����fǊ��bn�Ӧ�����E��% �6iE�m�U�R��m�Yޘ#��;2O��7:nv��������*�� G�^zd���0�+�im��Z�/(0tV�d��5�^8Qn��ڃl��cu���ԉG��Њ=���@+�����?�E�s�r�.�oQ�w�%f>yroP�x{�Q^�eA�#B��0P�Ln!@y����a+�G�ag�r�/r`�H�:���W�\.�E��f��-�x*�q��fj)}��;Z�9r��id�Ke{lK�42D�O��q;�)1��2��ʄۘ)�sPV�,�#����"�8�S��9~�:���f��FgZ��[�/s�X�ѧM68�?�C�yδvs�6�Y� ���8^��^���zlu�춓�m��p�#�H���"E䔶�N$HcvK���r����[��I�)6PTf�Yj�P���3}��&��>ݷ�o؉}�A>�oف[O����AP����U���;�����_������"����&o�ڊ�`�*j���(1)����k�:���D�d�.���,z��p��Me����&hwMZEL�U����ɫߝ�*.ϦΏ��ݭ
�vaY/���@� }f����J�r�r����0�/�b�Wk��$ā�A$�-3vi9�d��>=И�"���-��(�R/Xg�R��F^����=���|j`T�{���襧K-�\7�[?澂�Ti[~�ɕ.�Dj���]�e41�H&{n��+
ܧ$$��m�9A�IUf4��$~�rۏ���b�q�=r$OuՔv��R�U��)�}Rɵ�_�����x,����t��2���S{�`����:P����{������Л�5��LbGp��(�mH�K�Y����6�������=z�|�?T�f����[���bZ%�kQY"�J��7ϫn��F���ȓ%n��Y%~��Α��#Ѽ�y���t�d�}bp6�F2��ߙ/̝��r>~K��v����B������s*%�ظx;�b��Z����x�:�r��EH =���.����3U ƛ`���2NN��U�W�AY������:�ͭ1,Lm.~�#C1m���5:]n�8�6x�@�)�o���,�(�hϨŐ嶞

�ifvT
�Rt��H#����X��@�[��q�i���gwP��EA"	OM�g|ο,�."m��9���K� ��B\�N��{��%&+��|��ς"�֓�}2��l K>��al�ϛ���:Q�Rk��t�i�l�{�3l��X-�bW��ː=��������n~��LG�6 F�&�e�8��h:	���� ���sS)lc�������G�⌌݉��|��kAET9�(@p�����^��I3h{+&��-����ˀ���V?�s�f����'������ͬL}!�=��@L$��QK�Ri�%���Xb}:��IJq[��?�������4�ɝP��%;c�GX��JSF�,Z�α�����_2'$�7��qӻ�(���5��dZ��Fls�m�u�gF�l;	���Vu��Dp	�jl�m$$|2k�D�t����&������aw `BA��IC�ވ��3��D˺\�w�����C��<�4�cF9s50g�(�6쀽���i9��yu_�曄Ð��"+���H֐2�4WϢ�6�V�SYC��>;`~�#qo�~oJ�������1g�iM��0u8*��%նc��Q�}�D4?P�14��>�;-=���m; ����f-��'��$r�L WJn���_���=Qv�f����
[���=E���<�
�Ovg����)� �n<��k[D�\8����<��.��na�3C��r��:��k� C:��v� ���y�\TM0�lpE��{#�GGL����vo�X5� �:�.��t�����c��?�N��Q��I��ޗFU��]�kk2��1NiC1��'c��mZ൥��k�7w���B_������G^a_� ��߱�q��LQv�
ƪz1Ih���<1�=�8���q�P���R��������Aƅ�4%�Hʤ����bx����+��F�j�<5��d��ؤ�'ߵ��x3f����#=2�J�j�}*'|#Ĺ;�ݳ��S��c"vb���tHC�3	R�<+
��,�-�u�?��O�����uP�ͧK�LD��2bm����O�9�ڥ	�Zw�F�7�9(Q��N��<l�j$.�f@G)
�{��թJ��a�H�T$���1��
U����o�H� ^�E	�y�>cL0ڇ�`��R,/���^o���M��,c��3�V��3GV�8T���\���o����f�i�`u��@���c5��H4̠L&�i��my/�/jv�=!/V8
6NP@aƿd���yսa�#b���0�΃L*y�08�797h_~��m>\Z��C��M����ȋ0^�/���.A{��:���k�i_���mj:��D�YC=�);cl\�-���S��Q�W7����O~��-�>��>����$`vY���ߞ>[������)|��{BtT<1��2q�$	�S�������k/�+7��6`��VR��1�#��K5
t�O��QoiL�a�)�&h�/��d_k�"�j� ����-0��n�Ff�%`�ݴ)$K����ȰX����
6��n=xv�
O��|�m�N!+��win*��q��5>��$%#�t]&Oʦ������n]߄�����9�7H���K��?���;��5�C�D�Ԝ���b�P"C���t��7���/�wB�5�KS�c�7���I�܋�� Câ��	x�y�Y%�щ��x$����t��*����VO�t.l�S�?���sA�L��淵�No�!%�j��՜�Y��n1�
����	':�wDC>��g��}�CW,�ʵ��s$�"o���)tC�)E�n�3���X!�u/�q��"#��B:�_<�W��� ��1�ZW�#I_����C�m,���UL�Ƚ۸#�|�w�����~�d0ԛ5k��o�3 ,o1:�b�t����L\N�dmķ�#lO�QR=��H7�7�u���.i�2T��<�U���q�ލ>�$�Z��@4�N�/,�y�3:�eO����!���t�l�c4B�����T�H9K�ǔ�V4`E�1�b_ѱHd͗����t��Ln[�1�rEUK�ŉ���\I����Zb�Df�J��֜�(n����8�z늃4ڜh��	��j��������'�@�|V�t>�􅢔�#�QJ��S�;
�p��=��$�W.\�@���Y�\ͺ�X���s�[�
���)S��څ7Pw��鑌=��I���a�'m�wxV,��� ��|v��fk=�1Z-�O��Yb�xi������!�EU4BW���.�:�l����[�����m�V9Uxg�F�y�cSq/��V�%U��1��Ծ��z=�n9������vES��`'�*�-xM}ٟ�j��7{�nL�D/_��'�0��
�r����$h�l@G�zР�!�e7�3�����r�Ng����Vp���b�ʕ�5���r�$t�<�8Ł�?������!���J􆕛�OTe&P*��AaviV�r�.���X�jE�9�;��7c��A���TI`q?<<i��aN2�&���jt�����w���f�2�O���1x�R4A�2w��?����s� h��cip�g�sD��±�:���1��:�<����!���U�C����gl�x�hv ���D�C����T!�~��⺻b������{~+�q#�.y��M�"�����<u�����z�q���J���;|��h��,��Թ �>4�J�U��g���)m���ލ7.9�p�i��=U$ �r���$�Q���V�f�!�.�����#k����.ms����yʁ`�Ͽ����#�[8�ҍ��_���?!�E���_�����5&1��@G˘3p+�@��h��,�Ö�����y����z1��6Z�\%&�]#X���C��8*8�Q��7'���I���)�`y��r����w�=y_t������ �5�v�Hc���
�8��Z�^}&ħ���m��AA)��n�ڠqѻ��Y�����M�D�}���V���l����dFڄ����������,Bo�!1���Tb����p����'�jB���燎�J��9��΅oH�=4���t�U�+ ���u�-��,�M��U��pI�<��G���B�Нz+�b�1G;[JDRZ�g���R���ڊ�K=Dg�0ZW�Yc�.��ި�Od�ܭ�s�|my�=��ʈȰF�| ���6p8��l?�mgr�У�Mq#[���FM�{/a�%Z1dFl����*���(�M�7��㴌��D�����K-�*MO��?»"�>[��FZ��z��{���.{,�w7X)n%iX0��(k�zd���$�Jv���p�EGhAG�r�H��eO��������8��๢����ӈu�v��D=s���9����%B�Ss�&��a����bey�����w,<t{�.�-�k�{��jķ��a!_c��#�1kS<^~tq�(�U�K�wDaؙ#N-�" ':N��~�g��dr)�rA#QQ'C�����ۼy�-sz�`N��y�N�ꂘ��q���%�i��I�V�k�\ZS���~�v�B����\Y u�	骙���=���~���J��r����c��Ww���/?�@H�wM/�F���_0U�F�����<Z��9��]3e0h�;*5�[P4���>������?)0�J�WVU�B��"\��" \����@�³�$J	?(�_��@f7�Z�n�6)6Ve3mf�J2����l~��nFY�����Bɋded���~��}�wK�>M9�zߙS���]�~	| �8���?���<Ɗ�Ώ�ɞ�	i��*�^�)�&2��Dd
��r9�v��f�%OM%pKT\� �ͺ9��3Bg�Pyv��Ty��[��ZЊmtOـ��*T$j�� h"7W�:�1�Z���;��*�)�{>����&0L��r�R��y���0T�Xh���j�<'�C�{'��n�"�Z(_`G�o��g1x��wV7�|
+_��S@l�?�t���<��cG�R�y���>��?<a�_�,#(-L��Г�.�d���L�#��C{c��Aq�FK\�����=O� �~�xI�/��J�����k6l��j)�U0�*Q��7�!�)�����!l�*ϩ���8�S�T�͵�|W���˲�X��a��1�@��,e9�Ԅ�����ҒuX�����>�HF~��i4!�	i��+ ��hC��o�a�	(�w�� 	U���ZaH5b��h�v�y�}Y�:S���Ҍ8B���])O,EHs�3m���Fe�� �X��ޮZ@5_"�%3ңw�z�8���
L��]z:�&�7c�$�4�-����+�lm�6�Hb`*K��m�?_e3O�)�+��[��	H�Lʦƥ1l��Aa�jWID�)�i!6�m���� �鉊aY#w��䙤��'I��Hˠ5������%�Jh�:�l��@p�3_�3����Y"У���ca $͎;�-�J0ڕ3"Rs�E�p���ta;�f�d�3h�/��9Yԁ�E���}?>s�5��c2wp.<�Wy�2`�f��tÅ�eH���Ɛ��T����e�[�����d#+��FꇁOR�IA�U�Ap��&.��� �o���`#�QO	�9�H�5�!��aX�}B�^ټzP����`�@-���D��/ɕ�*�r���)i�S�\_��
h��1Xvu��y�8�|n�&����0S;�B�]�K�:q�K-��vs(ܰ�3^QY�z���%@imk<�/�~�28@���Rz��Fy����lx*��D�oo�^KY�y��5�x.^@�( >�E���25;�\���]r�1��M�^��="�X�ʅh�f	[I���{�q�0},h�j�?���(� ��Ԯ�0{��/��\j�F�-�=���q�hN�nƀ$�QJ>+"_�@��:
%]5M��T�mm�8�̱m~�Ԥo�c��m����'��5���ږ�
��0�Z�ڃ�,����S=�tԧ4��ڭz*j:� ��\A�E���E�I`��F�o��A��ڶ2��]�%\����a�a
(��c��ֈ�x+b�:��}��6�J�����j�����;�b`5�u7�z��P�{U���������6}��Nfc2q?)С_�Ƃc�j#}:,#6�͚zZp�;�����Bf� �%=�C�߲ϛ~�
A�(�C�z\K|�u����H���U�=��Ƣ��y�oc��#������m�+�7���z;b�৽���dTX #����'.i�_���惵�_ѱu�>j	��᥻?]��cP6Æ�鏣,���K=!��e���'�Ԡ�ET���c�"�����K��]�m��t��#J��x�ľe���]��6B.�i�>i%:��X݈1��.��P]���S\�7��U���^G����1��-xW;��
��F�N�6�:=���u�#G�/Y����s�dv��4ŀ
J��2E4~~"!ep8}4ֹV��D<R�Ԙ�ی�!^i\���6\T�PJ�'ḟ�_�������f�)
���6�mG�-� ����A�|$4�ܨK�$�^��0��UO�Ԇ?`3&�\����HmV��5vT��T�~F�>������V��S��G��5RA^G��Τ���2�#��U$��r�z�m�S$�\�7 �Z��"����֤il��D�»~�e�/�ͷ�7,@�M]���6���m-:�k����O]��n��X�6+���CD:�j�@�	��1�H_:؏�{g�z.����M�-���*�Ӿ�q^��u^��X������߭�������v����-eq1���0�e�'�}�2'H	�]���Ф��քW�eu-��E��,*BPY,c�����`��0^D	{����4�~Ed��������s�U$��Z�� 0�@�<���9��}(-h?嘵�����[�?Y�xܔS��h)��CBM�ш�|�Y\�Ъ�K��˂����k��:�~��X���*G��h�-#Lp��xh� -�͓9��\/�N/Ͼ0<@gWڐ6�,�C�������z���Q��n\��~�F	�K��YJYК��g�7h���C8+](��otN.7uȖ�(�2l?�&�Ih�G}9�!�y����%����s�Y�s�/g�%w�wC��y0��3����O�RH��Z=�e�hH�����:������+��kq%�)���p�.�nCw�/a�'�eت��T��<�.\��"\�_��0#�)'���q��p�F�kI0���}k�����:+���|�,�xE4��CH���]Nl���b����|B�N��C}q�ӟc@\�مQ省>�д���͟3M�{lv�!Y'@���v�f�3u�]��h�l��YϢeZ6��E@7�i2���./��4��~o7�i���J���f��[QjЫ�4�#�&�9�X�Ի�o:��I�5t#e��׉;�F���/�e�EPP��Ҿ2����Qf���-��H$D�F�`���ƪߵ�X���[�g��i�&>09|	,-Lg���>͔�'��Mʯ�X>:w�	"��g����
w3�����~�R�B7����8�A���@X��/�ժu ���H��)���Vhe�Q�λx�mkU������u�V�4����$�?Or����sJ��@������%s����5�6v�7�'Qe�}�	&�_٤7U�+2���˥G�<��jb������q(���Z�($���i�#xS�����.��������㿫�T.k〣�'��MS�����i�	�0�L֖�(K�ۮ7��2w�>Qn���N�d�����ez�3���1�����8Ί�w�yvp�9�(��g_@�4���)e����ޖ?}���Hz��e�q�b	�Q&�0��"P��#�.�c�� +%zh��ΈWQ6��T��$���;'9E���D�a�Fd�1?,dx4�L���/�B=�m��`�\���!"4D�+f�\+W���
�����j����|9��]H��'��f�tDRN�/�B ҹQ�4hJG�D���O������j�����fr:���)�)���$`d���+Qs�Q��"C�הl��!�z�� 8�re��w틲L�U���;�ԲD��J�&`���<�5nNN��$��z�؈c��w��h��mfL@F߱@S���L��+��"Ճ��}ʏ�~dO`,��k�'�
5Դ��țcғ�F^��Py�Ё�� H���\�[�����%�����o�!���#�4��.��@�{�
�ݹ[�ȦH�s�/��,�j.�������a~ٌ��KA��B�	k�~&>�ֵ�̢q�������]P]�&�x�k��'�#���o�BHe��}���)��H��>��*��lR�?���t�k2�K�!k�����4f�<Vq[H��Lck'�,�n�cB�&��g��`�e��ָ!+�K�@q0j?���Q�:?�6*?����慤�0�#�
{����1�ʂ6{m��� |2yh�	�����7|���kT�@n��`p�l7%Ɋ�bz{�k?b��ﳿ�d���2g9(H��!~L������G0�K��m��2�5�Y���,���֞��41��H��hmդLKY?���T�X@V�K�fJ���)���Ƹo�Z�!�EQ����-���l���tsB�\�<<�AX�Wi��b�w��(���6�g�?R���h�8�6�ج��p�1���C�;�/���\|VN��?�|�ѿ�G�È�.�@wb�#�Z�+/ܡ#
�H�_'�*�9��@�E��z�K�S���j!�����]�*.3F�?0�m�*��/��>̾�;�5�YRfkB��f��=���;xŽaW��k�$ySQ�������cT�%�M�\i>�r
�9��f36h�	v���`W��{/�Ů��?������v*�x�/y����g,yXS�%B1%;[���l��5�{��ݖJ7go�oV�e�W�&*�ܑ~�3�����U��󒵅w*�-=�L�ލp�(2����X���tp��	{��S�ٺ�����u^y�-,g�ĕ����=�� ��9z�����r�9}�G�K9�hyd���}�	�d�j�G����y�f����*{�J��=���GY�vL4B�ݪ��.b:�H��7t��(�}k�B�K��T��v�xճ�J�!��9��RA�H��y]�mA`�|�s��.7�#�~/�&��(໖��Ѹ̐Rd�z�$*���
ܱf]ڤ��J�:�+�#Uo8%p�K�ɶx�#�m�z���&�q����E�V��`J��Z�Em���S��(�2�V(o0�_��#K�W���j�Qv@���",9�G#P'1!PVV(P�RKM�:��� �
*���yKv�R���=Y��}#��b�
iUq������
;H���'�lF���lR��)�qzas#Ը�����#r��.�8F�֖���j���,ɉ���C�cӳZ�k��T�V/���V�:���5��%o�������^Ut����.�
f��t���3���Ve��Mȹ� ��!`�Ipti���C1J7Ut"NLe#Y���V��4n��d�1�y9�V�����b?Tj֝�]�zb���E������@���襐Oh�yO�Ś�.b��0Z}�E����&S����re���u�� �gx�	��Xtb�n&"�?y��b}X�݅�w!m	��rֆ�Z��m�P�a�Ĩ�\9��'��.���J.����4C۽*ց�.�3��OwvD�a#q�ƻ�1°����H�?|�b�G�~yC�D�Ɉ�gW�2��\��T�9Ł��F����T�W�oY�?,��Ed%U#�M؆p�{��.=]���QIS����^����Z!C�Ȭ���@h����"�=3�����ń�qL�ȱf�b���k�,���{�
U���mu��,l��3�g��	�["� ����E�AM~��ژYt�1P0��ʮ9S���ѯ��4VmC��sN>y�bֳb�Z,Ω`��kA�۔����OB˶Sێ�1� �Փ����s����NBި&��~�q�r��݌xZo�MjW+�m���S$b2o��g����_X�+Z?�l:_H/����Ǎ��W
T��5��tܿ�6%�b@#���
K*m_��,;�		��e�	�+wRc@/+<B;��T���\�F/\'M̶��S�=�A�wD�6���s>l��	>��ACѵ������3�(2����S�`���??�2w3��XV	�sK5]XHw�C�Z���<]1�P�y-�oKمK� 2/���O��z_�s����|H�7fo;���&����*��X�j��V��#"U�:H�K<�	�&����Y{#F�����-��������D��cO0�:d����#�d����G��D��6rd�F4�ڄ�a����vi��>VC��<�
�FUmj��~.L_WvH���@S�� ����(�՝;���>�kdO����6�a�"��Oꘊ;z)��y4��(r�i�3l��!]�;�|F���a��v!�!�����|�> �6�n��'����rY���/rΪ8��8����&K<�e���>���X�~��x����`��<�nb-�9���d�-�� ��Z	܋t�M��0rܐp�����c���*�\�8հO�Xɳ$b6��r9���w9���D4fr�U	p�rRF�8�W����'x�N/ ������HhsaQ�����M��{���䴎��O�&���]���{�T�+�kh�@6�f��p5˂ҵjާ-@"��_{���MCr�^ù�O��텚��=uM�CO$�F	w�c3�ij�aB����k����.�@��^*���̞2�DuA��U-7�����caX��vb@ޛ���d�?lp`Z��=��X��n6�e�)�3���$��saTq�Nڢ�79�B���"���2��Ie䵲�38��I	cUg�ǧ#bk=��x�����/_/���b���&��s��+�teAz�92?��)���W�< 2��N���O��9$-��s�N� �O�ET��R_�1��V�[����Z���o��I̘<D�A��P�l�)��t?���!}���jӺ��Ⱥ�ca��E��
g�4�_�)M��J}W�s�����f���_���� ���b�����
~̜o��f��r�^�eZ���U<�6څuKGq���*�hv$�L8�=��L%���)����OEfiOdN�"7M�\�Yw��l�M^���wjK�m����-c��EN�'~�巖�򲻁�x=��5n��.�C�1�d�y��M�^��/[ҷWr����|o���:"�fҿ�}�y$ę H���\^�}�+���/�I�Z��(�L,@��� x��{-���*!¤� ��|�
���Л�������-\).��/�Z��'�x�Un�c%ej�C�lx���ݻ�ˣ�I��ȗ:g��,�M|�EW��&�*/����o��Y��?c��}�YX����+�#Zz+58���2�>�Κ�R�b)L��{���&����c��ZZ���>*��zq
j��/Q�0} ^��3�,8`�#��SI�]L��236)8�2����L~��0�ȕ�IF�u�1j:��u`S��.�u����s�aƩG�e��am���uo�+w����S�t��	̻�2�^+;������-/Z|R��XX6����T��H�B��L�h��Ұ!�,��1HR��r��O��;� jRV�D��d�����3�W���t7�0�x�=�w��-�^rWk�q}p��]����C���W�#�ñ����8�2+c����j��%SL���A�u(��ܓI,sM�x_�;~��t���W�CB�N����6f�/�M�����tH����e@\/���ka2�\(�(�w�~��CB���-��<tp���vō@�J��8�.�L��;�_��|g���9\��C�F��p��ŕG�'7T�`4���N���\�^|�U�cJ��B�)�I��bӊ��LNwew��Y���S�%Y2����Mb"������2��>?��^5�q��������]d�,�&Q��~�5�YC��߄\'3\��ӭ���ywI���������2)t�S7Ό��5.���I0��T]� w�r�i@�â1�k��� [z���v�[�)�&��&�Aid�wG���u��̄�wQi0R�;�Y!�-����â���Lh��.�`OC#Xq�s�?v�`�+�-�F�cA�/f����t_��)C��0�@D��&����g���ٽO��W)7�>��PR�W�ŧ�8�M^�z�pu;j�EqV������sW)���k#n�[S�yn�%�^U�:1k���Xw��E�A8�Z6K�_@�S{u�2��*�QJ���ZKuKD;�4��`F-&P;�����S�%7B���\]�i�sT�K�?�?�e����Z���W�K��6�����m�"\�=���恪�N.,�Ų�Ǚ�C��*����-V��	#j��L%���5��%j�:��;E�eB	f ��8� �����vs�Ta+�QϢ�O��Q�pH������i]U�d��0
��S�"݇z�%C���v���"� �Ek"/����G�S�������mԡ��D�V0����ۢ����}�9E{��8�ZuS(��8�y@;]e�W}�t�\S;��\ t�W�%������}McT��G* 5�&˗�oمo����k��h����9�	�Ea8R��±�z�(��?=vR�^֠1���~��H����@���B�TE�N��R�Ǥa�*p���iK�S:���.3պ����]�UiY�O�a��?_�F�T�6�2N �MS��K^�C��g�(�TK"��l^��'1(�����d4�K�g��o��H9���y0�n�����y62en@�y�����$�В㸎��~t	��Ҽ��Gd+���s�`-�SZ�������`��l���̢�cT��_��3����SP�$�}�O��<h0�K����"iE-/��{:�ᒭ��/G�����n�]���(}�9��q d'�����p�̇	;(Pw����8_�����ʑQ����JI�[�k!sbw������CH�?h�UQ���P
)�(��\
eʫ��!�'�����3�U�8DV���dÜī#���ib7w�W�д�͉��}�1��v�oRj�b�3 H7����o>_@�O��Ai6^n�����7���
��=܎�Ժ�;�z��{I�ۄn��t���F�{?�������E̠��!��uZ
f(�a�2=[@�YA���7̻����Y{�͔���/��<��	6'w�W�[���u\���Z����`
���-�N��,�D5��U益��ek?����ۼ�,��n V��#�;s���p��N�Y%s,���٢�no�_� 6{�����eO?rz�?����f��d��P�(Sk���Z�����9���Gk�>��O�=҄:!�ψRx(=�i�0~��Ib�f���<Mu�$�&�Q�V0��kQ{f�z��J��&*�YKu��p�yw�o�]��	+����.R� ��@�w��[����ͩr��tJ'��54��x���u��H����_l�wHgaG�Gܠ"���κ攄�ȣ�)�К�)Q150� S�w�btGh�>3:�xo��Q�=�uM���c���(�T)��f8S��߷��֬��?�$е��z�oT��ě�Ҽ�'(�/T9�4�~�[/���k���Yl���A.2�+�G�$�t��]B6$�%U7_�(yM�H<�P?��@!�ïc��.#��/ƪ��!�k���9�1�1r�&�N��Q&��.�HTa�ce��*N�]�W����h�)�Ŏz~�i���F���/����5̹�g	�jw��a�!�|�'t#�R��)��i o�Q+�Jw�����0��ޔ�ƥ�zN]]2ΐyP��Y{�� �0|K<�zա�����A��,g*>��H*`u�8o.X�Ӆ.������>���wϺ���`(�B��2Vv9��ڕ!Vr�uG��T�Q�+� ���wK�_�g_���)��uTP�Dp-�p��3�\I9���(�(�_�|=_��UpJ�ܴy64f�Y]SU��������p�e�����r��Bs8���I�0�Y����5�N�ն��WI�+�$�m��4��d��	T�g}�d1��8�oa��h�E��.z���H���g�m����H�祥J ��0�ZS���X(�X�8C�Y�P���+����_ٹSmo>���[���m�nn�?a�ȋ�x�V�w���n��|��Ne$ʀ����1JR��F�U&&�j���r*��~�b��Z�^��|,D�����ˉH�M���|�Z����7]�Ǧ���'�@�����֜��-�a5���@7߂�h^��s6P�m�e�JE�K%iӋ����p&`�,S��H�
�ehP�7����r�
�E��b3w�q�����LV��#�{��fW��I(��I�*�Rriߖ�)�Z.�u4��/��p�o>��Se+�0t���1��>��9.��6Ni`�}��{Pn�]%�f�e�)�0�t���ڙ��d5\�NC��E�O����?3p��r��2�����=�꽤\c�3��r4�6��,�5�Q}oD)��M�J��;=�"kNg),I�#��^��z����a*P��\�5�O7��tWk�K�&E`mjy^�ɞ��o���æg��x�;{;�I�mЁ��DʓDz�'>-Z�T��QH� �R���
%��M�Q=$��O����_:��o̀�Tҥ���� V���hpb\qF���v�`[���a������!�_�}�ר��?�K�Ա �5�;��wu17��� ��3� ����)��+������+�+<��g�/�Q� �6�)�u��y�۠� ��� 7�ƯP�=�����dS��S����_tc6�"	~8�gG�+�e�xMY��o��ł�&M��s%��o4��ܢ�ƚo(
8�u8�%��i��*�Za��G7Ru���UZKr��w�j��0���[���s� =����� �{��-��I
�iI��z4^�5����7�Q������R@�1p��[C��!W<梭�h�	Z&<`��{��%����[��ۜr�@�͌����R�Q
����Q/wo#<A1��csY	��+�ԑ��Ã���%�;j���Y�	�b��F�������O&j��A�b�@�0!PO���;���V�{X�	<5�_8��?ݚh�p�"�A{�E������	�W���!�!ꕰ�Q{�8OcR�t�<==�UP}S�$i^��ݴ���V �rw� �&�V��e6�����ʜ�*�˰>�Y�ۑ�?)��I��/K��S���8)r5���6s��;E���l���߯]a]Ze4�{h�G���g�C��Ib~����#fA2��\nr���H1�f6\*���q��j)�����R�-(q��@�lCn��(�tn�gj�;�y��rE�#��E�)�m����}�)�8n�&o����}����ፇ�������WN�����)I3".��&��r�Q��f̑��n9;=U�8v*f�\����T��;�s� UZ>N�X�����'1�xo�.Tˊl����Ⱦ�)P��` e�E�:i�_8R�F%ˎ�^�YLم*�{����5ͼ�Ա��t�B_���X��]q��]���S��d9r|�l�>w�|9mqL/z������?t��#�,�C�C�&��kdr��`�Xܸ���a�6�>���1p�b6C��|'���ްi�J��R����5�j����ȸ,������Ը��E&�e�]��"�H��XM5]�R�D�a��ʛ���n�^�m\��OA�k�;����jFo�ZÍu��'�Ĩ�͚c���]C	uX��5 ��"�A3J�w^����>}�CLlw��ec����vA7ٮz+����������͑��qAZ|��@P)H3��K�6�]����J(6e����S��VƸ�; y�����R(���R�%B<��� ����@W�D ǎ{����)S��%�2�*A(�����7�B��	�X/q#�f�N�4�4�s�3�Jk�p9���e�Q���:topx�_N���^i���l0�wwWF;>9��JoD;�P�eT���5����;A	��<`��o�œ��`c�%_Ka`i�o���v��PI�Ǳb���s���`��/������]�˶گdq���b�)HY*"S%�EE����s�4���H����(�ٻ��S���![	*^9�i�μ��>�
������F�b/*:S5�Nm8sbBz�s������'������G���Y���*șZ6��g����ޤ��ï,�d��� O<pAU���e��L�yɮ}#�ē���ͷy7�����<N�h\N����E2&����i���G}a��ܶ���C�U9n����C���qψ$���(�f5�Xn�i��f�O�EWF���cZ�LZ,v>5����7�z�z�((©O�f�P�!/t'�&Vf�{o㷍��!��8#V]�Ǡ]Ek_N����7`6�V��;gn�x��@����+SVoct6�Wx�c�jIH�b��I�R�0Y��R���p	���`'C�N*��q.��*�A�{�l.c�Wc����֥�x�ڕe�\����C�֠�&��Z�E�U��b�߇7���M�e���l�����$/Ft�u�њ�~���*��Ig�#~H�K�^C�	�8ȟ]3{�Y���I!����W�lj+=<��t��,:���t���&�t�U6���M�2_��Z�Ā�	��Zkm$���*�8w�@��vc H �n�����r�wIU* a���S�\$P3A+=�.��U4�"�ŀ�a���w�\���Ks�JjY��bI�s�v�'m^�.�u�������.�:r��D��8G$v��y��G��{u�ѝ��֌;>7#S+�5VY 6.�&�9�����sE�ϛ�g�ȯQ3k؄0�h=������Yn�SFD����O�V���>��o��z&0��L3�4���2�gf,Z�7omU��<κ�mʬkl_a�����<YV��'gS���w�`��08�~Iبb�V¬8�u(,�g���y����������GՈ��B3޴��G��Φ��]�.����e�l����2�i���fd�R�%~�ܓ+C��i��/T�.ET�AC�u�Cl��wo�Q!��t{��Щ�^�� �>`4&R�|�ş�p���=�������ҷ!ϲ0��q-���YH+���/���%E�[�w�����st/�2��=X���P���~Q�d|���@6��(����e�����f�2q�N4p�־�]�7�ՙ�ګ��= H+V��M<a����&�0-� ���J���Y+n��%�EH���w�M�pan)��u��VFNu�/�_��/i���!���[����h�~�RVn��G�G���j:�:O^eu��Y�D����������c����t�+�Tk3);�8~V����1�C�Ʀؔ��W�IҔ� ��_�����P�'�Gi�����^"MR��"�\�wl�'H�1^J�?T(ĕ��2���u�o;����mE
~�޽�,y��S*�v
����[q!}�����%�����i�n����\�w����^��LU9
��'�&�2V�a�������l�A�eI�O�4@��	����v�ӵq��iUS��+'ɹ4)Q2t�6A�ؑԲOIjѱ�+S}�5
��v�?���G!O��j.!;�����qg ty4xB%�7�!��U~�2C�����3*�?�\���Gt!Bͥ/�G�)���0�m+؝�]�D���C�ͩ�#�y���E��S��
$Uaj�4��IK�0��Z�"�!���[��q����O?�1O$ %R>�*�S�3]A��%�Nɂ�R0��7V��ʥ���}�~$,�`�M,N�Ui�����'��Py����Z�wzO2�ݺ��I��T�jz�������V���ŒP�q��U��60$�Lb#�ҟGR^�� 2t���[A�oE(�gR-�V.�H��������`n��֊!R��ZP����y�/;u�ʥ�fBZC=�_��!�f��"�x���U���z�ٞ�u�ǌ���{�CJ��C)���8��1E�v�:y���P��]����\;k���\��\F���N�4a��u4uw[����:.�GǾ��<�>�v4,���/�!��@y�G^���o�z�.�Ӹ�]��}����ýO�e�@�g ���� �T��<�H�ĺ�)�w]��U��K�X��T���a�|����#r6K�	��v�/Tc�{���jTZ>U�������U���^���l�?�7/����Y����+��3���al���KΤ��x��@X�Nʣ�����<�{�n}�1!�>Ѕ��9Zl�P���e�jN�"5	���؀B~�Cwm�����T0l$�x�Lsu��ݑ׵������8�v(`�L��a�͜����;��//�FȢ9�#�jM�ҁA��Q*���7aM�[��_���I���{�͈$s��0�ٞ�b�#$Q���[57��u*���c��d���Y)��3�f�wQ����f�<�.�\=
�vhT�g0�RSr�X)�(5���՞��B��p�c5N�宂J���{��8B�Ζ�׳R<�;��o�+\�z4%7˥6��/UvByz�W�����x]�Q�f���Msɑ���3�4Ǜh�9z�i�ut�H1�|`�Q�%8A�ؾDs�FH�7���H���!��ט����\�$:9}�8|�vE>�[ 7Ҡ)$���7���>���o�W�,kNP&��j��%��i�ap��^�W�dC�j	~>`�^z-�W�@��Q��&���g�ƘKcz�'�|xh�H��S��ْ�F��u~�C��g���G�e���1WBk�+=.X�#q_X����,+v���M^R���$������b9^��p�[]�V��To��.m ô�{7���?��\�Vt�-t�����A�4ӤmHS@�{���S,���۵����P�ttV�L�$:�0�q}S�V)4ן6���.�ẖL�M{��$��F|��X��躠�*7��U�J���>1�\*t�6m'�0_�.ISn���:zS�Me˻X�0��)��2,��p�s�]	њ�e`�㽥ǡ�l;� "�l_��WO�H�h��&�^��3 �F'ܭ���T\��a�*��W3�t�
��c?]��s�MyT2`z������bvFzX����,�L|7�d��L�x	u�+�G�t��
��Fs�&RP�I�c�r���Q0��[��b��(�u.8��*�S�e��j�A��*�]$��p�耉�E�7b��G�R����3k<���K@��S҉+&�I;T�9��#��5a~Ҽ�����	I[�d!`'@�`� ?��T+A�2���P6U�]�Q�-AٶS�v�f�,A�f0�����p(��3x�1�E37r.1�jp�������%;�OS~�j����"�����sf�w9�%�Պ�u0
�T����f�~Ă!8>VkO��[O ��>��z�`{ �R�:Ĥ��8����8�oa:���/E��N���#	z��]B�7a<'\`�B�8����O/���^�0��U��ޚ:Uu���T���~�@���3��Ǥa0зV24���v8��e+���Q<�L�:F��Y!(��}=���C�K0���q�
��ޱZ!�.�%&���q�EYvC\�؎˳r���1l��mGS��0�Qn��K�J�«���?�&�[��l�d�)�|܏���ͽx����b .|}�3�DQ���t��NS�<�!j�9w��G�	��_���`�,��5�ܪB�>i�9aNj�׍��ν9+��B�����:����1}��l�po��vQ4<y�פ�x�Ps��j�p��
*ڐg���r{Y�e���wX���������L\�,��p���8���9vi��3v�� �~�/մ��׷ԗ��Z�*r��ʷ�d>\8�J�q�jc�zM��DoD��x��jK�H73T_����h�Q3&���J�.;��Ǉ8�'-�y��8�<���������B�p�k��sh��m�������8(K_M5��hϥ�"J�H�'�~�����[6�'�V��VC�v��Q����?"�.Em�,s�a�4�g��n$j����4~uB���&[vܥ��y���)�2�:m?wadD��[q� �1��_��I���@H�Z��O���*�/���<��<N���q/���iyO�����;�0�l+>��죑��C�؍���i4 *1٦���Ɖ� ��w���8\�0�8���`��^"���Ԇa�y{h�I�6Rk��y�i_�mњn��:���ղu�4��d��_�%��kY[���E�8�;Lh��T)����X�)��-��.}h;8LS;�.�[ȯ�����"6|�NL�m�}4D&�c�_~TT��Cw��	�尕�unA�6H��b�%�a�ZX�����'&���G���ǳ��I�E��`�zT�rB��I2g/t a��'�꥚)�U��!����e����g
$%��ڽ��l<��2��� �=)P�7{ž=��Q��x6MO1�N~Ҍ��Lŷy�tsy-��UQ#��R_ei�@�D�g�e�*K {���jR�'Vezv��q>�x:��ƣ�
J/� �U��WL�~�ْ �� 	ӿ�������Ҵs����ph���#/6�&W=<��	j���k�[��Lr#
wF�������m��dj,���&��o���g)�w�P��=$`�)f�^D?�.][�d���o���]=��1�
����-J)�$��j:�\՚��_�Ra��t�����U�#8����\_ ���%�g-�F�,u:?�D{�������~V3���`/5'�k���}��Y�GA�D�m��5@%ߙy�!���˄݇FfD�ۄ��}\�����b��t�Ol�J�N&s���:k-!�$� Ge�	���=1K��V��oJ��9����|�z�i!��(��%[��h�t�_�X^�
n����dPui����i�!�m��n�1��o�5�.%�B�GN��p�H��%�P*ؤ��q�f�ګm�X�MښUE"A;��������q��r5;F�OP���<�+��=��\�])^��A<Czt)�Lm���8��A�^��8�Dz1���X3��
+M�I}|w��C�DL��4�ғ���f7ùdC*[��e1�l���֟8���5`��A�_���t<!zé�W�VA��6��kt��xC�̡�V�w�&S�m����9쨜 ��GU��F�㒡Nű��רV�R�'�D>����2tQ���to���^��=��0d�pA�}�}��0�;�'�:����3�yP0��2�/�B��3��a�,5rIq�D����'��\j�(�^����FI��ȴUD��K�!T�o�r����Sd�+4䁕6�U�wh1�r�J� 	�-iC�i*�T�3��N�"�������d06Wc�~�^����c#����?Xb�X�O�I�I��)ɄK�P
z������g@U1�'�L{��]vƉ*�j�Ѹo<�k�ޑ�ЊEab%����I�2�_ẁ�J�O�_|v1,ޗ�IJ;o`�O=|D�h�*�����3ٳ����.�d�s���@b�a[�q�N�xK9Z�	5��O�?��D��s&v����F������&����g����:ta[&Z�&hr,qz�����luk��T���g~\�<(��GҖNL|'9��٪>|��;�z��	7��ٷ�!d�b<I�m�7�i���5:Z
��评��0>��Q�,@�{Z���R(V��N c� �o�b�� ��	s#X�KS�=h���m�(���=O��R����^@ů���p�����7��iz/(^���G��!tC�<��]|;5�~���9�9��Q���I8p�\fh��
Z�u�^|]_�&�F����͖&(���ЩB$,C�cT?��蛼9�i�W�q6���ʋ+yk!��l��a�sP�������Lf��4�Cƕ&����-ge��[��gv#���mZR���oD2�Q�h������"��]�=l�P��Vc8.(�F�*�D�����o<��sP�ϓ{d�ݞ���@>����b��56p>0;
ʖ�b�>7��Hz�ij0���
�SC4���>���$�9Ƭ_����|�j'=+��3�����/��%`ytޓ2�cHv��VAY ��c"m�6�y��hZ���k��+��	�]�/~�ȓTı���X����'U�0��MO�~�Wb�X�XQ��(p����TͪB<j�jE9��FPylx�͌弉G���_ޅzm`������UT�!�U���/C�>-��}��lb�%!�_~u9�\�)5��5�Iɯnѡ?vO/h5���H�#H�.8�j�u��3r��ކ�_��L~|`D�`�	O,#��� �Br��(�fD��_��O6A�A�:���?�\v橙s���L�$��66�y��.�F�~�Ά�T�QA�̷��[l��(��4��/��6�w��=�ͪ#|�Y��j�7Zkd��g���H��H:u����i�x��#����Հ�b�_�@@S�c���Ǻ�Ȯ����-�\k����ɗ�=鳷��]�:
��g�(�Ǡ����7�Ƒ��֮����Ҏ�VD��Ł�M��?��Ŧ���ίg�_�Af�ZO��J0��۴!^�PjuB�����G���@�a�f{����+���#��%_z;m>�%���$�V�˽U9�����`b���� �f���dfi��}S=\�8-����;d�9!#ݽ�ea��� �g=��u�KoS.����b�ٺZ�Ȏ+���-ظ-
��Ձ��_NF�w�A��]~�=�xpK�No�p9���;~����XQpn�V�T���*zON�z���(�\�ւ�s���3)���E��Ћ ��I9/O�p�n�DѝW���Q��NV�����X����ss�x��}7�s98��T[e�Ǘ(w�o��1�·���7 ko�T��-�z�U����CiY�X���� E�ɺk��ӊ�iݛ�w�Ű/-�H�D�{ʶ���Ox�#io[{q�@L5)��{Z�'���eiLJ�U�W�!��cB��;0��.�[��.6&�V��g�Um��v>x�N�"	��9|35�LSx����4~�*��=H�@��
[,���44b�<��O�Caem2��� �IvHnpڧkm�}7�@�f��B������Ji��$���C�E(��%.��=�x��X%l��;�J6�j��/s��V�r1��h<��n_wFq�0���Cb�uݣE�7�ē?�����\c`WK,z������vs����Ǐ9�=|k ������D޺b]C���m-�'P���N���\�V�~4�ժ�K�Zފn'IU�)]S^���W�P�VQ�laޠ�窖aoQ9��'��F���7�ZQ������"#g��R5eKvo�0�>�߸4X�v��d²Z�&*�UyE`���&3���̑x���ln��Ƨ�G��gS@�Z0�AI��t��o�f�ͽc�<%g�v\����%�&6��� c<�5}^��u}�1��7��B�v~�UY��]�I���Ƴ��D�kJ�[����@����kN�Ld�.0"�Q�6NT�4-Ɗ����?�V·�u�|T��jE��o�v1+c��;� +T������{��ɧ�z m*>�U���!��G!A��4~W��5�,4惡⚸B"�)��Р���P�6zO��y�p���Q�u�Ix	����MH}:r,����t�8�4�+��{���ν��|Ym�¹r4�Bdp�b�${�ڰ��G���g/��0�b]�D�P8k��f lnb&���8E�⎔��cD��b�U�۹���}u�f*q�+K�QB�K)��t�z��f@�`߁tG��1h4eCڜ��Sf�w����m5r����R�P?k�*��5C.t=�T��x�}��0~��$�9!8E�`@X�w��@�G����x����F[��?��[B�O�/;�1�h$��Z�W��g����S��p�C�S�¥'>�%�V,7�G^�$��y��>j�G�im#Y�p��*�tYU*�o)lP1�n�q������U�#� ��'��Y�aqZ���t�Q�-��&UP�ɕd* ����*7Ϛ�жP���F82�w�1�a�=�zє�f#��;r�˙`Q�jv�6í���O��oĵaf;;���1&b�GYKel3
�L0d �׼��7n*<܃s�X�y�����P��x>��҈��z��oO���N����0j�{Pl@��=��q�jr�Qb78&��s��gB��'�R�5#�U�Ƴ�i䯰=cd|�3��q�7��e@Ѐ����}����lB1���c)o��@�M�n��5�K68}��;��#MN�T�����?���i"�\�Sw�����3z�nhG�!~
Q�Nle_]��(S��JI��?�3_6�+\5�F��<�%�X;9�[時0�Z�B#�č�q��
 �d��=C�	�]�PMpX���cn�M�}��[!7�?\�G����:��Rß���My��+0��;Va��6r$����A#bܬ��	8�zP
�8�8�Z�Ay��;1�g�#9o_nH����d�����W��k�����=������XR�|�9��Yv������A�Z������"�9�l�٢f�2���Gw�1AS闵6/���e6�z5���9�T�A#�����E�9�E��oFb����)�B�4 ��Wq�!E��]��3��G��v�3�_��z7ʆ�f�U�@E�H�Yk��f�S��h�v.&�LvQ�fʼ����*J{5��"�Ip��4ణeţT޻�����κ�2���F˭��W��w �z$y@�<��,���_P:�֣+ˍ��B�	؛q�?h���d�2�����{3B&���݌�]}��;�$��S1���e�;���X������1u[����oCc��Y�b>��2�[[s��@@��P`\�]L�R�'M�l	j��W����Fb��#"}���zC�[�M��5��\v���������-�J֔�X6GkFa�,�2��&�dp�hrh�grɿǿ���f���I��IB�u�*�ܜ
���ύ��"��L�X�R�*��z��N��1lx�����
�p�����V6ǥ-�,rn��m�3<P��'�k�[W7<��F��u2�:̵x����l�)�(L�����x
�z�c��aqS��0D����sd`6E%q��Я��S���=��@��:�휡�˩S���#�m\����H�K��P@���4�Av�k��B�k_�C1͏�N�<3�5!�V�PG��_6�`L���Q)����3��V`�e�6
�?=7��i��C��½}cu�`�d�f��6L��1^�wL�����@���ѡ�u��K�����Uɺ�(����wB6�* &+:�����Gc�����KT�A<rAĝex&��g�Q�=Ԃ��z/j�ʹa,����-���|.Qq��Orз�+=�F���L��ʦ�Q+�Uk�����g)?(*FH��ئ�M���[dj?_uɅc�����j \8���Q���n\l�ܱ�Ouw�%�N0(l�Y���y�(�Sl��n/�d8�/9�X$m)��U�R3	��؎���1��M�� �я������b:�>����ԪZ1�y���{�"��0�캥�b��(Y���%ҴZl�������7����A8��=�NxK;gao�,�F����4�Y@d��qYl��Xn��(_U�#1�H��#q�P]�H�+�h��>�¡��C67t�&e�5D)'b�{w*@4��"���>XMsL��;��O���h��Lی�t ~� ��7H�K ��X�}Y��Չ*y��ꛒK���oD�������4l#W�&D�=��������l�xr�ǜ@��E	+iᇉ��p(p�Tl[�RZ�dT��~˙���\ڎ��45A2�Vj�
 �690�E>�՗J�-q���_΍���يn� P�R(%���������{#�IZ�B�o�\��@z��8x�|C�|w$�c�(�D,<���o��扐�����u\�ҴS~Yi7/�ǈ#�w�1l���L=���LvѽƑ�T�s��;�'i���L�w��ebhXP�x�i��9�T���S��e�?�;ب����/��9�ř��@2	���"z9YΩ2��:��R�j���)���&�I�-��ӏ���:��s��.��&��SɅ�?���p��\08�3I]`3W���Q�{�S;�b����m����j��j��X1ƿ�y��	ŋ{����k�
JE�J�A�r�Y�9'H����^�r��E]�Ȱ[�����J/k��<����o��w�ۢhU��!U�_@��F0����V�ܵ.�����l��� �&�ޖ�)Q�8}�#=u�6�8"���M�kK �2��^�Ę�>�R�.|m�|��Nؤ����VDY�V�t�~H-�����A*Cŭ�,�o�LN�ynY������Fҝӛ��K��T�iGgXj[pA�h���;#}��i�A�j��qA�ض�����pp���7��Ͼ�������t�N�c`�WL{W4�ܩǏ���9w:��>��>@0W*34`H���E���8T�!���9�Ԭ��&lHj��Ǩ:���<?B��T��4�=W"���=-dכ�DQ��6y�w�w�H�L�{7xT�M��iJA]UB^��铫�>6@��\��
��5)\��E7{���2j����Z���.h$���d{�2���.ȎcI�c��Q!!�l�_F�Ѡi1:� }y[��ɟ�a�p9o�Ż���k'�2�NDlu�X\Q@���T����Sj D�p���bo[Ěyi��ޔ�wF�V��=����4҉-"��nkA��PeF q-J�TixV��W/�^�9��l��
�^*=���h7kT@E�v�l�x	h,:�s*0�#z�}�����H`�,�}Grv �	]bj�Q�U�CLdǥ_,@Ho���O�i�l�C$�D����U��v�`g%<��Cϫ�7[��J��\b�0��s���rr	�7���@O$��jL��C �^?�'��{t|�Ō�V�ځ�V�Ŧ�@X��!�L&��l×{��=Iu-yM�#L\mY�e�?-o�q⠻m��%GS�*�E0Ԥ��5��G�QɜGB1
�Ħ�Z��x��+�I�����@]���W&�JCsQ���S���UD\6����h2��N$���0|����<3�s���G��e���uX�G���C��;༳s���\N�^ra�%2G��{�hl~�5J�{XB��]�.�vI�t�Ƕ�[$d[�¸��M%����d���sC��֕�$΂�P:LH�>�p!8,���oOQ�G-��j��F7Mɼ9DeD_�Y�z�t�EsIH3u�VaX�K���D�O��^�D!�]�OwD�z�3�_�h@�x*�!��=�9���=�Xs�`*"B�[ǥ�'��iR����-AkZ0k�P�S� �ՙ >�S�(�j]��7��؃�]����z/���\��T�����{zO�8�4z��ճU���1zh��
'�4�˺�Y��H�R����Á�����s��L�{3D�&Bz�h�L ʋ�9O�x��bs<ED{�̍G���C��,Q� ~�N��c�Ԏ_S:�+
eM�o�=������~�R�7Aq�e�j��FɔѲ�N�*Q�ʢа�0c���>m��AqO�^�C��oSa93��ؓH,�Z1�0V'*�\�'�j-�$���������~�$z�7�DZ5=v�0����~�D�� �~��m��E�z	�xʌ��3v��Q��c������ � ix 2���@�`�5��4���z���#�$�n�5�DoB�-^���|�I ��!!��u[�ɋ�ہ�z�	��=Ѿ%������ľ4���ހyF�8te���G6h�al
�}6���b��>;,�؇�֚-�A1�������eg�B�K����g�_��/:��.�$Zbw�kT]!�lH`����: �.Ρ,���.����Ψ��J�h��;�4qo����mz$�u����+��q(�k�X� ���~�TD6c]N$ss'q(�������3��ӓ+]�l�W���M�z�՚���m�d�H4�"k�![\�4̬=�K�c�Iy�##Bv�+c�=в��`�Y�G��M�����̹��H�X?�6y�,�F�.L���R������h���8d�I�rh!$!�9㇋�,Q�}��;��4�N8�3��_K�q���+������k
��6���=Շ�O�r�sqZ�װ� �pU:=�����01��q/��<��$�mKt��ġ5"G�-���c�ʹ�n�s�N���js�V�`m�Ưuz1K�/$aS���Mc�$9ث�hK���Eϐ�4�v=E~ă?ǀq=� �y"?�*_˰�H���z�"9����VZ����Mtj���^P��Mt CL$-��#��0H�o���\�P
贠qlQ��p�DFr���
�x�+�A+��/�(�ġ�J�g�e=*�9����9�-��pvN�"u�E�ս�#�ql�%�3�5lRa���l�ʍ�$a+7�N �k	���f+퍃V ��e����3��m�*��<Vk&��%o��|ji8	�Ȉ�%^	�"YC�e,�Á�6aЎ�mL+�����][���X^���X�c��NE��U����u�{�V^��)�#zb#��&x��tTĹE�+�uS��u/_ϨF����IA�Sz��%~1O/|�XH��"c������rʝ�U��]�>���@�	0/�w�m�~�Q��������6(���Z����2t�������'�3���+�E����k�*�����D�ږ���𮄝]�:�4$!���k�tr��4^h�]v��D��~�����F�Z�X��|��m��H�'� A�1f��`�	Hn-��fa�P[�{��oܲ�h��ãrK�)���__���ɯ�
<����Fc��k>(Ry� �5�b��l��3�<�:2ାq'��b"�W��>�``M�G"l�|"�->�Õt�ߌ���BF<5O�v�oe�Z18�$e�=�yܓ�b��6���X�o����[F�㚶�q���\� �{��+��0�������q��q����1�Sp�)�i?f��IIK��q�z
�|��Azt[��6:d �dy����`貲��"��2X {w������3�!D$�$(�ꁿ�ʩJp`rj�M'H�4!*��q���I�<P�f��-���5�_7�m\kޣ*!��S�C���Kdq�������>D�UaK�u�F��̷@�����R�4�>0���G��ꦀ
��#���-����(@Y�_-�}�_����_�%�����h_��T�F�5'�L��Fn�7!W�4]'�Rp��-�fb�頶�.�q2SǓϊ��"bV�)�m�YK���S�?.A���:�W�|��� �Y���z�ǅ�3EJ�"�C
��@�xx����i`����ZL���ccP��ޞ��!5d!xV�Wj%����
K#Ԯ�Zo>��p�9K��%GD2XN Nd�>6�r1\A��:�Rgt���<[T3���m��ףqn;�,���(L��gUnԄ������G�t��fq�Z��&��SAY�T媼m~�J�+V�/3@Y�M���,��f_[��%5V=�y�W����f��1G��+`A�J[Id���	LZ�BHxVt���%�|lq/�	�B<z�$�	�l0��i������W���I�h�vz+���?X��=����+�B4,*J����E�,��G�VD���!��	�
ƃ��56���g}/�x��	(�U4��`4�������^��c]�
��\�_�%pJ�A�X9��AgzB❒r��M��\afm�f(?E니�_z��ݝ��.��z��C�P����	2����v_��Vv�vy��9����vo+'a��,ꖡ�e��LV�|�B��"F>� [-S[�'���`����+��0'N{5�+�����(�k8~����n����^a5�A%��,�p#����isu)(�DiO�k�ıڕ���㖌�nI�"�*x���P�m�����j��{����ݖ��pDDq��G{"r���=;�4~�C�T_ȧCM����\!�wr#�1����O�Q�Wiݮ�����Zl�i�a6>�*����b �.�l�] �I�㞝��G�8��H������G^HMC� F\��EՍ���NW���MUжZPJv̉+���54�ԁ���(k!M�+^T�;gH릈��pe;�ڤ;Qm�?}Z��/��]C[ۛ�����ܬ�?�P��QY;����J�j�V7��{�y�te�9���S���=�A��z�e{΄}�9{�������&��`�����wY�2 �]�q����5&3^�y�f���%Y7�(�]x|;!�=�^�4��Un�$��k�K������̷3�iB�C6����ylsxaLOZ³��z"���T<�뀍���Ћ2�����!�@��|�*��[��)�lg AIm@-�v'�	��a7����@͊��p�0�>�,���cX
���Z���.gDa������Ȯ3��t��3�~�`g�M�+(r��7$��]���K_�P��d�g���!��To��r�/Wv�bz}�`�����s�QR�@s:����o�S��k�:��ņ�eX=Ú@�49�b�zg�Q�>�����8-V�[\�=.^��f�%�;$��V�n�C���	a�a ���2/�?:�����?%{i��Di�f;�1�#������y�&^ӯlK�,�Xn������'4j��[F����������������}Pu��=� ��f����S"�G��� �R��_]ݱf�����M4~���ltcD��VRg	T����U"�����8�FN��\OQ�QZ����*�J�ʆ� ���/\vd����V��c&t�ْ
S;���Җy9�x?R'��諮d�4ڒ��Z�	�=��:hk|7�X1�_%��<�Ƞ��&#6_���@���e��.L�4Խ�MS����+)d�v�ckƣ�&uɱ�����t�kfo�`.������xv� ��׆�}C�|Z��6��.q+����3#vl	�3_�ꆅ0@F�|�%{gНz2�la���״��C�[̕���>����Q3�3೪��byZ!�@K�GX��,��52��sl�1{���;��O����~�7pf�0�Z�����j���4#�1hS�^K����*��o*ܹ�v>kS�B�w�b���,����r�X��t�s�7{(�[��87WL��r�A m8_�`�`�f;����;�Z>�O\�W#c/d����M~��gU8�5r�8U�7xw��+k�-�&���M%E�l��O�/�!��^��z�|*�e��ZM)���uC������I&�g~̵����G��c*K0�93����fl���UfV�i_��UuO^U}Po��1`݇h����q���3�*I�7�^kX��0���m[�>Y�����`Ĥ�qi�$ʽ�#2���Ʃ|�Uy������*�o�x�t���[��t
��c�stk�ME1�-yR�!z@��ĝx��1��_�8%��@l_��ӼsP��YӴ	G �Vb����)a�˝u�0�-?b�E�'"�d�;����!U�)굙�>��<u��r��B�r�h|b�y
m�%PJ<y<�B[�F�̤O"A��7l\)Tm�����0�>�8��d�%�+�^�)��))[���h�\���
b���1�s��dK��1��d�!~1Q"H$��h�QN ���p��{��(C��g�^�G� �:�����nA��|z��җ��ӣ�<C{hv��B��%+��c�(�A2�����';% ��ˊ����/an����,��fp�@�|]���7�Kd%R�#�:�f݅��pY�;��(�̢�G�-��w� N�!e@�j��k��H��{�Ҕ�r�ն?����:���)nVL�C��]ݡ^�?���1�k����V�K9h4�8�f�C�І�Fĵw�n�*�d�M�;���&���Y|�_������V�1��,�܂-�	v��Fh��Dx�sz�Ҥۛ�J�]����&��D?D�����9���~),�Q�&�K��X������%�������#�;��̴^�+\�2@����~��>s�ܯeP��K޶Ш�r�Ys�3̰4Ȃ2�}i���D�:��9��D-j��G2}%����e��ٝ8Ƽx�/Is�aLT���{�Yn�K"��}*�L�y4���G�~jI{��i9�P�F����в��=�)��a�N C��Й�~o4�~M>��׾w�%.�xg����w��#��H
L���1���f��U[�ށ�6����,���6x7cC6
�Rl���/"~��g� �z�dw�b�����a^$����3�����R�J�a���`���4����ZEа���&#Dg���^N ���{�H��������H5T+��	N�<Yq���:/�^�Jҥ
������d���^Ґ#o�9cXg����oɾr��?h�t��A�A�����e�0�y�5�-{���RPW�4��[#j�,�P���>��v��zdf�F�=��~��0���)ж�d��_�9�f�*�)`�3o1(�f~dE�Q��Q*H�)n�q�e/M�����)�I���v�t3)�v6����|��2�6r  ��#��KO��:t!J�ｅ��|б��M�O��IH���;�X*����n��rm+%�"}F��?S�:p�x�:���	��Z�[!�)j��D[?&3����4�d�����[^P���'���?�0��4:���"i�p�X�лV���O{��%G�:~�2�~g��NL��LJ�/ \@�]�z�(Rf����	��lr�"���T<߼�)�D��J�D�ώ�+�"��N=���n;�I�)��|K�?��#�	����`ǘz�еz�.NEmxD[6+����� j��>��97$Gm�l���� }U�rk�u�V�zi��z�?`OIDKե����^���������o���\9a{�:[3A�r�Z�5L��^���j,�x�q)_�UC�W\.�OT̩[���֭ -��J�3<f'N)��Q	
� p'c�=�(�SH��Tw	�B��(�|w?��*�مQ�R�{Y����r�*�����iqI��]n�f㶁� �1��Tf�-�F�scA%���]���4,HymK�+�ܡ>�=������w h���gCiMG<��o�+dj���ׇv_�"��[ �6L!P��z�Ѕ�x�2�2�������΄�ż�v�Vy ��3.�ܪ{�M5SV�[����E���)-Q��&1l8��l��"�q�M~f�juo�1���l����'�0u��%����0�[��S�ʿ�_��5�颏���%�2�|4��]�E�1����������6H�D�{q<����}TE��D;r�Q��,<]06���m���x�}\\j������U���r�q�`�A�uQ>A�b���ivFf㛮���8n�N�%��SE�������楷�UZHe��0��6�}M�a\$��B��_��t�P�~ɭ$$�r�J���2��~@�&�b�v�����6�G�k�Y 
d���ι�5ׁ�jk�ӓ��0<L�L��3�)oa��dJq����^�k�{��Ѵw�"�oTTS���N�������!���pm[.¦��S�q	E��R��Cƍrb�㥇t9��^8����#�L���7�9�ի0��FOxH�?�Ǩ5%�	���w�L�8��A�\mU�ƞ��^T�^M"��$Kg��e��сñU�]�.j���'[q��h���9T���ٴ��+&��qZؚ�I��{��%!g�l�a^4;�L�����w�����s��qg��}���9�Y��"���Y��/7�έˎ!(Lch�y*���e���R^��9_NL���$�p#��A��sQ�Qc��>���E9,�l���!�h�M|DY�ʁT���s޳��e_�
"���y0��Y�K�Ul��`�8�*w��ˢ�����tuD��q�v��/)�5L�u����X|r.��Qfc
��)�V���
3 �O���"�e�{���\Y�(�0�طE������P� ��QV5�M�!�c�J��R�˘4%g����� ���*\��؄�^RP��n�Wo�I��������x	ð�Q��o
�ϫ�}��1֩k�ubL"�3��r�[��]�1;��0q�o\������AO�$�0�R��)���:�K���v�m #�'/�qXqF9��׻@��lR���e��=�T���ϧ^q���
����}|�����=/܅5�=�;��x�lxj�
��ǡ��F,� ����x
��kHt��H@F�v��W>�,�WG	���v6�������^�~cF��$]̽���&�"�}	���2����ď��O��'hM�z'�<��˝
8hQ�|�!��jDt�,�.@wJ�\138Zf�'X�3�]����Ϋ�ux�#�5LqW���_G}�#빚�9*�Ȝ�0����ۜ����{fյe`v��\����S�����P�H'�m���Kj�4��aui���{[���i���t�j�!T����L�n�0�V;ؼh����^��P��ڙ�i�i�[��V���tr<u�A#�8�^�q`�f{cK�2�8�3�K�l�{Ǯڳ��	%u��ߘ���g�w��V:ί�6��0�&��Y/l+���B��B�b����p+��q�:,35��h�r������V���a�M���bҍ :u*��������|MsUW~��e%³��='�S�����s�R݋rEL�ݲ0��]лq�?�R���1�)^���Dtk���t�0�6"�р�9T�`?����;��-�@��P�.�/��?��#��Wc��h���59!q�²�x�T��P-f.^m���n�w�q�31S�s[��o�Ѷ23~����/��H�����V|MQ���X�BKg�(��V�{���q�q������I"2�H�=��W.����g�NL����� ��2"� �lK��H$�����AH��wJ���e��˱k%�P�7x�$�S�3���B��a��>��'��v����L#���>����q��ɑ�J6��+
���>,i;�C=xX�c����+&�܅���6_\�r�t_+���I�ooh](ʕp��ew�kٶ�ˢ8�vuq�k�P�*��M���^�,2L*�=Y�K>k}�u��(��hNm�D5>�éV���T�k3z\g�� ��콵��2i| ��Zsd�wlJ�w�Qy[6���ػq�?E_���΅�,�w㫥"SX�
]�+R�yO/ۂ��4E��h[�ݕ�������/t�����Q�ty����b-�W��,��C�>�Do�̰5)��Ԛj�R#�{ 81�7�T�|OLΏ~�1�$��YԂ�;���B�sk�y��rw�}����84	z������X�JB�sk��/�8��Ѭt2�a�����0�o�$�Y���p
�yߨ��QG���H�Ȩ!p��){�{��q ���(CU�����ͮ$3�Bp����U^�=<�F�>Q��Jo�e88͋��J�$��C�*]Y�,$V��Ig:�ˬ|����;�FO��H��a$�SJ�6U�F�ܻ���ȧ����6K�M�ۆvUT.GB�F�FY�d�Vo Β��Lȇ'�� �����匫J����?H+��N�[�8Z0�� ��"����Yi���H�ӡ������)2wH.7T=w�r ���p�=�Fm�x�
��ѿ�H��c��`���O��z>P܈{��cu
L����$)L�W�fн�T{�?�����{��P݊��27�7sP���¯�g���us ��s���mʭ�V��� l�'��?&����f�*/֓�vX�P���K�)����M�\9l��|�I-?��k�tPD�fSU�J_�����y�,3�C�F��\)�Rd �f�AH;�du���.�l��V�eh[�ן=���rvq~�wR�V'�����ط����E�`�o۵΄�Ǩv����d��0��}���+��b>V|s�όF�.��^��YJ����Ί���x<��8��M�i�N ��{w-@��0���2����}���q����C�O�A�5Ԙ�ԣSlb�U�J͒Gz�Uں�8�@���$��Q��k���+|'ͮ��9,2�odtE�v��6�a���ee{���49w���[G%9�՟�H�d���_(I/F�{D��Κ��{QT"��O
����P+ Uv�"��^�GpL�ä��֖��Z��+�$�uҀp�,�"����Nc��(&�H��V�_��{�h��Y�~� ��*��%b�K��T}9 |2�@R.������ۀ`9φ�y{>�,mv&xf�q��%�\g��)�� �GǏ7�ؙજ�q��*��󲲀�6|]�����u�M�1�J_��/ME��
�~.P��FV	e�1�-��p�V�K>�󀑖���I"<�.��.��3{)�hI�S�B�6�\Iu��
^�(�ɘ\���L{�ŧ�?������s!��=V,y[V��í���~-�;	��:����ʤ�O}�S� �s'1c�kc�˛SJj;Vi�A��F��E�>]D��q_*n�L+4JaC>h�\Ei����'���-g�ŵޭ���c+�� ���xD9�Gyڷe���B����x*K�!:>�dP��,�,d���@��?v_��
Y�4!�i��
��Wy�t[ƿvm@@��/���f��S`�Əd���Yh&��5��������Նڼ���a�`g�m��ܲo���gN1����?�m�-?)��"5�k,����*)p������;�r5����g�x�T��2���>���]˂j���4)/P��tM,�VKW�ˉ��Sՠ� �~J�f�xK�?��bFpg�/:z3���������d�.�L�?�y��ĺ2��׼)dLf���6�g�M��k=G�~X�{�P�W΂�ŜPo�"����淃�eE=>�{�����bq(�m*�{W8�n� �OgU�t�Е
�t���)I� ��}h*(N�Ź$Y�v�r]���0B}�*+�.�$�[���}�a��-D��LN��4z�L��֪Bs3�GD�VF�S�Ġn�˕�_{T4=�-�eɮ�}K2���!=���v	߁�������@g��e	���i��Z�l��<
�Ģ��6b�����B&`-�m��NQ�:v\��ar�/��fS��̴����~3�ȓ7��mڝz*���C+�:�Hq
�([�j��E�v��҄ÆJK�B��O�y1 �i7�R! hE�(�-ił���Y���Ա�-[�m��ڐ��I>2��:&��kÌ��T��y�]��G�(⎷�����2Uc#�X��?Oܳ�����ɖ8X�Rq�"1C�
b���1��}�ю��U������&��]!�8�\%
�&�=l|�7h��ηc�H��7�����9�^�.�푽�@���^?�9�Z��M���y�26_q�@��ڪ8����qY�:�
3A�]�P��3Vz�Q%�ؿ�#�$+��B02-��8����շJ�Ԙ^�V�� �3U:g�Q��V����u��-����zne�U	�efJ��lQ2�] �p�V/�98�f�$�������`��2���F�Ca��D�����)���	Ջ�����)��ؖ���`��z"�.n�f�D�
1{{���E�8�`�;\ ul���O�C��b��qdi���󒵎=���<E��/37
���{��Ul�BEH�cn��t�A��5�
����j~��<4��$�.�
<�cP�?B~�I�?�慸Wz D=2_�d% <������pI�w�h��;��A�1,۴�	�g���Wf��OT5��0��f�\��a�;T��bB<1��� |09�%�	sy�\O{#� m�72�WOC
��1�R7L2��1�<C_��,NdY��o-����nsS�N���k�����F������?Q������6v!"C��Ow�/�0���A�c����YpdcS)_F	����µpZ< v\D�$x{�a�D&b���~���@�e�;�O1��@-.%D�:��E��K�a�
5�9:�i�+&����b��W�b���f5�]����qx���U���B�����9�/)z���X����)��R��,/7h�@�a�XBB`�:��^p��D�Ȉ�������*zV�w�Y^#d:o�_;�|��=w_mQtac����{P<��7Q*<`h�{ֵ�zۅ��'�_��ꔧ��E�}x�%Y����x�gW-���}[ecm��*D��_�tqz�_��b�O�L7��Iiy�bp�A�zj�S.JѤ�'[F�ok-حĴ,�`��"��ަ�p��NfÐL���"��Ю�>���0^��&��N�*�����I�f�uX�ʞɪV�S��C{�9&L&��L�?�"�O�����0)2�����
�/�Dˎ�&�&XT��]NbZ%���E��Xa�&P�=(s���k�ԯ���l�C
.� \3g�Wm� Y��6�� ��#ۃ��۔�0.�q��k	5�_|���u��!�MY���z�,�b�  Fp^~�2�n�|]cRA�����U�֮�Ժ!��/���X�+��߷D���t?�� ƈ��S���p9�p�L���;Z_dE���;�\"=���!?/`�� ��l�%��۱��kPqgj�f�X������� ����3�T{L>X|���+̝R�����:��n��k������cl��:뵚I<a����1u7H2�YK��{�z�ϓ'��b@�% ������fm���x���9�!��#E|;�>�xRpʜ8r*��C����]7�r��?�E�%ϊs
5-�b�s��U�T@b\ZOT6]����<�
�V1|�"� ��T���c��Y��l����4}E�g_+( ��.�q���u��u-G����$���ﻹ���!4�C}p��U#�Z'u�q<,{�ѵ��7�[rp8(���@��g<9g��� �>��@�v�Q��|NE;��P��<-ױ�Y"�a�09��ag�c�����U�G��4���[Dw�w\z�V�mI�6�크�Ԙ��-VEi�D��2�㋂�i�4qz�w��7��2v�s�נrUZ�H�Y&��G���]��O��DkxG���;18)V��L�[l��¯�M%����n���G#U����1I�Wj�����+��ަYZO��~���-d��ӡ����)�A��"�q'�(�?�җ�]ɸ(�\x_�?{*bP�?�eܕ�o0�]���0W�_[,��.bE�z�O����~��F7ȭ;Q�bW7j�v�h���2���'|�5F!��8���< ����:���aT~�\e �̇�ǭ�<iF��v���wzg헗���� �,>5L��dY�O��5��P�?f�G�,�&�İ����+��_�<����t���A�d�4N��/u��X�v��z��p6��& x�Ax�2$���h�iR���㎖��׾��n}��n�,%�ƞ������5��R�G���(��\��S�m���!�ui=a ���w��Eْ��#|�@��c>j܋��4�z07��s�L#�0��ִ��̅+�*ϸ//Y-�1�4e��Ű�IYТ�ɀ���ȋ8����]�=���j�4/���]���4|�8�0n���R�⟣Şpa�}���$���KC(��XβG*���)�0R��+�!���/lPŮR�(|(=�@b���nk~m����U��kT&q��؅���7Ixax�5oG:ɏ��Q�,�'J��^���%�#��*�?f]s�P���.	Oh��dQC���֧S:��x0+�[�K���Ό�$��u\]�Q��U0��\�"�X� 	YrbכRѨ��� �h����b���&�A�E�Vd������ͳ��&�uE}�L\E%D�-��	]��͖�Q�I�R�n�]���o?��/KT��e�pA�~�^"&��O[s
E�H�Č˖�ܳ��X�}�3�#~��_16ɈD���]i�����i!(6H��jҼ:�'�Y���P�L���C������?���r,�1��^���T�W ��ho>q��%���pv�G�v���hϕpÚh�CK�-	NF�+��Cf���~��ݏԗ�Q���ɀ��H�z��*}�)��u�z�#%e�y�[{�RF���&ݸ�ӅV)�͐.d���G�Z�!���S�/!]V��$���+a�$!�>
-��#�z�����f�6��҃�k^�}=��I��83Je"1<[���"�Ve!�2-ߪ��Y�ӞxHK��P�K�����p�p�&Ι;y���)i�)D�3W�E%��0����e���Cf/���pL%�l�
�A���w^d�P5���e �n���g�ӠfuX0�	�(�3�pJ�F�X�3�C_���]T՜�q4`v�;�o~X
�x]R�t�ţ�%��6�F_J��Q�w8 ;�Ȼ��v�+�#���`�˗��v�ECI�L���jC�}s�N�t6��x졟�e��$'�hp�4ھq�T�Ue����(���ޝ�(,�-�V��@5��r�^ȇ=E�_�U�Bz�|�W���2A��t8�H�=���>VT�t$��3��9z���~g���U#�t�ԟ�����^���Ġ�����t9?�Z�!~oȵf��.�F�r�6�X���C�u4�;�':E|Q?)�u����b��	�p�����3�	��R��������%԰9���'r�RA�D���E� 9���[�]�#Rn�]E5�F����s����"I���
s��Z�F��;H�n�v�����6%�p�K��J���FdcUً.'֮��m�vQ�X�;��z����J��1�K��XRw\D&����f�}o0�b"�v e�feX�͖ *��p�.���o&�Ɋ�Ny��Lw�ҴI�o��k��w���)��V.,��up����*J�8���R+68�#�`�ʜ�����՚(������o���t졼�%V�o�\�7L�)|zФ��ܠW�4|ʹj��y*��ľ�~�[��Y%�D�7*�,}
�����W �BlxJ��df/ߧ��>+zH��[�%G,��Y��J�<%��$���;A�N1�Z}���i)9!�n��RL�O8k�7�[�j�|f6�M!��O�pZ�R/�V�bL���D9��,QT0�{���x$C=�k-$	|�P�lm�$E���l\��O]ގ�Yz��k��:r�h�&،��d��h��������(�Rrq����� �	�ݮ�q��`E�ʫ=b۠�������>a5�b�g�5��r
d?�;o(�1:�Ge���1!�k��0�\<Ҵz5�=L��l�f^=�q��e���'w�d������Ԍ�]dP\��2sX?f�פh�Ke��҆?��[�X?$CU>�A��[x�޸1�P��w��Cx���kn�ja��s	D�R�� D4CHz����k2.m�����n��
�$����G��A��;z��GO�����[�����v����g�ȁ�������&ʰ�i�����W��H������3�g~�=w��K}��7 _���D#ͣ���H����ʙA4ڽ?��>��'�c(��������q�voB$uW�;�{,O5� �Hkj�=�y�%ܩ?�����, W#ْ�	���M!O��:�:��n�����gݼ	��5�Dr�Z	�U]�]<�0�~����LZ� +&�M�ۯ��![讗��I����N^)�F�QTҐ�����/�e��8�Ǝ����R���S�P���������CX,�	N(��av���4m�4���[jf(X��Ͼ؁��T�*�_�c���m�Ԝ�qn�*�o��!gl|��������&IŖ��uum�w(��C�.��*_*�Ln3-����p�?R��Z/�`��6�淍8�v���w�[˕�=�'ì5��,/bYd@�?�M$������=�$#_\��m�8=���\&ǜ\X�y�Z�X�Ss��E^ׇ͐����e��(i�h3�Υ��ܱgd�\�ؗd�G#�� ����G��C���i]���g�Ke���70O ���̈m�X�rb���lĵ�ӳ�T�P3��?7��`����Z^� �{�&�<�*�c3M�7!,%��-�K��+ W�kQ��#]����E�U�(�� �N���%��l�U&F��U��<�C���a�Jۂ��Q:b����]�hMW�t���t�����4�[r4�1<f`��3���\X`ww�%F�K$n%��!"Qq�NFgg�uM�غ��qc����洓�����c������[��b��<���d&P��j�Ę�~�N�~il�c�a/�%A�$.�"����;�9�oCE�w(���:�͸,�c�
���rF�8�?&�~��sw�y�z�[�����:3�7�6>T�pϋZ�MBU'�ޞ�YCQ��~�E�� U���rj$(`�&���5�plG�����H�	쥉|0^clø���r %�JJv
��oY4�`���ĈY��w�멸� ������jE!��@�2���v�w���o+K�{�bDaw)��;�S���m�<� 2���^4������U���Z�9y�?�2�A:ƹF#	���CZ��w�q86���5fm��jm&+��Sy��KxR��D��N��>���QE���]��v̳S�BQ��
�lIc���54"�`�V	W	�4��#UmF�j�є��z�.��7�5J���-ZZK�D�i�6?hSt<��7:1���J��QJ����O6����k�����O�1A�~���r��%��>�!'U�#R1|����مyK�\����G�p���>��P�f�$j����}ܻ\nVʣ�x�қ|����C� �f��C�ƧV�����n[˴N��S|��i�`9�P�nø�󈶜�ʣw��-����szOAߊ&���.�**p��둈=��@�,D�u~x@	�����>y���[}��{T���Y�I>-��
�]�2����0�f�C��#���1Xo�ܑ*[L.�}o�ޝ�#GE6�ֺ�+h�Y+%�d[m2Z�vE�?�����m̩��+��:�n]��eZK�����e����V�xZ���?$HK�b���r�Cͥ���#����,�`��p��0��\�A�&��ǣ��b'��Ɛo[Q���4��#�|K�6~��7���Q۝+�_ɂC��I��,�x?P[F�H l�����Z0�Cq�k��ZN�˶N��E�̨��R�bC)Y�B���q��fS6�kB�*'d�e�����7�z��Uh�~�,�S"x�l^a��J�����{� H,ic�o��W����B�(?�L���23Z��SP��Z>����u���f�s��� ��Q�<�Be1[����}�8;d`6$�.L/��iӫ��a��}Ju�Q?y�����T��I�G������Q.������>�5��q� ,����:��D!F q�ZD�� ����9���]X/�H��Ǡ�����m~U�(y�F;p�����O}'��f��; O������ ����fo�b5sL�ۑ���������'�َ��a�+��[�W����&׼g��uA}�+l'9�r�`g�Hz�!�fŕ
�0x�_:�'��*����ϭ��^��Ү}���ɂ8�R�������3C�DS6���k(�����j��r�@��M��3�J��^��͹N�ns�-�E"C^w{��*9 �W.�����aNX����"�6���*��/z����P�eAs���G����pb���U�����k��������%�ц�T���G���I§�$�����
��0A���I3�\D+.�$!�{=�q~h���:�,��Z���?��w�W���(.��� �#����6�`�Q��&o2��Be�}��jʆ�Pb^��Ҁ�ؖ;h��� ����kM��Z�Ǹ!p�m�sϷ���;
�-UkQ���潽������v�F�M�� ���9����p�;oM'�^�rj���&�� �p���|#���p/�h��{���cS׆���D���x	�	:��dX�<>
�%r�r�1H9޿��3,�sJ�ȷzf���T�"���ڴ�d<yV� ��U�LP�:�j��ɦ�`���ٙ�#��gJ�O��!`�i?`p[��~�A_�l}�k|��e8O�*��h�=���[��E��k�E&c�����
�8��8�^de�g{L��FP˩ML
���?6ƒ@�2�i��>K�ww�k�&�I��s�~S%�]'�P�/N����A,�؋���]}��k��W�#PN��U��L~�����6G���h]�O؝�2�P�F�� UF;�����*|�s�ИsMP�z���z%d��!����O	��g����вnsk� ��J0?�d�T����}�2��
��SL]2Bt;J"ݯ`٩Hl�}A���۷ۼs����hz�O m�(����09���G�����o�w�Q�;Ce��q���~��Qu���S����!JT�{�����t��|o f�
̨����A�s��&�:��ΕY
Q�s�-��flեk��w�k��x~K_��ڽ���p�a��" N�%AJ�he�����N?@�64�+����p�:�������H��+b��t��rpӫ��ߌJ ~�������Xe�gudI��	#A21����`)�	e1�%��+L�e��+#{y����:v�>pf�Z�
��Kz�J�j���T癗aD��g������yS���ۂ��lJ��(뉋�LV�;�t��A[�qL�:G��o���c,�=қ����U�{�ř�g�B�u<Vğ�"��y��@�>�	���X~O�T٬�m0!f���D⪋�B

�;®76�{�VG��Gĭ�[H�v��h>�N���z-���fx�U��!*��\��ӆ�?���Μ�P�b-�_��E��\j�P��e�eZ-�)���It�om��wZ{]����pm��\m܍>�dy����A%UMh^�r��w>����a�(���
��gt���?����0�a�&C����T'}S/l�)�|i��`�K�.��L��iÍ���g�DE�zN���u��V�~^e��LZf�-K�b5I�0A�W3q���$q��6ڿ�Z��S�M�G���{���v�s4W�p����w�}J���Vpd��a~DQ�X�����ٌ鲤KV2aBnc�֚��8��YI�i�&r��>Z^��س�-��vp�2k)���7�n�8;2��En�B�V�O��b2p�bj��_*�s?���0C��~�KVv�Ls�U�^o��ݲ����R�y���{�e����27l�Co���]�_5�|o[��d��� 1���P���AL
q�%�(B�;p%<����k����EΙ%�J66@�7]L�"z4�OU^�дl����(�Ԓ����|�e���&��k%��F_���z�~b��;�˫>�qӭK�����By W=
���EV+5L�F��xn����T�*�&�ѿ"~I�N߀��zt���x�Y]���^z��L���۟�����,xđ��vZ�3�{� �/D/0R�בfؑ�lp".pz��REu�k.�����lL G
��x���'�U`z&��
�ɡ2t�W���bȣ���z���w�q�A�p������ׇV��Y1L����<�ӌ��q*�jR�W�¨���`z�n�H8���\����Ц�� ���ά��s�t���On��<��桼=<QO	mM?`�_��
�"N��q)9T<��Qa�'0�&�6KB��#,���ų���`v$��!���yI{�BA\��;�]��4�h&�Vկ�� �%k�����]�O�;Lg�pg���C:�x�9���ó娮����zt�G�m��z{�����0��˂�'�;�V��4,Y7w�1Eːs3.c[��a{�R����1�<�n3��gt��$��*O�ܸ烺�i�g�/�LQ�����J���
83���b�m��d���%��Ӆ��ď焔Ό��C0���5��3�;H�d«�wsP��8w��pp&��e��hW���Aօ�]�C�7�f7�D�.w90&��;�3��H��ׂ��@�:T���e��ZB�����_�`�U�ZGr+rQ!�4���`�"~�Oˌ�z���n��+�T����4�j�̌��h��:�)�X
n�����#Kϥ{視�ٹC�X�Ȣ���0���B�Q?x���J����.�Eץ&4�BMM��Ɨ���X��w�!�O��r9�KEx��ʻU]L�5��~7te@.u�X�����}��v�O��ld�CaY��#��K�u	Q�C�
�J��)7BuQ��䓢UOP��C�1��Qߣ�E*R��'�MW�9���,%^���Y��z�x�e����?�9<-4ƽ[^#�#��0�~�u7$Z���f�mԢ� �6TѲ�_���	I{� ���>�]&k.ş*\��F�Z9KZ;x�~偏eeG������
,����̀z��:k���l�Ѵe���?<�D/�`o�M�"}�P�T����!�["�6%�v��E�3jēw,	�_�R#�Mt����:m)�I���e٧Ӟ�u�$�_�$�X�!���o���S��,ci�Ԉ��;�r�O��$��n��	��$�í�w1%�-fE�b�<S��{t�`�'q�j�gG���4@��hc���ء��C� �%8��{�
]���z�+��'v��x�H����%c��uo���?K�����(*F��iz�)|wi��sͼ���	�Ŝ���)�irZ��9 ��Ӹ��4�h�k���߫�k۝�7E��m���e�Y �"o&#�@���?�:�Ff��<���e�-�I3��j�0�B��C������-��Z�4�`ek���٤S��`�������P[�ND�u��+G�&gBF
%-	�j�X�]+�)�����g�������Ļy��@���\��U��"{��"��Tou䮠��>#�ӈa+�k�����S�G�2�v	��:W'��z��On�����~��>�����6�U���$���-�Z�T�]<�C��F��L�$@�F����:������)lw=��0y�@���֙�����Kɏe�l��sR-����{6��&:$8wp���g�?D �V!_���'���n��A�0�;=po=�C��x���Mr5���;,��̰#ͤ�;�@�K�Т�c���U�BՔ��ǖ�j��|�T5���Ԃ8�rc�s�O*D��ϸ�Ply|!L��]�"�7�f�N��d����(�*��"<�pV��G ��&��$�6��9h
�j��,����@�}Y_�Yi�E�����Q[7��Ѷ�d߹��3j���!{�9�u}�_�N��
���I��rX��R%�*��R%��H�����YS˗����-V� �eH���R�9�ϊ���(mB)���U�&J�J!�:��!j0���C��Wok��97^�����mĔ�+�$�~�)��{O X}/G��Uu�P
��G�l�I-����ҿ�(�d�f��	����\����S^�� $y[Aί��W�<$e\q(���{	s+�>�%�ݵ5���K��/���y�x�<��,�xD����˺%8�8s/ |*g�$E���M��a�I���D�uȺP�N���\�x�u�K�|������A���'I�M�'Zj�����Y�瑖뉊3V�J��ň4�>"d3�r��<����,�D.����E4g_
�&�k���O��qw���qF$�C��Or8�q��(��^���:(E�3a#��l�yZ�n /�^��},��l?.s�qhPn�j+��(��$Ux�\�d�eK6�� ����K���&�t�ղ:	%"R��A	WlL���Z;Jm~.mӸ����e���\z�E�)f� 5i�h[�+�Rm�����$�]��)�@�;~�� 2Cy��ݟ�+����^a���sL�DrU���j���n�t%Z��-F���W�ܼ�j�'��M
W�L
�S����l���(��S�����WH�.dQ $_h>>�BVTpJ����w�����FZ5$f;??u�7�X P�.�����(D�3��V����:K]�4���0Ԣ��ӿ���8��i��^�>E>QJv	RxҬ���R����a�vs������2>ᕓ�H���u M��Jz�}�PT̾0
�t���̗���֣nT�1� �������W�7A�Gij%�uMƞ��,�}c�3E�gdJ���d�˙O��|
4u�)9��n�&Q��u96�m�� ���.A	�vǊ8~�J�|��?��[H�� r���#P�`����]��z���{��wX�U�D��Otw<��ğ�֩�Ӱ'-ʏi!�,��0�˿��rko%
�^������vJ]6,�E�����Zd�-x"H�黿�gP�q��d#��¶s�i�\D!CП��N�6��ܐ��@,|��!MA�R,+�e�S(\��������X�ZKY*���1�w1�]��)sN�����7}��:��Pm��h�w\�-�y�����B�kt%Q�f�![�΀�}����v�O�;Y�@�1}X2`�SA�^~��-����i)+�qGr������(�kP�4��B��#��n-�� �S���6�7V�h��t�:��iMT3l��'̍��dRL��JU4�8�c��Eā�ʓmj��B�#�e����nN�ai�ڊ|@��F�4��|]�MB�3iڔ�§�(����������#�G�lkr���CY�f̵
�E��]�qGڶB��Щ���&?�1v�(�]��sm7xw�YW��_�|ë��G�R�]CV�'��Jꄚ�-���au`T)��W�$<��1��(� �s�G�%�V1p&#�NZ��(�4*QZ�J���6fQEWI�N��(�dX�;v�/����T�#����H���j'�?w�^�i�n��UC|�uڰd�����i�rp1�ή���>NJR�U[͏ ���㞫�+�{�@�V�II9�/�]jF8��9��N�Qb8��,�$J1��5��[m>	�x�7�������Ⓡ��������Վ�(�J����W����E�����
T:}�{�A[�jOk	�K�P���"����<�ut�����N4�ܶ�ԕ�֣ρ�?������`��Z�=�dc�V�#�[�e������&���yy%�������t�'�P
LY��Ϥ�,E2�����Oau���r��8YH��[}�VQ�פX����ʬo���ll��R�7:����z.��W���8;�.1����ma�+����)J�u�(�w4T�wN���րDY�W�ڮ��gyF�-�8����</Sx{y��a�v�(yXBJ�qM�=�XI��n}j�-��ś��^�1�$�E9�9ڧ�Q�Yqj�K26p����̨���O7��u��V�6��R�����l�'W��Hӝ�*2M��r�oh��`�G��q�]U�i�*�R�n��+V���ܕ9�g�1�Yv�wR��� W��(��ҋv3Z÷���-Z�՚u�lFd&�(Ԑ64�N�w/g��h��DW���_����ô���)�Zs9Y�RC�DV[W^����+�R��L�]��xg�*�$2;�b�i� �>�f�w�66�q$R9$ݖ�\�� A{~�Z�uy��=���,� 2��"��z�g��Y	�< ���d����f�j�Re�S��>C���#�3��+8f�g��ӤqB�d���c<0K�q���P�IU��@�;,��"�T�����ܚ��%�9���^rr�
3e �h` ��2Z3�J��:�#�,A�B�K�*�H,a 6�B�ݬ�W�3Ũ��6~�X�z��im(�]�;�	�]ыw^�v=mыi8�0E���I�Ý���#<7n�_��FE�ˏ¼:=A-���s�3��re�M���`��('|Y�Q��v(�
���9�0}��A[C�[��|����pZ�]�����uީ���	/�u��2?Dʨ���r[Yפ�w��Y���Yl, ��;�4'��#`���a;���;A澔3�<^�U��>�^���*�5o�����r�{�b�u69܀�� $F}Z���௷��t!�,��²�z��e�l@,�2�L�9^�*�H�6�;��D�tAa� �f�8��]	y��=�k��q�Ȃ�)�GI$���� ��{&���+#5`k�!�Z��?��c�ו�F!:CV���oT��p���L�y�a��))!�]����s���������̓x��RU��ȓ/e|.xW�_vK]�2��^w���tjQ|D5to�kn�UqO!�^�F�XQ��c����b�j��%M��n�mD7e�r����)�����$A�ZN�pÏ���o������0���|�����#���lٰ}���/�`XOɎ�z��ř�ӯ4��|~�%�ޖXD͈��簢����f�X��b��d%��	�٧�C���9�_;	��{�v���0ӱ��`h�b<0Ud�+�=� J�����F�F����I�m�b�lQ�,�@6X���*�WgKE�������/��� 
_5/�bkH��E�K�߼����[��L�oCɚ-%�?��}\x�EȨz�
�Lf	�9(�x��t�9�Od��aH.B,Q�ٺP��'t=񯰚?�L$H�((9D�=t��^]��M�{�
n .�1T� ���:��D>���nt}������M5�����{���Q�z�ı�Q�П�)H<w��q|���\�MH��5����s���H4	����<����ڶZu#�Jy�,����j�G/.Q���jT3��3�{��?�MOS�Y�#7'�enB~�|���dݡ��?|��+*��#O@��ݲ	��N 26N}�),�;�=h{���g�Ϡ݊���3�,�� =��W��	{��7?�� ��eM������zn�K���@P���L�%�����C#�n}�F�x�=! ���2�l�r�tp��V��z��#�CD�]V�_/n��z�ن>�>���&v�*p��I�g?��m��#~߮bS�w�� ��	������%����o�L	s�����}��8�(hY��"��{b>pL����S��?�lr�t�l��~�A�ދz�8���F��4/�`�Q@)c�F���v�=��f��;��ݵ��x�?-ٖ���YC�P�}����!��4��A���+Bj`�2���^�Z�yZ�{�
v߬8�ۻ�C��J��T�����]Q�n<����;�5 ��ˤ�G�]t�V�0�	;j'������S|�I=L�
#�h���M����V<B0��!��(%����8��MBl˙���Ge�;#`mM4`p�����o��S��9:����MBW������r�CuJ�%߿J�#;�]ԉ9�<��Gi�I@�٘@xw"՞ZBFDj{� �=��3ݴ�Ⰼ�/Ƀv��d1��Vm��l�2�D��@�����ew�@a���)GZfm��cT�C\��ȳ��̯�����k5�h��3u�%J���̴֥b�o��Yip�RщF�<���w���d|q��]��]�΍�0��މ>�ES��b�����@ؿ|Q����D��	h�(�#�E�}�h�DF�V:1A���� -Cs{^�%=KW���˦�9 "���/�5P�}���4�����^2=2]]�hT2��r��Z��s�E.n��n<��Լ��;Ԥs.��c��d���u�����%p��ǐ���,�2Tï�T�NG�.A����O�V��Ġ٨�Ͳ�\;R^.@FjW�m��l�ծ@/չ�&���X>t��>d��L��Ȭ�����<B�:�߄[6�B7�~�J��]*��+�k.E�Z����sX�h��l���}�b�3�h���e�6t����,�_��� ��l=�|�H{�)y��ڏ����w��p4D�6ڎ�P	����Z�L�U�O��U��8�T�.4�4K�ӝ<�(����Xm�S������F ��h�/�*}7A�I�ޣ�)�wKr�GT�0Z$L������.Ag_ǣ��1�������Ik������ָ#���I$��,Ӡ�Y��T��tż�;�ȯ�oAmsyb�+X��,2',������������5f16��z���nj�Y�1��V�	9�>[\�1"�c��2�jd�S���S�_ٶ�`�LEf�������ߥ�"�����떉� mb/@
ns����&E�_L�<����l{���te��"ft�|P9����\�},4�ᵤ_����k�T��3V�aJ���p��z�/���n������)�^UY2������k���7���Ņ���.r �"C��錘��{.���)ؘ��:����畂]%��S�B���ρ/7�DN��4�(�ў�˹�k�ĵ?0��3o�	��	k�.�qI�\ e���|��8���H�02��YE�XM��E@cΦ�}�x���q�S�*�?Q-ḧ�>����(���(Bk�^��J���-�g�D_���@���r��4�'��f:r.���`_QC=��e��pQ~�ąՆ�ւef�Z���5���@v00���HSp��"t[�s�	Vk���=�<�ȟ��Q����^�T�JC�G~i��O���/��ܒ��x����YxR��]���P}��&�wh��'�&F;Y�f8�m�T[���%hpN�Jj�N�oX؏��~���n��0��:;��������k�v��\��w�����SL�����^�X����N3���R�r05��"8"�o�'fJ��3����~�ƣ�d���1"~���"�~Y�>��C�{&�,Z��v��Jy�W7�ZnZd���#�_N���Z>.~��AVn�����Lv���~v��&�40��cRO�nW(`����Tg1��5O�R��n�6��{��'���#�5`��XV�\(9i_���F�V�?��	J4P}����~ް ?��P�[���;
�3
�!S}@���"�{�&Uc����擬�޸`^)])��k)ذ{����É��k�])Hc���v��p&�����nF���q���Th6B��媢ٗ�(,��\1$"b��[�g`�m���6�_�?27��a�H��VC��44��[�nG���ׅ�Zg��['��\�i_o��NA�@m
X�0w�i��r`�-^������ݜV|B�KF�륦���sSc=��v1�!l2b�wj�ZG(܃/��FĽ��
�yH�rIH>u��;+�b��mɈޑ�g8���y
b=�J��- t!��P9B\\������ԠK�G���ɬt� aɍ���EX��a*r5ƦK�j�o���	K��3&�r�w}7�"�����歉z��5�^��q#$�������:!B��������<&�c�<�\�>�!� ��J�J$�\��� �(j]I6^����=��.>��S��n��>��+4�#�%a�'����ݏ���n���H'�ߊ1�����M)��e<t�gu��,�K��T��'[��xr��\���W�L�&s���g���8�6[�-�!7=�Ʋ��c�0c�[9�3�>�߃w>I	`^tgi�
�E|n�ghShF�i����4Q-���m����q�����z���~�bSUwEm���H�&���W{8L�.���C�w�����yN����?�����h��-���m[:�>x8�F�sKK�@�ҕt��W;2�7z�e.29J�n���.NC�U�\��c)��炬_,X��)��T؅U��&�x�^�n�,�6͔l&��F�M�h�#�\P���*O~�hA�QI�m���
���x"��E\�6%Dnk��+z*60���y���hb�6�����zV���~��S*��K)smLSj62�n
�W�P�z�\+gYG�a,ǻ �K"���9f���Y�}R�{����`C�&X��'�ъ'��M�i!� e�6a��Ax����w$x��WW$��ϋ0Y����@���JS�Hj6��c�R�r�t��i��*�s��ݫ�R ?�I']Ӣ���Q��WbHe�!J�
�1�������e��� 3a-�_^)�2�>����
��cӄ>,����ͬ�Z��6�T"t�:;�����g�#GV><�ܙ�Qx�u3� �oٕ<�I2�v*�{�6�WF7�w�82�����wdǼ;�C���!��� en����㤐L�����5��-e|V��P`�=��m��w�%9s�����ş�?�1-�F�ԅ�~o���7�M��b�Ͳʠ��Mmy�7�+�N�a�ç�=�1�����Q�)J�[mP#��v~Z�rȞןd�4Sa����K�����Mv`qH/�'�H�?[_��J>�r]5��N�`��n�/|1{V�!��I��\���3�*T��1�r�S�2]��m	�� ��l��MTp��4EZz���jE?��r
 ��7�����t�NM�)5j�%C�`�D6�E�C��eڱ�Ѿ������"���nI�1'��竻�~�����bJ�3k�T�p}�>�1�Na"��{g��~��/�ɝ�|�n�����m:(N�\%�A��	2��K���E��H���sm�vOQ;����(�&9=e?�=�O�;���+Y%	<�k(���F`޻t�ܖM�l���1�֎��$n>R�M�V��vֳ9�&����jQ@t%Qw��.wpe��l�0�]�ޚf-�󹱎wDM��\<��r+o��R�ʬ�E4[��l�_�y����"̽��,��Xvz�?$Sd��Ɍ����J���w���
�y]�E��:�`�Q�\��X�pծI�-�k��3D�<z	�q]���qB�E��~�'��� �qe0f�h�vVE�[B@�/�^�����Gu����b=�}h5՞����0�KO����n�ϐ�}�)<��e{!�5s
<�;B�#H ��#���it�1��.�?��b��M,}t,�ƞB}��p9}~�31�m1QQlY���y;��į�DK5�����Q�<�O���0�<�wC�.4pUA��tܑ/�]��}��U�A�H[���Ѭ�;�E8�f^��E*���8�`�Y�gP1_F$�a��'��3�gC3�--��b����'@�T��	2��6���k�T��p�Z�͋�xg$�B�FM`w���U�G>Zz�-	op�����q�[�Ոnrܝ���!��qЃv�� cر^��#I:|4�Y<�e&x)!�#�k#�ŚX���Q<r��2���n-������Z>jt�3\�^sIۜ[�aB��<COm2�x����0�JEӧC;i�9�3���%��z�Mg&�j�ۈ�4�-mR�D��`�����?�;�cɁ��_�E��������~�S뀙��y��3�^��˛1�qY��Ń@���nC�廰 ��MA��V�e�z��P���&�w&0��]��OM����`CzZ�}D��ԙ<ꊷփK�ޔ�Bd�Ú�}���s>��h��2M�˧s+D��͵����>^�Y�qX�rЁR*&ڼB��t���lt�ݸY�%�ź��Au6�_����O�aH4|�ˬ\Aw��P�?�9p* n�� 2��~,e���e�M_nʶ��YFU&�z�Y��{��e��%$&�~�nq���?��乹��D��n��2�����DV���p�O�RT�ր���Gr�`7~/�Ͻ��(f~��`�mU��
��"���Y�A��r*�Q~�z�&ٜVf�^A��xƞ��
m�ZMNw�m�N�d��;��8�!�d�pּ�@��׮'�.�F���[��������{[�������ͽ��fġy&�_�H�U�ܶ��XG��IP�2ׅ�{>��7j��L�4�+��V���	P����u�bC���4Z|z�6_�p9�(��l=ؼK"�r|��(�>%r������C�,;uH��o���g�
!�jt���J�0Rg�	XŖB�笀�g+f���R�z:�Eg&�[�q��� ����3��w���\�m�zG�)J"��T�56qVU��2��o}�o���D�8|��<��]�{��ƕ�?�Ib��x�Ú=��,�_	�ѣ�M�.QT���䖇}Ի�?Ǩ��][+�G=VSV�)B���֏ڄ��p�g+�_�J��,!prK�$fN���3Θ��*@4j�f�\ �{���I�����)6:�A�n�g=Ə���{%j�h� �q��n-v��l{"p�-;	�5��Dx���t��y[���M�`z1�KG�D��^W��2ꗳ��X��L����v9�89^X��@��"4�3Bx˺���6ޝwK3���+�����R�,�!ev#�JM�ɡG�pc�\$N_x�{���r��g	 ���.���w�58{�唫Dv��\r������TfA{Y�u"Mة@�T��ބb�#a"��j��a2�
i�\���A��IcR��}��Cd�$�ZsS򛺸4��J���0,sXI�A�4�D�@��iGjq�L�b-N�(�P��Q�WC�J<���`[�̉�$ߘ��F�m�Q�����[�$�x����M��M�(�{�L�9�Spg{ �'g��]����.Lы��id�7W�Um��'8i�%g+-˩J�'�Ŷ(�_����S������/`C-������@�+I�k.����ײ��r[���B+E��������d=/ə�#�.�\5������)�aB݋n��=iE=��
ںAF>�|��d�e�m.J
�D~>�b���g�y�QR��#�;=n2��?�u8�l.
G��U5��4�4|��Z|�]\����[Sa�����nb_�yQ%��ވZ\Ֆ��A��;؍��OHt"_Ṧܰes�3�v�a+�'q�\��z�_��!���!�_3G	�F��.3@l&��㒃gK=���G����ɤa��9ɱ�<�&xm/*z}�z��NL��mꞫjM�IdY� �_�����[ݥǔ-T�n��C�"�.Q�2�Yd�$���4��)��U���*�8�ʰ��J!Ē��&?ږG�!�;�T�O���c��._t����������z��7X3�H��������q�:HO��.���l��6���E��Nǂ���A!�;�ڂ=����X\�4y�f�`$��9��.m�[	�&��G��>�e��է�����q2EA`�����&u��|F�K��K�͹���a�K����m���ȏ��p���]9z��0졠m+[M�>΄�3�����ʿ0�Yh7hL6K��͇��3`}0��B��xm�Z����Ag<������5��gU"�WU	�o(��C/m����j�3W��8ͯ~[	���D
Jo�����N��u���(Ҿ�>
����Ɂ�j�,�ӌ�Kr���2^OZ'N7�|Qyf���t�7>�c�bCvKn9K!�g�s���S<�E|Bf�\���n��m�t0m#���&���אK�d�P/=,�z��)�ҡ.���iW
�s�5J�DF�&��ڼV��ɍ��E%o������k�d���<;��W����ϼ�o2� �R�f-.�i&�lP���Q���n2���PQ��^��s�x����h��͋��~.�	�S<-���|��UT���`����ؗRX�X�t�>Q!��=v.�P�r�d�[,A�&����H��]��j��ŵ>Ϋu0^��B'9V6)q���7�<�Kt=����y���_?��I~�r�Cն��~	�g��P�\�0�6���;  I���h ��ǰV�l�K�P����)�^�F5g��,pG�c�y�bE��:0C���T�YYz;s�m#�\�'t�I`���|�b�i��D �j�\�Z?��gY)WUV]b�6�x�R�~N����PÃ���Bq*,��]�8M0�*Q�"�CQ��z�^���lۆ�"�1��%�R�k�8���N��n
9x�T�.��-ċ3�����l���? Z�L�r	3�맰��F�.�Ai����2��u�������$�A�;��B�̩��k���O��P74�#t�"��Z��b�O/e���RGMkԔ2�Q���s7 �R2�e�����U��I�ʓq���^��_I\ж��>E�����G�&eK�e�����̉v�l�7����P-՞Q �gK�>�R6|����b��F���i��y�aQ۵��6yt��΍����?�Q��\�K�����*��=��t��m�μ�0����+�v�i���5dLdH��Y �&h�ǈ�j��OP@�f�g��X�Ns�){�V#zѧ��C�Z	"oʹ���E��"��x^x\�\�<%���I��in�8��Z/Z8)�KZf8��G倥��S���rT㰜]::����&0�hKS���Y,�Pt �"�}��>������m#������ixTKy�-��@�ǝ09OBe�s��9	�0���=��]$vo�TP��
� ���Z@Ir@�-�
~��0�]?���������O��f�dn�=�B�B}GNl��(�)��P��ןVhk��O��F��>��z,�Kg֐W����>L@?����i*2t�&b�^Ff�|���T*d� x(3���c�)c�(C�Ze[�HϺ�/�|� ��R��.TA%9� ͭ��ek�ݿ�q뭻�z*`3O��>&
M�:\)U�-�)��K�!���O����q�-�p�U�G�{fE��&�y���y��?�bD��������+0��&jM48�1�~4ƒ�=�ʞ�-�Yc��&��7��|L�7��Z���-�m�R��}���3�,��)�S�M�I�0`i�x�B����:���������L,� ��f'��ɨ��?��3\��m�,AVJ5v�+<B��сKCօ��=��^g����.A}��&��&q��ic�"��`Q���K2j���rY�s�#h��~�~�?8���4� IuC`��rh΢��%pM�GGxY��rl�B��C^Z ܤM�0�E]�6�sx[�)}J�2����t/;�*9��L��[P|�O|���'�+���uc�������5)�L����-D��nPn��u���5ՖoB����б�����S�a��<��?@l<�
|��K��J�N���D�p>��"�JDM{�e�E�u���1�ܪpg�/�Z��h���dtM�g��xke��]L��ty��S�8%�C:	��G��cɅo�v~�9�-��,mI�iz���A7}�����z<E
�h0�N+�9\,��K��޹��a�n�}�lb�� V�P"��00�~� vN�����_
��9V:��|H7º'6���1�'4���сER�'?cz�W5l��m�p�0j
gn�^���~�th�4f�.����4��Uv�����|��L�刲�f�)`�WD�˄�^,B���E���H�W3��"Rzbli�J�A�v7�Ǣ��mĝ8#�MBP�u�<ُ�j��}�����N�-�6}��C��J�O���wܖ^��+y�hms�CC�=���h��dq=�'!�Ɣ*��[�r_��e���
��ۚ�I���rc��K���ٚ�$z�b��YY���l�G��!��ĵP ��󻭀��r�<������^�P�6j��FQ ���3p���ZW�6唪[��/s�+��2w�^�Ϛ@	�Õ�/�b�V�?	�bnRi�A�va鳟{���h�cbG����Ps��s��t}sB$�<�ݺIUۃ�6��X�J�����Lw�9z����%�Đ?��������'݂zҀw3i��ɳN�[W����kH` Iz\�^��y[m�Dˤ`��Fpg���f�C �-��A7{���C��VKJ���ͻ�M˥,��Zl��Ŕ�7ͮΒR�dt��kt]�T9,�H��rr�tk+3[��� Aw\B_k�C/Q�3�e1e����t��E2���&*� Z�+c�C�{m�U!iP,/�;TiA�6�(�8��=I&��~d��8��,v�� �z�p@�O4��@�?�uw�^�_l|���S*b�cM>�w/AL�
��/�0�1ċ��
�R��1D�q͌��07Y{�!�.�G�	l!F�U�w�:���*���&_p�)��Tg�I�A\/E 8���[���ѳ`S�\xM�����4+��mD�9$(Q�+���>�%%!#�Y�.w,��2�N?�JB�B�H?�,�T�)��0�+��_�GD O.�>�+	t˾;�b�WIJ@6,v'��o6(�0$orA�l|�>�rK"Bͽ6>�����Dű�h�>nY�WSJZn@�|�1��'��=B�񁢇�/3��чG����IR[�7�;�^_�F8)@���,���K�ޡ!(�yE�p~B��τ0���_�<��|�X�"���1� w��)���2� �d�QE1zcfp�ZTt�~�9��ږۻ�_9,'�����J�`��i��>�=GG�)�=wW���@eέN�Ҫ�N_j.�!2с�����#k���+�,�,b����a�o��O�������\��RF=8�pP)մ���_���Rm=�F���9��F��dC7X�#uD��&��1π��4V�s2<�G(T�^#$>ݞp�r̓On��N�{�:��~9$i8`���"~���O��~c3U�"����F>o���0��F�t'�t}&�Ʌ�t*(gBWFT��vl+)��d\��8�̿��z�y�9T;����/H��VJ)9��j �65lפk��?M�`Ja�J�sܱ�ct4V����5���?TibN#���D�wt�y����OF��d�O�H�,]ޣ�.�\�m���U�(���JO��G'Ȱx+��Z�U}�!Q�5I��.�����jx\��M@��YI놼M��9���47_p5�(f�H޼���iAX�H�~CD�U^_�wH�5���\j^�-��:"��������4Cy��ș�ۺaN=A�r�s?Z��Lϥb|)�v����<潎�y�1ᱥ�5� �/�!�;$��׆n��0bts�̆!�QY�+ݑIx��x����ݯ,�MK�j�p?��'>a��{ܧ�5�A.k�@�Ԁ��W>��A��{HC�|
ӓ�����[I��$)�$'���6�=w���-�>�a�׼�Zo��5H=%,��d��]��L�������A&�#~��p@�,C�Ҡ�_
�o�h1س
���|�#�41π��|>��;��Q�� �FA������"hM�=�åɛ��_f��3��x��L	{���M'���@��]~��!�[��4������s�Ӓ�I^Ȍu)����)�Y�0�w������"�_�6b@�_��!�u��A�!e�W�Q�qj� 2�: jwb���>K��~��Oc���P ����NT�sD(CcY�!a���_%skV�ǻ�2��53��a �,�.~�fy�H�5F���O(�t�"�
I;qZ�c ��U~L�S���ﳤ�څ����%�e����E����plZ'U��� ���**��of�@�� *����@⎾��3u�[{��z�z��k��aJ����BK��%�b��腟-,,ط�qܣ���-B#:joG7'�L�8����mݯL�ܸ���I�"h�� &��#�����I�I5�%�A���}�^�����?�ɖ���
w�'����i�أ��}]_�`L����g�]_�����,�I/{ �_۸gL����6ա��BՄ��}����'@w��`3R
���KG4tT-(��O�:�a�L"�lQZ�����/7Y�r;��^_�	�=�NFH��y��#�6+�>!��
�j�I]��LŏM�sbwN���G�+�zZ�(��_"��j���&܃=��� ���5-[Ve�dl�j��s�[���H">Ġ����|FШUi�5������aXN��Y�r����7���Ce.����o?E�Zl���X/<c��� ��6 -��n<�E���Ǔ >�B�$ؓE"��^���8�9W���-�[�2g��ܜ��X�C�)�i�����4m8T���H�lWG��_ԅ�a��o���[�#G����L#[^��W�d,�DK����q�L~$	-�B�;��.+�8=�=�^���"F.L���,��?����c��Ȋ\u��FX�N��H@-o�^r=ړK�Ţ/6�fln�Q�����P���bK�p�����*�R^�g��D�E?�="���K�i/nl�~�Ƞ�i6��[Kp��+�̟���X�	�O������e�s���x�=��!�t�J Hc�>U�pQU(�D�Ąc4��n���v���i��}R�bD\�C��n�6a� ��.a�9�K�;�3�?�O�����^�����1cAĿ��	8 ��Ҡ�v��)7mQB ��$��̎_`!հ��c�l����T(��M��A����04�l�P��S���k���W����@�N��[1e�T�U!�F��C�_p��_Y��`s�r��LK8��ݹZ8s�& H�v�E��鰧���Ov�[�pW�&� `ᯑ��	ߢ:Z��\�8�4���h.˸Q2��9�P^���==r��P:��DyPqap�V�$�@x=���x_r"x�ŝ�4]?���#���60��vq6�J�saA�"�-'�ҸǓ��SN�&�� �t��e��gҵ	7Z�o���vɵ�hR��J�de�2��s?o��g��+e���F�k�� ��3��u��f ��=�ܒ�Ǽ���G�?����*�ͤ� �5�s���іAV����)���?�k)�mȓ,��� i|I�a����*k��=�ٓ!�Ԁ���c;�qD\k�3�QI^�>o�<�<�9
t6
	
s�%'!��A##潱��"�\q���݊� )���xm�)��|Ӕ����3�k��B�L���;,b�d���4z[w(�B�G��+h�޷Y4�ݹGaS���ߵV�?\�d!���B�����j���6�dMյ���%��Є73�(#XJ�a #U#���=�֯�%�T�ǁ�I���}ǻ�]i<v�	��~��F+�_���4u%��6�̼�4��8���b�1<�@�#`���5��W=E���ԓN���%�1��w�ֻ�sB�&�����g�#e��������R�b�`M8<6�)�.殰,�T�*U�n�(92�!\�J�S#=�{җ[G�g����$��x�<��&x���Jl^e����TH��?�o��żP�y����}?���#%>Q2�<��}�,PR�H|m>NmM�o�(�i�O�5��e�ǅ��ʦO~��4%�](~9_�57��U�|e�̿�E� �B,H: �ǁ<]��9�Ĉ?���b�R{b����މA��G�:	`�+���0���x'���?e��jt�kxq����RMP�G�ʔ�I31����d;��ë�}�Z[p�s�\������b�0m�]�̼���E;�6�0��6�fH1���y�����xs�*�3��������bkY�D��R�MJ�.�6�*2�p���g}�[
���z�� ���/��'U嵨_V��S?
2\�~4��3��D\�5|QV@Y�N�0�M�j�T�l:{��A	f���,J�Jㄎ�#�J
�����	�S�N����v��SGe�l�5�T�VW1��eDIl�<��9��	uX���JM���L[�r����G	��slJY�L�I����n^�����r�����U�#�[�=)�&p)#�\a���������A|�Z-ySz>t/�z���2D����vx�	�:=���`u=�K���YG�~�v�O�*	�rѭ��7�θ�9'�`�X�����Pz6Rv�����f���+�^7����Y���e ���OS�_@��4K~�A׬�t��o���q��,:[�&�C�2�*n��������x���^}����m-�W|l �q
K�JoO��?�e�<t}���Q��y��f��.Us��:��Bn�'+��=Ҹe7�y,bi���H���c���ʌ�\�^>����{�C��ح�Rl�MR� 4y��g)J��lvP���<���#t�*!��.|������� u��|羏c�"�~���)<��w��d	��Ҍ�B��S�n:��wcZ�D4J.��K,ė=����c4�3����߂�y$�����o� ˇ&���k�S"��̔�W����SbJWq���R�K������U�ￔ�#妅^-�j�`G��dm={�3���pn��qe�a���n���+ֹF��4��0j>�M��Nƴ오P�H�"i�Y�N%��"bψ���F$�����f?������;�� 	o蒅~"m�0���W9,p糘mf`֮6�]6��1��Y�O�l���ϢN�����)��R�ˠ4�>%�D��Q`�A�n^�=fh{�j�#x|荶BDT�h�7ڲ�ڥ�a�}c��?�஑��!:*ō�B�'���	~G�����	��n�a��I��a6�}��Y+w�:K*�w�2��-���?��F��,�o��ޑ�0��p<D��)T�j?&���uѶ��*n��N�W�Pe�/!e�x�wE6v�뙪YCP���L���}��'��׿�w3.ר��J6N��R�7�uܰG��א�M���$>P�E�R�e߱���i��$��2p���-�6�λ`����h_��/���B����컻�!�+�?�}�%�bURqϾ#q��*�Ӯ��-�p0J���	i��ԝ�WӋ؎�$�j'�:GUL�P������(�y�
�`!�{��wf�;�T4��9�"��ˬ��F��hu��<�-���rJm���-T�����]�������+5*Q���üPyg_���y��E��%�V2mT7ǿn*� 4��Y�ԺH)~׍b���˱�Ĳ�1N��I��`������T'��-��/'�zr�$�bNa�\g��¹������H{Q���z����<�N�P�����L��,�tBo��x���崬��RY2jQn�DĺX���.*���V�]*	.;Z��c.%�=��J���y��	;�7��2%�>�ċ�3ES7�[�M5��rl*���۱�=����D?��?1d��c���p�����y�2��Ф��|��yD�ܯ=eڼcm��dn�S4ɉ����gLS��rǢ�Ě� �Y��[U��-�R�1j�S@Se��S-9�a���W���S����z�hwL�%��^�>/G�|��FjE�'"���^�xgR'�C�}���F"T.��A��2���%������B�;��T��z�".�Ժf���6��8�Gd��V�(y�Ȍuv��-0!s�������!��`,`O��7Z~�ř�{S&�w0���n�.��TN�=;_�H�^:C�>�~��Ֆ�9�vْo����\��_3l=�Q�s�IY�`��f^m��R��.�A��;����yԘ���"HQb���V�[����w���~��!��K��<=oo�7�Q�A:⩄�����ϸ�(�/MdeA_:���K�����#_h����Sp��x=���B�	�?���B�J��T��l��+m_�}=��V��t��ch�n���: ���j`���~�>�H���E��ՙ�߫����63�L�V)��~2��]��[sU{����I��X15[�*)(���0�`��M�T��l��l��Nݾwk��]C���7�����=8�/ْTMJ��׾ʷ(u ��rM{������ 	tC�]�г���]p��W��.A���.4���j�3��0�Z�TPBI�d�[�:�2n*�����#��v+�]�X(�����z�;�PƄ�M�R�i�	'�c�l�(GwT�����ХձiM*���R@���;)ƒ�M�$7T���Y���l!��dxR���eɳ���:��3��0���Խ���1z5�$��ux�|]�ϊ�/�Y������!�2��8%b�56�?��m����<o�j��A4����n��W2*^G&A��^�����|r�i@��l��|?\����c�WJvZA&��\f>k�ʤ����х�}���Ǐc�ao��t�z�,���IW�{���˪!�b��Q��Ƭu��� ,YHD�/�+Te%�f����w�x��<��2X�xg���JG�׳�U�v?KF��ѺEK�b;��
F}<n�ۖ("-p��ܜTMsW��|m���b�-P�3o�	������
�8��dd��w�q��H��팊� �6yҼlQql 4�f�ڣ��brP�fxǯ�Ȼ�w�8�%k������0����\ѵQ�H2=5���[�����ե�*��<T� �F���n��e7D|]f�&�����;�o�
\�	-Ä;��%��:�8Ml����	4������l��&�p���.'N�@�.y�t�����brlB>�8{O(���� .z�D�U��w��I����s�ÜbP-�k!�Nh�w���32��/ ������#\���!$�h���2M��]��=ef���i6�R�s�7i�bHe�f�r��H��7={K5Q�4ˊ��_2�0����F���W��&8�f;9 ��k��ɤ� �JI�B�#�u9���cS��������@���!�A@���D0��k��V!�1�T$F�p�G���s1�K�B�IvPۊ�\��m ����k�bo�u%�WH�v�Oއom�����:����I9i.�OҟP�O��h������{G��\�B~��1*7��}�
��U��� 卨Z�Gy��#ɰS-]���.�9[�\��R���֫��6��ah[[B�'������W�o̶c���ڣ�v�KLq���H>�0,额b#h�uP	��f}Y�2
���љ�>��Çj����y4`��-�G�&t"7	�	�7|FJ&���H]�u%�̴>RH�\�BDړ�{����)�Up��Q%>�g b6�D�&J�f�K�!�:���9	����N�؃�?�̠�CM�	����;W���g�yD�~a�12��������]�����`"6�}�x��-)���y9��K�R ؝�.b	�rjf���Ŗ����i6�A@cAMW3�q�����=�49?k�j)f.9pԳ�V�"�]C������ņ�y�AWSdy�A��u�,<�J%��;�Y���G��`���ηWƢk����,����U���S?�Q�K��|?�w:=>pQl��� ���K^��uuߑ�����oF����{���V��]ێ�F�3��ũC�Ν^�(�̊�ׇ���@ʋZ�T�O�kӼQn���"wt�>87��>
�ĨX7�������s�ϝs$>�@����R�R��oFu�U$��eM�d'�̱�8kT��c���{4)^����������\�dw�f˯�&�q�GK#`��o���f� ے������v��	;.�y�>��ӷ��� ����y��sk!��z�D�,��V���i:�L���
��\��~q�b۩q<1Uˋ�8Ug�i%��ƈHO���-;eUzC�)��3����{���Ć()�ZX������-q<g��,r��Ϧ�T��I�w�C0XB�e�����2ش��wD��#"[�6���*�0?d�ySX���`�M�}eg	-�dW�\�?�Q��PfG�ƫj��ݞ"�1���jS���;᪳��`K�pQ˔��٢�`�»�:[9�ɬ@��?|��M���aCUߤ���{�. qyi��)F���	"E7JL�)}c'i�Fho�����bv��<��E�	Z5|�{a�q�*a7�t߆9���@�ڱ
���f�nE2�E�-�wxCQ@_L�[6�5W��@�n+js��а����U�Vp�2Y?7�� �f��l�n[�	h��dEe:�]Qᢵ����?��?�Tڛ�i��������8���{�����/*.�m_���+���=ɔk�7}]��Ȼy��:���Dw�HJ'O���;z;?-�D��|3J�.���!<S]���̝A�9Y�l!�~>R�3�����/z�^�0I4�B���P�)�a�)t�g/�MݕWc�z�z��(�����~�YF�4�g�'�x3� G#�Ns��w�2�]��X��uρC>�oU;w�2�U�r�I��l[�;�T�B�~�`z��UڸIb(���0g��y�O�?��N?�8oۚ�]潥�[�(S�t	�Ǧ��SI�`^�6;�<k[�%1s\�]��$p����iĬ����|�>�/Dd`���62��ȶ��6���N~�4��#�m��oW�W����Q�/�/.`w�Z�Lp����E#��>�1s�A-�^ӷ'Ԣ~��=.� ^������̇�Z;z7�3�5�+O�؊����m>W��D������[��ާ�Q���ku�7�1[��B6��&;Q�!.��(x��{��\v�f{�����S�\���:��Sv���c\��B7׽B���1�f눎��	Z����z��]�>���wi�W/ٟ�'N��?��^������Z_�qO�����<]���J��N9M;&Mjb)��Wf����`@��/y�H�կ���N��w�3h�,{��*�i�h���$'ղ�٦��]��ﳕ���i�~T|�n��ǐ]� ���� �S��Y�6� u�f�(t1a�%�\|I��d23�+y]��R�^�ˡ ����i��5�8u�I����Jc�v2}�wt+;���68�~��&4����'�hS?W�J��,�iZ�A$_�z�f:7]�PA��D1�#��쉚U}��|Y]:�
�%.ǘ����\5q��9��KJ�����{�g�*q�i��G��N���M�t�o�3��S������o��I��D�4�g��BZ'�p�0�o�O���E������NtߡB�V8Q�ɞ6&�#��(�@h�H��EC�m�߆�Wd_�@b�C�[�wd���N!"�N>��������w�f3ͱv.\ 4�p�	B�Q�g��qS��C��_��zF�k�d	ǝ\Q�.��%���tg��wK�6��*%�'�Uܫ���m�x$���!�ͪuks��Ԓ�4j�?ю?�K��O� \wM���XVʈ�_�&�>�^8��6K��\7p7[�:������H���^����II��
����kTHܓ��3GD�+[���j^!x0�9G�Gl�{J�_����ç�{=��q��� �ʏ��z�fl@�/2v���T�P;���	����w�6~��N��L�g�F�0ZJ�W?�kdx��,�~����V��bf��3F�"d�ȷr1��|l��k��)R��uD�MF*�#AX��z��c�X	�db��,X�ѱk����Kxi��^���|�a����q��\�@�9������!aG�3	I?����h���A$��d�H[����i�W\I����� ������2j��I�}�d��m^|0���h3�A4�4��$���if�hP^�6d�7���\S+
O9�"����v���EN|va�;�)З焨�."�&#��+c�y�OL���	���+L��Cm(�έ�{�W$�/gn̋�]���='����NF	4��2���ihy ��� ��-�
�p-Po�s?��/�tX�յ���R燝���GS�jV�OO�^p�# ��m�j�Ұy��HOmgg��2c��$�|�(�ځ��˥Jv8[]#��� J�����Ġ��U�bL~P��!��V.�ؘ�U�zA��nB
�r�?��m��H-�U�%z�v�G�=�)��3���y$?U��J���o����:�-�
�M��V��K�?|�`>X]h��L����+5��HoE�y�x��Wliȗ�%7��뭑ze2;s�򊜄1�4�J�������V+�v�����&��I�ѳҷ&K� 2Q��"�Ɂ�S<s�+֊yDƦV�H�P�W8:�E��p^/�=��n�+lʆ͑��v�!����%��E���2�Tg�E�C���]B����@/-����EŰBQ�G�4�Wd��x�k����V����Û_�EK{V�Y�����+�;������pҪk��*�����i���i�^�6 .��&V)�<q+!htA�4'�̙������4.�Y:�R�}���<3@�I�8�2��D&ބ�GKk�-���U�Z2y�Գcg"�E��[U}(��}���^��"��@6�
,̀�,x�2�$����7H��h&�������3����v),y0������e�o�C��U�y�NJD�Ǖ�c�?R��Ju�J�ז�8�{ae\�J����c�X�nA#��2�7�'z,]��ܮ��l�r�K"�j�A�)g�R�
��ퟃ���ԅ��7u,*{���3��-~�W9�����bQf��Q8⭍�W+������I��v��f��3���U�d�����q1ٔ q�����M�ԁ�������y���>��L� 
���$qY{�я*r���TX;���(�����U>&���%ݳ$2��mD`6so��7���m�=,�Ʒ���.��V���&�y��𡱮�zMX��a���0LMzE-\�=�J��?;�x�mz�����k�aX��x�)�b*y(9|��?���{�-�&�x�!F�)q�4�)�b��ͨ�C�!����h+��> �8slOW=��������=WZu�u�37-E\��l����xf:8�I;`��Ӆ�4!����03�?b�ra�b����\�<\��G�J�$qp��Tˋ{f�8������^N
!�g9$0��p�+X��|b�6�?�z��f�(� �1z �M�9i\�1
��!e��GGS��f*����tp�1q�b��=+lJघʨ�C�soE(�qv�D�s��1"ޅ��~�/�H� �47�k���r�vn��1��I�Tp�1�<a8z�e�g��F[_)����rr�%���#K�8�m��4@5c���x��vt>J���d�q��	Lt��0��Qk)PRF� g�ǭ� ��1���%B%B�p��8ꦲ��6]d�6� ��������b�����cW��9�r
ۙr�ø����at�lY1��M�e��m�q����c�kK�o�-%ϳ����\vѹ��[�nX,�oʯ�!!Gؠ��E+U����:R<�
����7[�pҍ�\-��F �0��I�&?�Z�h>�g�sZ؂ڂ%�s�Ʌ,v{�+*�m�V/>m�(o��h`d�uf�0G��2�ĳ���u�I����Ԉ�(����ʡEа�'�<��q��ȗ,q˘�4���l�޳��ģ4�[�̕w�D�ǱS�����рV���tnA��Ͱ�j�z�:?�������o�xE"=�C�WZ��e�p�|��w��~�:��+^��%���Pb�d�d�Ks���L�Emh2m0f���x+�%/ZgϐR'#������G�Z:5�ύ�|���+�}�kRw!DX���«Aܕ���'lѳ| �$ 3XF1���Ȧ�������Qa�� s��b��b]�"h�2GL����ե��D�#������4R�=wp��D�m3pqy68G�	�+�Us��",pU�b�-טic�7�M�>���O�	��mC�����t��Ut������a�?����>2�6�0B)@�^�	���l��Ki�>zٰ'{��CNzކ��3P���L#&t����|�y{���J�rx9�/�s��u����;�2$�W����K�F&��/���W!��<���X펂�� ~�m���_���m�d35�������v=\d8ǓVZ�uA5d���'�s&���h;^��x�G��j󍅅n�%
�3��\�)����O���=*���^j��^p�E��l��_�4B��gS[~���0f�B��{�4k��Eo���^��3H��\vCP�#Ai�uL�g���Z-�^�������+K'�8 *b��hU��ƞΨ;}o�q�hBmHZ�=N�w| �r��\�>kK�� ���3@�ِ�=/����a�L����~o���ny��;x�ʴ}�*���1J���~�nH�`��3����p���6-B
f�+�b��<*/:(z&�b�&�ʿ�&X�OC�9�)&l����VA��y�HA���l�4.<7�g��w�p���.'���@����<?i.�>�쨖S�׈�Yfм������U��+�Ϣ>g�k�>���2F���*\��fu��ߏJm�:�|K(�Bwļ��gFD�l��ĒH�G�7mf8=�Y'RǬ/���2���O�#=��k��e�
���J�/ޣV'�A�6�?����_�C�f�gO"Q�K�!	X��ֻ�`�Y����u遼�RoAe������[�oH�[�ڻgL@?���ϒ8N��x���[��v=�w�y�˲j�G��A "�C�r��	n	`�GZ��G��I��l����yI��}�i+�[B���.��8"�����m(-ㆧYН�Bj�������?�=�|�t%R�5b��E��o\>�j,��Lv{�tP� ys��^�]�c����#�2��ܝ	y7��+X�҄X/dR�,�T0�X�� �8o-`9��{"�+��-�L�u,}��O������zQ�I�o�Q3-����V\�>���'9�:G���R��w��� 5E�
峯g��t����u�1�v����2�q���b)����i��V �?z�7�Q<i2�uDys9�ؚ�IY���b4�}�5�g��u��~Eȹv��h�����j>�3�'9?C��-t$�C�����rŦ��o�"(w�"��3q-7�a�M}�^&b�<ImAa��A��Q�X��_��/t���[Du�k�K'>��C4��.F�cp��0�I�|�������_��"�vD۷���H	�AA�5���=����ۈY6 dbw/&O�8qS�jl[}�3Л�edW���;�&mc�\��'0�������Y�Vw�$��$]�����=�{���������]B�v5OA��jVMPs��3��ͨ���l"���S�����ƹͱ?�M�x�h#���e���4���J��6��Ʈ1�B�io5'��6�J2�H���崵p�&GR�n��KZy�~�^�v��nR��2bYdZ��SAM�멺Јs�d(�&�W�d>^V� ��7&q����3�������@i��F���AM~�b �:�+��R)˯���g��f�B��ITŠ=�Ń�F����ހ���.&�6uQ(nM���n*NTเ�C�"@��:q�]{�*b���gJ�ލ-~x|7�BG+	:��:i��9����hV��
m;?W����[Iz�!M2zz���8#�y�FbV�Gg�9��6�̚�M
�z����S֪��������D���G�ӒȎZ�}m̂����_����	�mNQl觘m��I�Goqj�j'�a�f -1T�kŅsm�ǀ��~q"�k�j�d�a�j��U������
���g	����ZK_p������7y�|���NT콕���+�8�����.�l�Ɔ��|U?�~�h�|��Z0�$:���{�dld�C:�O[�%���f�2Ć�y��YWO�yv�ioq!���:@.�M�TH��w���\�`�񩐝̚h:�x�s0+y��|Z�I�X����Ϳ��o�9QyI �9��Ԑ�x��k�p?
� �QX��Jq��Msp)����a.5����z��jD`����yYS�#�5�G�A&���A
k�Z���Ro��O�<�܌+�2S�u\��k)R5�;a� \�<����
S��D��ݢ��b�xL��ն'/?->��xӐ�璢#w���o���]E�B�D[�1\�<_�k�E�����Sh�Mq���'�[M'?���+-.,�-�/�<:�`L�.�f׍}-U�\	Pdo�Q��-Hdǟ`m��Y�_H�5��7X��[�}�d'?~I���K��z	2ߏɫ��wsz�y��(�
,��c�MlŔ�9H1��x�n�%-S@������W�-���r���/r{�9V���
����0�Vw6^���u���i}���밎��@mQ� �b8:ă���'��X��	�C$�{�͘P酳���ѥ����~�x��q��nH61}�#b�x��Pr����N`�v�@�HC�^g��BT�ك`���d���!�����, *�`�L~ /A�KP?iy�"�h��.���,�a�u��/|�N�-(��dڝ�ScSu���=�}��Z�{�����I�vi���i����&�'���f>���j[[���se�[���
BoQ���m=�A0Z�W6E��V�C�O��0�y$�ͪ,) X�O|��F|d��=%��uʆ�Vk��.���]��X� ;��<��P��m�#�jᢗGڛ�DR��9E8��Z|�m�};q�(�n3o�/���8���&��5��fk�S/��1s�+����BF��L�!44^�yo�bHO_)�,ύ{d(_���dQo&�
�Q:��1�=q�mc��C�]�Z�L���_{�j� �Y
��L��r۞����� �cN�:Ý���d�<ޏѝ �"����0���;����R�s�7�G�$�d��i?�y����%��kP�t̖�T�O���a�MFs�w���5W�'v�RA�-i6�U��3�4��$�<n`���߯��ח'eH^�Ptq	��c�������|����
�g�C���2�94��ɑs7������V.�%��?��F���1N�n�P��A&�{>��^	8��s��g)�$����J_�nq@��۝�61����CI,b��%�( rk=�1N毃�hSƉr��<�R�&>$;x�W��%�e�:�fP%�g���f�s�I]��Aƙh�+�}�D��{�G�@��s�}�r�ca�Q���o@�k�(�<�n󒓲�Q%�t�Q��t�$�Z|�Iz%���e�#�I��:����׍���($&����fV|�߂���E1��\m�x�m%�?X��̬ח;=V�0�="�E��mW�8X����i)w
b�~�)�$Q���g�Īe�M�2g��̲��\W�Fv��������zH��n�Nꝍ��"bõ+Kbl6���������XFD١��8ԋl ��Y�Iɕ�o��1�؜`��9�-C�O���"/�佅�xH\i�>� ��!�B�/-��Ԯ��az��01�� ^ݿ4WT��ƚ�P������b�d�,]~�>����k}x�-�V�W|��/����@�}s1����%�� ��ը�m��A���S��lt|Qe������4���$s��?l�����.�'���L�!
�GJ�J�:���N�3`Xq9y��� #}�j�	V����En:@@���D�V�t��C��KR�5�)��ؽ�xim��vVOF,~��u������i>ΎE�84h���8q_I3����Bk&IE�3$�I���!q�Z]��}��T�a�
z|<�0�6y��7�f<��7?}��Ϸ{
�I�]u�.������	�|k�[�/�:���h���"��|���'�R�����_�"G�&!�h#�W�U��8��<m�Y|������Cw���[����k�T�#�>�I���e�Y�n���>�7��X�0���[�{';8_�.�jM8�pJ(!̟sp8.�M��_��]�D�Je9��吉6���z�A/��a�prKwQ�;�6�`P�(�z`�ה]�(�d�9���S�g�h�J풹��D��rP{��0�u"1�l�貗�t�s��Y��8`��D9����k��KX>~(�N|ZT}/#��k8��i��˧�ʩr}�zg"}��Pc�ݺ�"Ƶt�/�QƆ����$z��'�(����x@� g�c�ДR���-�at���L���:�*��l���WtO4�%�R2wy���Jt�h�V:��M��w�9<V�*'� W>��>ˆ=Cr���`gnR�Gy �#�H��8&&n�X)�}�l_�N�?���`�H��1�U�`��)���暶�^f$����H��ܫ�݉�Q:Uw�������9i�yq�&��m�^�q��{��aĵ���x8T���P�����ʅ���Y�����P��5�����âs�g.=)P���^� .��q���C%�����8[�-���<b�*�hx�5��5�`~A�+Vp�_G&"���r!�M�*R�f�Ed4�N�Uo�G��k�g'O2V�}X��mZ��|����W�Q.��1�5�I�Ң�����w ��S�;{V��U�*#�ĐB5"�M��gzp�[����s%�6��]D������pr�N�dST�k��E�:�=�
���Z�t��r��Ik66+�ҒL����}�%��!����(o���5/��i�t��?'�e�iA�f*�޷�-_�ƴ0�/N�!���ˀ��}J� �6�c���j�q���F_'+�A�I���?�q��4��e��.7�g�H�4�kDT����6��Y�ضX���Ǳ��톃���e��^����h�Q���R)����W�I�|xB��|q�Iz��%N<3���BT�=<����4��qE����f+�G�B
�8���9�+޴eŕ�9��Y�C{8!7^�c�l�J������($���ɻ�G��})�OH��_m](KYIć�5\ic,��v�Ӑ�"��`7<������X!���]���k�QUG*�9}���gIh�p<S&�ݶ^,6�{uEx������'�%�ڰ#&��I���n�f1݆<�N_ ᎘�mO�ֲtr[{�غ0l������V��=��G���3�2 �U��Z�t���n
�5��|��Q�{-L��(��o+]j��<��!6AT��턠�k�{��-<�2FJ���@���ٱ�Ir<�3m�`6�p?�Y�2W/�	V��J���ڨ��k�z�_�;�.�8�
���h��)�յDҧ[�em��n�Q�+��A�k3O2��=��Ѻt��|��.�%@�hu	��^���]��Q@���=���%�5��I"��\"�1ۑ�Co���xQp12&���$9ك�z����p��X������2�Y�.�i}�e�т�>��R�\f�B�ǿòY��AwX�=����F є�rߋ Q����Ύ1�ݖ�=g�����U$
B`m�K�����;�uӁ���� ���ˡS=%�,�%�E�S]u��{��O~=!�D���5����@�مC;Y�J�!� ���{/�l��d��0�F�f���5+��
�^k#�X(W)*u����D\o`��bՁ�������J�|��wXe�I�{��(�p��Kd�Vp��+����1�O��EڽE��Q�@���{���7e�[�te���a�&�h��%'a��G�����`�bi��dz�{��91���ϴ+����ﺎt��������2��A���2+�LHI���Z�(s��Z� h"�!�
�%z�,Jg[WpxV��X��p��eR̵�@Sq�)�S��>�������,�ƅ����Td�L�a�5��(o�^��-�ʋ]������� ���b�c`'R��B�ׇA��0Hpx��ˉ�'����`o���!�{��u��J�*�>�H����UO���dUjƖ�G�	eNW�Q�\��hb�3�|8���KW���P�#U�!��b!{�]�v����x�Q�iM�nV�(�IzV�P���}����Gu��j:r��d~h�P
t����pjT CW�ݜ������'}��n~���G�>738m��~��bj��>=��ӌ�)uV+5�fv��"��-���oqR��T[�.U �������W֮�Dc��lV�E�ֱɆ	'�jz��e&߯�c#)L�	y���q%"t�w�\��elc;d�{I��<h��w��;��-i���p]K�嫨���~��c�[$J^��tW5��zz�R�L_"��Vd73p�迄(���8�t��!iǍ+*�R�I{�@����P��7�*��{������ߒ�m'4n9�V^�x�&�x�� ��B?!�_,��J�ʬq`?\�0������b5�y���1?��K�c�Z-~!{�N�o��]7�'��J����8BR[�LͮK����~Cf�m�j������A���w�H�����"hX3 ٯ|���c��2��Z7�@�ED踎S�ׇ���?���Kۍ�o���6J>-�
���*X&������=������6��@vEc��Ϫfr^X�=^�%oZ�C\N����b���`�tt�x���]_7_���(�Գ�I1Pۄ���ӟ�}�������b��Zmw�a���g�;�q)�߂���
K!VԴ	Ҏ�"^�b�Nr���q� �y��(�J/��%_f����iJh���F��-m�m���k\x7 ��?��>��3�ٴl�ҭy��r7�Q#�muR�&����։eU�9��?�����9-Ό8���Z���6Y`y�f��&���dl�D�BR���mor�����Ѓ�d���������]�W.�Z fU��5�~���i��Q��âsfH��Ku�̎���m_�Y���~��q����D�@Z��B��:���!R#��b�r"�U���|^�sϴr��W�TX�V'�?BMi WU[��,9l����~���|x�0QU�Pd�����ՙU�y"!�2l�eo��V�*W������& �_�KSZp(c�!��x.��7�����O��%i[#Jz$��[iX�81v�L���^�z��
]�����N�yx^3*�O��:P��H��n\��.z�*ǺQ ��� !�J�:���R� ^��l#�s\^y�sޗ�u�����61��) ���D���	l��~nI:��uaP�z�w^�z�8&��A�m�!K}=:3`��W��b��|!C���f�{p���)q�i�'�D�v�����yZ���a�k�kňY/�h`z64��	���d�D�g������M�	Oh��U�K��A����%�5�D�r��ԙ>q%���;+�G���T��{K�>�?8r���?�8:t���)5Ƚ��R�f+�ɉ�����������M�C�#�0E�[�W5ˑu��[=)��x1���������=�!+�yq*���B��x�������������V�h�v^;"#X)�ӽ�Y���@�-D������l����uVW��Z�z���/��s�mA'Ȋ��*�r�c���ی���Q��. ��,��~�@�.����6��֐Б��X�'���ƼthWݽ�q�$Ϸ`�M�NaUE�W���$X��ѭ�D�]p`p|�p��踤�W�����	��z��c��jKΦ�3��j
Rĥ��J`��}G��wo��{�:rs��3-��m����y_"�o88M �%4@��c�ڳ����v<iڰe�9u���	d�vvy^��cǼ��A���j�ޝ�1�³�m�ρ���M�i�o��L��vs�sNM�!�q��f��ɱ[���(~����G���S;���i7�V�͋�5����X�Ȗy���7�(�t���T����q#_����A"t-�7��O��Lܨ���8a�������cɢ��'2����݇7�4�T��Y� JX�b��!�T:���?�M���2�L�C�%_�L�JzJ��:�����b>"��[Jh�<��_C7V���SH��U�
�;ࡊ.��[�|٬U\�*4iF���^
TklhIo�G��_2X��.�߂���*XS{cD�:��K��� <�<�~.J�/�5cђʒ�zAW�\Wz @�s��E=)�����0k���o��L�����%_�9����z�5ɲإx���;E�P�-+�0�����4�E}�}�m� ք��r�eQk�PH$�f. �xp���{\��VīE�$�?�b(G��`Wo�1&���W���L5�?�M�3�<���h2Ne��@l���QRKڅ����v�r��$Z�*i��}�6b�(�l}����a:��!���	�̌���|���D>˙o*�%�`QW�ؽnܠ�!Z��T=�#?n e���h���E�ׅw#^�*:�kL��̻Z���T�ŚgQ#&A�b룁�䔀�C'9;����P����ٱx��L4��?&c�Cy�����|���ˊ(8?k�J �ЯI]\�����.Kr
M��2��EP�E�<�|t�,�=�Ȕ�!u孆D%�x傺V������a!�/�����З��H�9��"˻����-�?��YC-yu��sY�m��1A�;I���#	���_��j�-�efK��k�Q`��-e��%�B���*�#l��U'����L�'dw�)���o�׻�eK��5���.�]�)l�^���4/��Y��6��챈3�?��H����s�~u�!�R�HTW|@W�n��s�0�X�g1����7�uٲ��U���B�)�/\�#�|���&�L��9���	X�Q6I��x����s�i{r�v缶���4�m������`(�促ЗtE)�h"�.9�00�9fҿz;,1�����g=�G�(^���z%˺%+$j�ޥ��]V�;q�A�;�N�meԘ$��~F�K
�??&K�]BM�G���9"�7��ց&��E�]����B���n��z��[ ��(r�?�
)M��Fo_�1+�Ђp�X�_z",��.�Q�y���Ӻ�N��Z�ĹL?#�C���5ɂ�D�$"��n��7�J��4��l�SH��|[ǻ���7;�B9��-�,VJV1k� Z+�y�����)zN�#;}"p}��U�<HF�ꓤ�Q�;�%m��16DP��ml�����l�N�E�����f����,i4;ʤ�����qI�t�9;����^ci򞨃;��<���A9����z��e��f���9�7�BX}�i�J>�	��]*�7������n�WD�*���6=ƀK#V����Irs�����D(��9ey��#�2������=��uYW��M�Qb6h�O�ߐ���g��?��y��vҴ$���S����a��E�Vzy�e��_�����^���{Q�Ek)v��5�5I���$"�+]�y�1鷘� �����k�n��Յ(��$�ux�H�`.OQ�Z�����I��Q�д�vZ������Զ�ꥤ\�?�T�k^�N�R�4�x��vnNy�����;�V�M�x���N[��ɁO����]�}�=�b��1��V-�!�$eSĘ�-��	�wyG��]^KPw'�E�����n]S��� �#,z�F�şi]���0@���J�}����_�B^f�Cʲ=�o}30������(�6x ��3��g�����kh�\sqsq�P�d�hiu���i� X"�?�w���SG@�\Bq-�3�]̜������	7^�mh�I2�L��=o�%���%�;|*�����/n8h�`#;n+�.A׮Ti�&{��� M�̇�f�2;:"�-!�+�d��R�z�5�d�ev�V��|���2����dZw�)���T�`�7g���/Ag�n��B�7N�3��I��`��U�r�Ǧ�3�o�C&�G�>�;������{��H��΂�� ���V��#����t��F��L�k�q����ئfM؇�$�)����(�3�x�(��d��#�}K���yV�9�/�T 8�	�,�05š��h!�:i������?>�b��-�2��������nG��yr2�.���|$�cb߄ԌV�W��R�:HQ�bL�/�إ+!X�a&f4)����6�U�z�_�6yu	C�d��֯+O� �D�.y����qZ	���������/�՗1���x�����۾SF�;�:\�*l ��������c�!��]�@PAUS|V9���l*א]��1UT�X�I�gA����E��Fg�a��:����*Ȕ!6��x�t����A��/o�h���K�L`P�SSZ�IAi��?�j�<����Jy�g/�|����l�בvY�4g�z�arSr�P!�G� C�И��;�W�Gi%�o޺�u/d�0������&�8g�{���=�<���6i,Rį���'�n�wƁ��J�@?"T[�I��Q���0x�[ٝ"��pWq�d
�K� ]~6�̽mg�O��όQ2���װ�eN��'	��2��}��tfl����ل���"�(�ZX�8�{���с'�5��ᣨ�Տj�	ǞiG�*����p֊�[+b��W7~�O�~���s�ű-ZD��&�=�~�n�֚�y"�S����c��W�1#ő�F�_�,Ia�S��k)�&.�C�۾�X�a7�xǂ~�Zu:Su!�g\�}�b��wihk{��JZ� ��7FM�����(��_4����~O:JA�4�}���'�S�>�x�8�F��b:�⾗"�L���F&�m�Z�PŐbо�I� ���
�-;��wt��)������4++J�")hY6�C}���C�ļ�ҽN;�N)K�3e���O��"2��Z��)zj��n�![$�<�� 0��XP���GHW��'�Aaza�DE�mX=��)�t-�2 X�7,,�d��L�߸�N-^�lQ?���Q�
�}����EH��(�5�j�Ļ>A?q��R)�qo&�Ojߢ3�ѡ��������g?zlðΊ��<����Qf4��
Z�=�&��
������@�Y�5��b�]���TQ���Ɠ��rz?���j��6�T+Ir�J�Ƽ"O=��)������!�_*�.�����7/�#��ҧC�ӾN/�4#�{��&R��͝��i�cvs)v�ݡ>\�o/�]�+V�<=ՁR��?�4򬩈c�p��c���2��w����3f�a��\Wiy�XD��>��\���߷8���
^�¸�J-1�@Z�A>u�y�{X�r?Џ;�Y�Cr��Ӊ�b)�0g����?�
 Y3��>����I'gI�=������\����L���jZ�7���B(	*�8$ϴ��F`�+��-����s��l�g����������f��9���rh�8���UZ:(X8�M��Jh��ω�QH�#��G8�5l�r�"������~/��;ԅ�HL�75%�i��T7Z����,�Nv�MC{�*Ҫ���헭|��?�4n`�`[@;X��2��F�g�9�y�	7�^I�p4����Fd����3X�!"(f� �Om��gv��&�������Z��C�&\��]q>�q�p�W�8�> z��j�@��=t-���$$�Lz)a�2��;���i�5�L@�5��EO�0����h2�ivþYٗAec����;���=���.��5��e��E��3FD�H��%ߺ�l�\X0VoL���'�'�1�o)?�
�'y�,>ښ7P���Fq�6��M݃C�w�� 3�1�y���-Svg!?+���l� ކS>ۑ3^�����l�K��^�z�D|����N�?m�9a5SJ�	 $������E�5�2�=��� �4JM���#4�9��3v��&d�b�@?[˞�`[��7��"E�� �Ԟ��ꖡD��hi�l)�N'h�B�3�ܧsd��B\Pt�=��lp�⛑��I*�GA�G�N�l�(H����Й]��
�wIqP*A8����W��X�L�H�NE>6�`���d��ب������A���\����;ÿ p�����O4\}��O&ĳ�3�!]^�ȸ�gf���X�_t<6!�� IRB��}r�mAW5�10��~ۚ�	�D�2i�m�z{r��P2cK9wx؃���9��Od���Z��l����?��2P��4�a:)m�Y��<ڂ԰]DP�*�$
2���9_�&aPIl,{ш����7i\�Hx�T88	��q=IM�ah�C1��c���T�,,���KUQ�Dr��u��iJ��W)�D�)�q�]$�р^P5`�xo�n$g�ydߣb�K`׌Q�@q���y���[�=����t$���,�mH٬j�م:Q�����������
G����r��B��ϳ�R]G5�^��C4�pO�s������zܩ7[���|?�T���,��tQ2���H��K�2@��3`8K���;��O�����1�7��ù�I��:¨(�.b����|���A����ԧ �%�,����� ��L�
�ծ�/�_!��#-�٭�_}�s�ce��9�6��	�[�����v"m"��0�ԝI�;&�P�#�r��y�޲_�O�e��5��4eI��2�V�ON��ė.: d>��3GI%�nD��P7;��jfH)bfW�K�uo�Lwh��Ntӭ�j�vξ|�J�u��4��W����+�W��B�8�{A���$�:}[��;Mkv���M�>�eu_&����伽zň�̆�% �gij7�R=|ڍ��=����h5c?��jc3U��7���V�0#}�{I���-N�^(��I�:�\���M�?H�o����&
눅5�_ā�ʅ��J�8tC���F�<�8^ΤX�$��$������9f������K���Q��֪v	�`V�RvѺ���pN��'����1�,���)?c�.ւK~��GD���?��z@�/ɇbz<��#�6B�µ%H�<�E���oB�硖�@y���P-��.�)� ��?P�"�]:(�K����ɟd>���F��
ð�Ed�O��Z3=�L�ſIT�]d[��o��v�E���|uY��~7����_U�H �Dd(=��V�ZVo���g��#�vF���89�Q=�kR%���ZR$��h�Wф�"n������.2��t�Lʅ��m��Y���|2B)1���e$��=�H7������Jhut��z���=�ݿ���^�^�7�a���F"�i��(n��[����,r�/�f������-�ku��������԰��.��1�$��%+��9[���|�	�C�ۙF��a������?�8�w��Ƈf�~A�g�4kҷ&��A^C�'c���=��;.���6�3g�@&?s��΁�Q*%XYdl��0z˾?}������b�$�bt�r���։�L�.ߓ?�;s��z��]-���5ۊiIu[(�p}IBJ�"���:�L0���W�b��Pj�O1){�E�K����c�1j)D^,Q{$7�2�=��Ԏ!cJc[ړ#�A��^��U�� ��f�W۫��^EU���N��X����R��p`�y�Bd^���5�&<J�D���Oq��!�	��D~A���c�^(�ei(Ka5�j��D,�:V5л����?X�t����8�:��i2�E0�����Ml ���#Z��A�A�0�(�R �1�<O��E6� �VvgV�F���̱)����1(�V-����v2�0�ᅫ;C���6�F�S5�b=��V0u0X�TO���bu/B/��z���@��Ym��\Lx�b�z�3_z�Y��p�nʏ���N��_W���X\׍���­� ?Ȟ�}�&�B^|����x��&���Tʫ}kB
;H1�|'gMF�N�/�����_f2>T�-:)����)'w��a�&�9��>�c+�D(2x�N�.�_�s"k�֛s�5�2��N� �!���藳Q�S	�?��	�i[Wl@ �RF�e�BٞG�_��K�v�ƀ6��`Up���!_t��b��x�6$��n�i�C�ýG��ҁO\���4\Qj��P��B���[}�>C�"L����=&����il>4�+�wh�W�Q�$�B����	.���v�Ƴ����ֲ��h���!d�f�N�b��b�`�p��U� h�E���dDva�K����ڊS�1kj��S�~��[��Mh��Tjh�P��x�ly��?�C*&��j�_��w����|��G+K4&�z�4�mc�����}}���'t�h]ac([]���n��i�71�����hCSt��v�=��KB.E�3�C�)!���6!9Ns�^~'lɐ����*8���ө��ƫ$��������H{�c ��Zp�U���.5�C�P,V�����-�˄��ҕ&��h���� ���c
B,��7�(m�/5��������r�NN�8�b������������\��\30�D6�	���%���P9�Z�Ұ/pSo�x?哳xa�N]�r��\tEb��/��[�v��bV[��Q�}�1��z�
�����f�^L�[�6��T��ed�<��ϩ� ~h�c�G��K�p�X���ι=o<y�&V���%�G�J��di�k��ТN,�JI8d���$�9��.��Hbk��g�vMOm�zsh��I��n-~�����-����dd�lzq��`g��u��
�o�g&����)��9� 0�9$�䳿_�۽Qq����\(��]�MZ4*<��~!j���l L�t�4B#�$������N�r&)���Xސ|� �>� r7�銄�u������~�[�Y*E��fe$2%�gZ�.�U�Fq��|"��$�GZaAI}�Ƅ��v~�B/�P�\���xr�8�o���ر3;@�*�H�Л)]�����t��4������=B=w��F��5����X7hMo2��|3�</�Cj�(�@I�SQu�U��u��]+�@Ě�U�����Ե��I�'N��	�t��ס7\#��ƽ�hs�:V-�{nN#ai^�/�р�=�@�r���٣� �����_!�'*QY�
�{3Y<�#e�oV+���w��m^]Jg��i��i��A.{bIId�)�yi��E��L�z�C^ll����h)1� ][3�귗R.��ho��H���Zj���S��Ie�@eZ�3ė�.��̎+��j��N6K�^	��|��sk
^�����M����+d+���f��AA0<'����OI��9�>x����p�c)� m��%G��T�͜�{uԌg��w1�A��?���K!��K��Ӗ@�5��[s�rW�iL����w �7N��0��}��q�����(�Ζ�dύ<��S�q�[u���pE�z�sJS1.1ny��sժM�<�Gv�|7+�ӵ����<Ak�tL%���~�%G����6��(����d���\U�4�؋�z=B��L��*�C�i��
G�W�=�3�Qh�,D�x���a���s?� y��	��@���|�H���!�%҄����j�,Y)������$�U�����=��#���,?^�fھXr���H���+1�Fm�p�c�+V5�X�!��/�/u�11�8;M���k�p�'��j�3�]�|k������ң��	m��̋�U�O��%ۯt���pa�	́�lb�pl��i��}��!��S�|E
c4��"�Ό���MS�V�<���0Y�7�5�œ�'�2��O[r��̻�[]�G!֧�� f��P�[T�f�2�f�Ox@��e@�'�(4�{����B�P��s'zrJX��z�M'�!^�/N�����)����A1��:g�H���7JF�oF�\,�b9~1t��_ �g:��,��μTi.��S�%̜�C-�,[�T�-n��;��Z�aw�@�Fcg�R�n�d�c�Z-���w�v�-������[��u7T�x}"}���{��~�-�������[��k<�/&��E�/9�w�;��(?u���P\K����i��
j�'qZߊ �j �2r���v�)S��S-���'�SE80�Ғ@FB@�P+}$<�@�lW����M��������L���a��pK��R���/x����#���L<ܢ~�{���K4N��Ӆ=�Mr�F�����WG.�
���b)������JG%�cc��,��B7a1z��a�=Q�hZ��\�fm(�/1�~�/����`�y0���ڝ*͇�"��2X�Ȼ�ݸ�[�]��ҝrX�����1	�J�!ٍa��}:� re*��L!��BH)��՝�����ƶ�Q�S�1��������w�]+E_f�60,�`���B���%]>�<<!��3�5b�9Y���}F�O��K�S�������n��TߎZ~��k)��=hm��8&�V39c�eփ8��wɑ�J�an7�<C��� 1I���T("�㲬�����_1g��3���d"ty�p�؜ ��9��B��9�<+�O��_nk@��C�˞eQ��q) �0��� ;R�N��[RG��©Ⱥ�)@
f2��jA�?7&8��##W
������,H�)�Ea�:x�D@%�H�ud�y|&)�<Feo�s�8�;U�-�����l�4��)^��N
ρ�j�JD"��G�������h��N梜�ڀ�T�����}�\����!�y��u�8-O�����ߩ/j��F���-�\�u���Ƞ�d.X:ЄXz�
H2Pr�;�J�)���T��36Y�a�w�s9Jm16;>�N[ ��w���R�!]�
p���D���b� �*��6H{�H(��h��yǽ��5�UU����^�+����;�)�u�I�a�㻚@v�+y@<Zg��튆J�
<�=���#^.qs�Y|48���t�i2�$HejW�,�Y�����sH�[զD?���ɜ�mP��S�lؙo���K�_�B߅5h�X��z5�7Ö`��u�_�i�	T��~�n��
�]�P������1����`%o=���D�,��h���Ƅc>=�;�z��dQ92\ؚr��b_¨�nj�U4��g�A���>J�p��)�ݵٹ�\��oRl��^� ⸧�aՌ4C�"�����#�'��+dy𯋶���Iz~K�U���7��wU��X�-2�&:,��%b����tD�rA{�tf�*C�v���0��.���sbն��+�q�ޙe|'�e"� M`�(ɇ���0nU�<{,
O�����voMe�����0�m�O$����Ŧ���b����񕑛�s|��"Bߣ�H�xC.apf�z�3*&��yr,�,��zzI.�,=�Iپ>-#Æm�V k��4͑��Yڳ��|9D?w���a����]/���RV1K�FZ�öksSKa9gW��ȷ�C�F;Fcx��Ov�Q��A��P�I�����龺���X ��_���$���ܔ���͚Se��`���D\�')��erqq�����&��_e�S�f�@�<z8#_9Q1Jz1'���u�����r��>�[w��F5I�ZW�0�!��m�qRv+�,�+Θ�s`f�8]FU�)$ƬV��I�K�P�:��D�����{_���> ��<��aZw����p"��Ix"��R*��ܣ�Z����v��g:�0=�L��2,��������x�s\�B4�?�����2v3�U�����v,�+���qe�9�°3�h�|C5'X��|����2��J�'m�q�C��A�<�`��2����nG��f�u~~"b;�p�gUAI4���E/����{���Z�>[�5Vx��S��q/N!�V÷�тy�#��c�E�aFC�V6��'�!��x�2Ie�.|NY������$�Y��Ƿ"�-�� �
���͈ �^AL���X���5Z�D]M*����C�H�3*KG�h]�վ�@i_����*�"��a��I!(L�����~~�8UM����hɌ��4�XF$��������<a�vd���X�ƍ��Ț
*��BB�<X�׈�[���a|�A�|�>�x�?g��P!�R�G[�ȸմ�/!��� *��!r�k�4����=������OV�Ö�'�˖n'4Б��l ��H�M�n;�>QQB���I+	�~�ل��Il�zz<�\�[����ݖ�[�}|Jm�؟�#�2�	������p��*AZ��L�g�_��>��BM5N�u}PK�����ĩp*��h��Ek�����tm:����ԣ�����k1P��sJj)HOά0Rt�ԩh`�q�z&�H®�[!�$Pc6���C&��q�w���[�ȘUN�*v�l�eO��	��V�7��z����,�美fX�c�� !�y�:B��$|?��s��XMT����4\è,8<���Y���Q�[+��[�l4MX)�!T)����)���i��
j3�ɊĹ���G�Z;v��c����o
��]	/�,Gڽu`�����:4T��*{�e�m�A�,Ӌ5�ٸ�.s�`s�S��C�NN���l�+��G17k��6��Q���+k���`N�|��1�N^��Qǖ��2���LO���:=����h�'�F�0���C�����F��1*6��*n�a*\���S��d��Ol��Ы�x�X��+ 
M�S����U�쾣��=�'E)�5z��w��)* ��+�Q+�"�<d�\\3������|y早��eW?��p,'Er����e �ݨ��[�W�f���qG���F��E�2��1f�,�Z���C|�c��:�`b�[5��9ȥ��L�#bLxsI�Q���}j~���Moy(�b�M�Ti�:y�U�˧%� st�U������������;~�֧�5Uz�5�W��~㇜ǋ���E�ԅn��l���\'���/�ه�=#��b�^4����@H�aT'�����
&�d�����C<'�>����L?A3��(��������fa�G�͇�Yb�h#(n�$���ա3�^��l���%�OQ�뗡�Y��v���ja{�|�X�vގ�1���"`, ����!3
�6h���tl"S�Ĉ��%�7��t�����}]���=���$.Ap��~K��/f8�M�T�p�3m1�2�4�yǭ��:Yd��� �%����f�n��:�ͤ�ї�qn�+`G�#
.P&?�� ظtB�H)S$�g�&:�ڟp��`�gqU��2����-p�$C@��2�I��4;�ڤ�׋R(@�OYt��/o���a��)i"58,��[�Z�)��2*}s�k�S����a� \�ebj���e;�}�����E}(^��y.}
�b75���O��r\W��W)��Z�܇Y�\B��s�����@/�$���I2�����3g��}e�|[m� Bؙ4�T�k��n�T�R(���z��9T���,��[>�mmu}��ߍT��Eh��W]97� ߬f�{�J˹���z���'_T������Z��vLuF��8��;zldA���P�J��6#G�Sj���M?@o,ge��zi�{Ǒ���5��������n?�q��x��Ҳw4Q!X�X�Ε�nD5R4�/}�O������|/j�]��SS�z�-�L��.|s\��Ɲ'�W7��?��f��l�esg�<ZSЂ��*�,�*� �>1�6a[�2�2�A���b�Q[Ʊ��̓�<mE�:@�h��r��kpQXi�c�3��T��{� i}�nV!bo�DZ�QK�Y����g�6gpw�1�孀���"w�N_�6RH��3hp�� �HɄ
|�"�󵽟����M�����T���P:ʣ����7� {��b��0l�����!S��#�[���g�m�z5�ӛp�/�]���<��[#�P�4qp�+��
]-��D�g��_fn�i�^���}V ��[`�����N��+	����s�XŶ���+{(<�]�T~S0�Y��a����N���܃cn@�G	�>�?Y	.����ZOC�h+����Ͽ~�F�ț`S� �7�:�(����]��<6��&�;�cG��e �a#%�E(@�zsû#�# J&�I~�&��[��8���Ь%W,s}�!u��o'@I�y[y�;HN@`�3���6N�5�p;��z�R��m�Dx٨�}bB��[[g�C""^n�A�P�-'7�c��~+��kHnX���1��q��"_�W�I�Z��>�U�:�c�㢦Eb� \����@�U�L��UWX�&�z{��G��v?� ��A5412�ב
l���F�Ծ@+���\�p ��>�*���4
��0%5�+u��4�a�?��ܪ�����l �	�5h�B~y%_T����UFK��U�E�)���,�Z�9����ז�uȺI4��^B�L�k7��-|���*��6����e�e(���U���eКz |0�2��q���f��K?�-Â���DzU�����0����'��Q���p�b��ާb�����t�v�kR�����u`�/>p�_+�:<Rf�m�򫍮%|��ō=�i����>�<F����P=
�oqTڡR�Ʒ�J5==H5�z�\븂D=�WN�BX� `NB�đ�"#`%��o�tg�&�~�S�2W��z�JH6�"	�?ee�}�qq���w�bJ៰����d���f�1�3pйl�g��O9B �=>�ݗ�T����\3��9�0�<81���
6�a�����G�����Z���66�N$�
��	+v�da��[K4�[R����im p�
���{��esv��n���nrN�U������,�����U��B��v� eQ�N�����v��?r����QL���~W�N�p�	��9}�2+�:i����o��F%����Vʫ��ar	ĺ�r={��_�.ʢ{l+�*P=��Ǝv�6p�m�/����,&��ꁄ(۬n��t�xGx��i�����3��|���1�#8�pZ��X�35�3#���8��,�(4���3!dT�C�R3𦮛���}�QQJC>��Ar����j)I���o��'�����pOpÀ>u�zRK�>9�^�r"[e�y�K��%9��x�i�n��cA�e�Bn74!Q��k�h�د.�$9=e���e��%l��/�M�$g�7d]fB���37������֡��Ҳl�n�b=s����`��s
'�d�Wv$�� �REi
B�. i`>O���͞���[�x��!V�d��&}-�ۤ�#��s��M�x�W�p�}O���d����*䰭���41�}��o���J&6�����V��8_��#[�������]��g2�=�~j�߄!�4�����ޒ�pBc��l���K
�c)�!}m�݉��6C�{ŤF�����y���wtrdD��.��@|���?���@�6֛u����	�g���C�6D����y�=��Mq���|nuQ��C<��o��i8AE�l#bk�[�0�j	E&�v�9�S"Pq�`�G�>eF�y~�E�̹��z$�Z�}c�~YC>���P@���*gXc����ϔ���a�(&��*�� ���袷 ��f������n��hD7E5Y�V�����3_�*xO�&�T�#T�^��8*V��5^C.sF�<�y4B8�䔶�Hh�s�PRu��%���	P�)�ж�R��Ԡ�`�-���-J��ֽ7��t��8U�����[3$S��l�y\�-�'�ɗ5��QH�ѓ�5�4��LܺP[��F�J&�����(=�ZXІ^�K>��ӄ&��؏l�����F���^|&3j�ټ#}F�QY�__���û��lv�h19!����S"%����z����n���)L�e���*~hY�1N
�e�̮]�NȽ�`A�]��)��SJpG��F����i�z��3��׺_�#�MO	��?�z��u~1��-�HwE���.,�]��+��!CD7�-W�)z)^3:\����R�l��$H�c%>c=ܺ�o��;K-��s�ƚ�"2����P;��&�7Rp�Q1\��m�=�L�p���|�h������#V�ۡ��J��ܘS�Aݩ���$��(�eZ�ޝ��oΥ;���:�>�c��������C�ݕ��I��Y�H�²pC�pP,�+�O�r�BM��l7�P�VdR2�Z`6G����g`2ء@�۫�M��-�l��$�3��i,���Ĺ1�����~�No�6��~[���ǩK���I,V���e٫��bb���az��0�}��76��WQDn�s";d�+���OC�21M�>7��"�Z� ����r�}��EF�Y*L ;� ���=���<F@ہ��x���2q��wt�MkRL�2�+/6�o��c��8��X�����z�۰>��-b%y	$>��nQth�6���5R�zu�>� ���)�� �<��A����8�B]���,���B��+�?�]��ȱ��i�Z�hB��MR/��B����J��]���q>�k/ `_�T�9#?���k���c):��s�E6m�^�oO�#��N���$z��x��-����ϭ8� H
uf<p�WICLv�Զ��7c89�#�� �mheY.1KG���x+�1�8����X�R@�/��@��3������Q�ov9����W$Ƭ�爙�yucMb��t� �]!�Q�n�􏏫��a�����|����SQ���(�˵���׍� <�^�e��~�K�I�֌j''9+c�����/�h����\����᷸����,�2�j����I�ʭQ3��6����9�i�F��]��B���V��W�I�7�IggX1��Q�xq��@�3�U*[��R���}��f���l��XU��W-1'��37��A{�S{�̫��>��p�H�(�QY���)���"�����5�Y�>"�?&}����"$��Ǹk� � ���OX�����k$Hș�Λ&�ʼW�>�菜#�s�F&V�6� �JC�4���8z��00"�;��?䳵p�J��+�7`������>*�?H�� P�km�c��������B9v��i�lIr0�����%����F1�y�V�ޘ0�r��@bǥx���?Y	c1��.#ku�� �x����YcZ����u��bòM}�?�� �.0HbX܎�c�R�I͡y�	r�s�#}�g[|#� �nM�j��xNH�X�7�@ᖃ	x��Z��O�@�8�^�C��[Ĝ0+j�//ҩ��5��+�=U%b�C\,}�)ky=�BNgx#��F}�;������t��&����VB�e�������Ï�3����Q	��=,�DUh-F����L��5!�)Q���hg�"�	p��,BB_�����q��(�����+��S�7x8�PQ7A�Iz�j��0jH #7�ۍc�D"B o���БF���g�C�N����4K�8�CQ��}0�cvW���
�?<��W���'!��Í����z�s��pq�^�+"��
���-�� ��6(��݅���M�'� �c��t��hh%Hta�le���of���ܗ��k�������1�,����Z�).!��J/�EЧGjؾƆF�|ٙ�*7B�ڽQ�")��䬸��9P�|A��ӌ���p�~�c�z}I^���60����#���$�f�N��ט�u��$gi���hd��O	ֺ)��#�Y�,#��΁��Ҵ1V+6:��e����ِ���ٌ����4v(�'��υ{Gj|Q�d�̺U�C�w]�ԝ(m:a�W��
��y����ʬl�I�yu��]`�۫ ���\X�]zT�9N8_4p���4�ע�E����G_"V�S�M*	ҡk�����yUl��6P����C���g�����g<=X%���X��k�g�jb�;>��m������ݶZme�ޣ0Ly���%�p�X���ز�S�����򦬜���R�p��q%Ԋ_T�r��	n�w�=�mM-s�ԔN1�O[7kP�5ҩ�*s�^5��V�c~��:T��� �^ ��q6i�$��?�dЎ%R�"��7^Bxc �s���2z2!�$8.�(���^�R
��d�=�<*Uy��d�|_���?��_J�jgl�q7�NZV�&Ѕ����X��	O�!��Q��G㥬%�]~�r_-f���AOR�7ݥg���Y�q�� YT�H�4� �5J�;f�>��?9�����l�ה�!h�(����9�'�j|TQ0�o.G���J�d�v}�T'=cg�u-� Yj��n�ݴ�LМ�
�M���0Q���蠞t�x�F�?8�&]�y > �E�1 �(l��*5{��z�3+Ս!��K�
�������Q�]3(Zw�N��Mx窈�-��f;J%6&�$��0����q,U�ʕ%��)B�N�׍M`����bƗ)fſ8��${�W�q�Δ�7ܻ�ݚ�/��_�����$l��Ix>fN^z��1�!��K��N�2ǹv���%��4u3��x�RH��:�?y�\���D��n��%/��,.�F�x��9*���g�Β�+G��GQ:/=��=l^xlW�#`��:��)ҵ��q��ĭQ	���A�DW4������#��J��x��K� ɘ|#h�d����z�|�k�u������Y*೔�����ާ"�YԀx}�@rsܟ^?yrP7DWJ��3�58��<��H�w��[d���!}3�.3)�.vNφV1h��p,�jvK]XNխOdW1��$����~5U:U�2=��vţ�����	�zIH�p�q�.�~�K	�Z/�b<]%�D����]�0���[jdL,k�/1��Bǒ��v?��d�h��_��h��
9�E��aL��x�D'R6��4Ib.����M��}�j&�����L �*уd��iV����1�ī�5|N�� mc5�����V��D�*��K�����N���q�^�7��H���PHO>s [�Q�8̝]ya ����,�z�8̐yJ����i`�;ōʞ@��}�Wu�()�uX_"����ם�A[�A �nD����0�
c���Sͬe��/�GL�\��
�����4�>�6�Z
n�A�X1'��KE���Kz2����z�2b�`㰁�9��Ŕg���L?����2�P�D5��[4)�OH���GontUٓ���'^[��4'9Ť k��Ƒv@<e��$���9��u� ��P�Ԕ���4�W�Gգm����v�%�/�V
��vƘ<Tȑ���x��Rb�{�1 a�\��e�E_�[B��R��_���������kQzL������]j�������p���)_³Q�"�[�fL��r��Ǩ �#�n1�㣣���V�ʄ�� �V'y��b0�c`���Ot6l�o.}Ϭ�&0,)%��L ��Ң��$�E$��ܒB
�É�+��]�0�E��sc] B�����l�B��Ԓ#�H��u�p���Buw��|�uR�orz�/Z��
J2;����rFtPK`P5���EcY �݅e�08���2N+'�:�<Ơ_6�\��X��8/��v�����0J3�׹�CY5�H"�z�M����bȧx��L�*�_�����جA:�ҩ3�O�@�,TM�Be�^��Ϙ� �д� V��^Xm�ظ�7�]��Pg��<��Ղ�cqE�H�o}��̠������_Զ-���d ��Q��8�<U GK4&���5O���P��"d�E0�<�읕���J�l0�K�Ĺ���v�K�YF��z�P��^�8�jfw!���Fd�6��.����g(�lo�!�	�d��#U��p��yP��Q��F����)��**XZA��*�������O�{���e��oV4i�^��ra��mq0; ޮ׻]&�df�s�W�#PZxa�>,�v˒Z���"eń�~��f����A:s�a�NJ �m>}3��Ў��������8{�aJE�l|0B~_J��8V�O(=_%�VLG��%;���:&b�=�WpPk���ԥb8�P���<P#� ��_AeY���^>,&�.�Ԝ�*ã �܊KS<hR(�H�gC*���ƹjហs�Db�������|3�0 �ꮦ�U}�Lg.%`X��r��5}��r�d3)�I
�Z�����s�i��J[��R%dRc1P����E����ؒW�@�e	�g�A���VI�9�4�l��/�H�F�B:%ϓ���=�@��4�#����F;"�S���̈́��=��*S��p������k+1���| N9���PȾ��ȐK��fiu����>l�Lu�b�Z6s�D�����6�S���ۀ>;ηj�<���vH��/ٞ,�{�a����U��<��
������׏$����0�1DI�(�ӑ5I�ŀ�
�`H(޲p�Q�m!��b5�$ ���b�tPjupؗ�U����2��pu�}lL�j�Ha~M�8Y��F��N1�B@-kRì�t�0(���QK*No�Bh=�R'��U%� ���`� �濺z�.^��>Ԯ)�d쵒�u�OZ�e X������"ဋ�H,R�"B[J��U��.���� 4{7�QC�/k��v[�֬U��/O�4Z��B!�Ct��MY�N9�y�J��;�������%Mq�_E2����z�m<U�[��� �n�W�c���~[[G�M�u���O�h�
�:��O�����#���.y���	�g.�$-s������+�g�{�����ca���}�@Xs:k(�ᖼ�)u2�DL
G0��Cv֍�e3���b������y=�X�ط�䥶�Ğ$>(Z���q����6K�Z)�E�^��l����>i8{���=�$3'�fg��RFx���W���&�N�D�W�y�&<�?������C�զŕ���ժC�7��gcd���@c�Hc@������yW���2)28S߹�EdZ7H�Et��{QZ������ښ~��Z����摪M����9?r��A�� k�娌U
d�L~U�e�6��g]�%���k乵�gM4��2��'N0�#Nt�o�T=B�^�f���\hI����1�f���;�H���'�ҹ�AC����u���E�l=#�%j�Q���,;s6('n&��;����-��q=ѡo��t	���	|eqH5�/L��j�D�����;1y�*���WW��@���BR�d�C�	�,O���N�@�P�����A�=�g:�=�n�&,g�q�W9~�	Oj�n��:�[h�P<ҙ�g�>B�Y:�Z�m�;�K����dMZFNZ�̖�U�}���y*`H���R;��,���D�������H�0�E���i�PxO<��,AE�qe�4�D�w���ʡ�U_��I?�-��W�ҿB+o�E� ~{r��i`����X�M�R �����ț2�T�q\ǲNPΪ�k89�Č½��#Ɣ;�>�}:����Cr�����j*�ha_89���[�"�Ao���wR�nk�	F�g�b*B�E�0�i�W��ʠ}�Y��#��{gLG��ɡ�շ�>�>/�@ t�m�,���v�D�-��~5�e�1�b��f�{����u���y<(bp�����+��e�1����/	ݻ�����DS������н���;X�r�4��0&�p�ډ̥7��G����	�˞Hk��
���A$#۱���}%�{��>�/-���ɜ�Y)&�o���H�OmK���Ï"ꍇ4�����t����O&w>��F菠�xI�!`D?Q'�|��8��!�
 8�E&l����EB-pwL{3+������v��Y�sxZ:�{��`��.��T����R+t%��"���
��sK³�B��R�H�*�-�c���:kTB(�ڏioN�yoC2b�1+/�)��*�Mn���%e����E;!��~��,}�`A�pXy2��M�TDd���:���w�Ư0�,����=��Z��fuup�H�!B�n�ڼ�oϕo���9 ���R=�8��847[@%Yd`�pB��:Z�"&��:P�[oy{k���S`�-a1��R�c��;C�qh��M��Ӎ�SLS��V(��~uY��O���(�Wg���"\y!FR[��1�����ڱ�#N�P�g.��
ī7��hϰq�e�r�8�:���)�_
�Ȋ��W��;��=vW�!�gz�������^�% zFut/�u	o4Zmf�I�L����K@ђ*��4�����.ݠ��`�!ҕ�w��TI�,����Rt�K�N�\JcB�zܯWb&�|ڌ9��n�tXy��`s�BE��I�1pJڳ���������P� �Q��!El�Ǫ��n�R�j|�κZ],���ڶSB^L�y�@�0�%k��!��L!��i������z�"pNy����)���}ڌ �%���jL�_;d��]j�ˉ�S6�t���(}=&x�~�&�2���dÂvW-��g^������M>Y,�?��Шq��!��í�!cA%���ߚ.�+(	"ű�opL	DL[���oFcES&�yq}ʧ�L�#%�^sv}���y�K��;��wc���ѾeO�.���˥T(@�� �N�F�Y4�Ń�F����b�V*g������䯛n���R���W0g�\��-!�k�I24��NC^�o�uG�e�d���sn���~�����a�]�)�Vf�f�m�w^Gz<�����͘(��`\��	A2�M�WB�N����ѥbq3���T��O?������a[�������҇�Q_��c2� ��������$#3t�B�왭�kuQ�k@�o��n���T���I�=�p_�D���̚�0���Y����3�?�����U5�Yo_�4�&Ҥ�mS�W����8���
�Lfi�)�2������]���vIΛ��z�L䁤]]kR~kM�v1=�q�W�GX%?q�:8�-���8�zv�\og�-c��%��XT�	����ci�)��}�,�?d\k��Kq�����תː�_q��@u[+��~|5W5�\&�ɑ��o�l7#)%M���hߪ���R(�_~˴6Ȟmxe��mBt9m�2F�E|�()��\��5�`�v�[�[��4��*��n�⧵�Mr����.����+��+�p��oM�n��D.Q4u�x'B�
B�֛�%�S<f�A��@�[�.����m$#5�Ec�ur�^}�T�7BfA�CCf���_�M0C�T�V�I��I���"� �^@
>�Z��V�����6�e?n������Q�m\t ������͜� Ң�__K�Q���@�`3RxJ2��ĺ��Um*n+�]��IU�v��}�r����%d|G^�C}�"
c~ �_�'�h����P?��Uw��:H�� v9\�<.�8����5�j�2\I+Xu(�i�VNՖR���b���Oo��5sX�"��) Y��4WBt���o��.-�5C6��?V�~��G�gr�'��\-_v�`?�]5����S��r,���x��,aڐe]j����j�C�?xw��iK"�\�}��N�/�e�	ϋ߬�U�J�m��D�����,jV�4���/�F>s���E�R�vb9L���[�#��'5L�l�X3g�K�nr:���<�(_�PwWga�1^P�� ��)4/i!ש$���4Y� |�vn5�h�฼�uh2��*�當�C�=Y�����*AU1�أ[�7fE��Q?�1P~�
��x�A�{����DPD� t-đ�HE�q�L��4P�-��C�Y�KqL�8�|U0:�@!u36�z8����`����_7��t~��"���ѿ�*�3HR����5<�aLh�t�O����<��0�z��TD�1��<j31�Hb���������l�}��٩�����X��,��v��8�Д��qR
��Meݦ��Ti��ܒ�-2��$����a �Q�dBU�.�l#fG^���oZi�.: �=�2"�.�vϬ���o���ƊIv�(ճ�?]�v��a���Z��n��d��b�f�5�uhgA������v�7R1N��0>�Ј��ѽ^��]1���mWsA��:���Y��'u�|�����?-��\ɿ' jZ���ې�*&�W�Y��c���nծ�x�i����'V2�J��?5�:�=Ʊ�]C�B!�@���3�y.#%��͋|2=�i��_Z� Z>���D^d�Ð"��~���J��Y���w�}]M���4MX�S�%XL�����>;$�:���菍^4��ye���FZiý�&�FΟ͛؅DS�D�S��}Lۉ�� R����;!HZ��o\��?��ǧ����PVE�x����� �
0�S�*�D�
/��'�e(U��&H�/B��?�ov1-����RX�m��gAbE~sO�dZt0���:��S���PC{aE��\;�VڨY��GU-(�Y;���"�'#��� ��[�wW>�7�e�3p�� 2j3�A*b���d��D�����[��'�Ʃ��g��9�2�.6C׃��O@�1�M��5���
�GR�eQp9a"d-�n������l%|P:n��q���z�q�4��|�|���}K�$]�MfvX?��4�_�k˅d�b?��Z"[e���u��k}�J��f@C�,M�n�]ey~�5��7zK�i#���P\j�+��q�����,L�"�d\�y�B# 7��9+B�u슣5~��ha^'H��[+]�I�����P	yRI�8u
Or�C:1UB����/�u�e~|���2Sª�s���i�z��3��Q^L^�t/qQ����OWH�R�����������coU�����#1O�Zye�<lb܀�j����4fH��ui��k=��������A�nF��94=6�Q�����L����#huDc��7�[M�_�&y�W�
�����[��+Z>�ţ��
��HF�7���3��/79"|�W2a�'�IF�M,����7�R΅��,�[�)�\���.�`�u"3�
����Ak;��C6}�/E�;�5��_�@��W�_�ֲ�k���廴R���]�����V�ݪ���TQW�T^��P�Eܧ�%��z?�����t��M��&%�':��*1la_x䤏�fb��Mr?�(��K������M����K�q�JX��DSs,�h����I��̢��ի�+l5�a�-�Z���#4,�,~�����|jU�����a,���ǀ���ｄ�ԫ*��m(5��V��� �D'-d�B�=�:o-��?3j���BH"1����+���0/e��u���b��dy�X鑕�<��/H��&ۚ}�߾.����D"M�=K⧆�g��-���'J�6�nD׼ܟѝ�4�y�.�T��E����6o�g;�jGt�� ���1E+�^��/G��T8��ޔ,ߴ��}�,��)�,gC�ŕ�`I�Ϭ��������e,�O�t�����eB�i4�U�Sw�K� ���Ǻw�����׷MI3�4�{Rc�3hbi|��ӗ�#?+U+@	h�_F��`���,�;��4	�+�����e1�#�Y.O�0``\8��ogN�bq:[♇Wo�J������%?/�v�9,���/O �'򀛟[Y�J�*[��$`MP�~	w���\�^r^΋���^�r��v}��>����p4o��?6C�	�N���'��b���f��"&�{�4���y)�N�HޱO�h�#��q��k��p����T���
�챋��	�@�%����d��Ƥ��S�^����EFG-�s�^�QI�g�R���Ǻ��)A�(��`�@j�s�M֡���%�NV���)&��{5h�r��&�?�Y-,�)ɟja�Ӵ�~&���2V��I���B�����`�g?1���~BO^~�Fp���L�A�N�K�4G�&$1��rt��,a�g�έ�J�h��=P���0���FKo��_1�J��(�Y�� �h�6�����D���$�>ܵj���j��1���y,5�t�sמr�d�<��K��3��Qm��󭂛��3�/Q2\��\U~��k�>_T3��t�1���Tj�O`Y٭|�!��#4���}���-p
݁�ٝAZ��{���[j�g�
��Ħ�H����qKl����V��#��?	����� 䵣�5�֕��W��܅X*A�1��hC�D�l>���=@�COW�o!h��r��]*j�I�+^m��?�,v?�֩�Ϟ��=p���k��
���lS���d�MUP(~Oۯ{�U־�SP���*��%U6MHn��ڽ¬D� уI�X��R���{�b$�(w<�:nܡf�?Gt�A{=���O�I�8�]�M�]�D�p(����nm��4�ν����}tol]�*�������>�k��=[���[�Dp[�E{8d��y1��W]k�� ��d�$����fT5.�x-?�����_-Z%��c�\����!�	r�q�Cّ�ֈ�рŲ��5��ڦ2b�|�'=f�0GWB�$�!��Y���D����s��w��º.�x�b��� Y�i,{L�����l��`�e��;�D�`M�s仼��'[�Q���-"�9l��'3�c���X>|��Y��6������	�Տ��o��B�N����B���
U�s(�RO�q�8�U����n�wy��tї^$��=F�+��#("�gL��w0N5,Bqe�[A�7�=Kf���ezc#�I��[��
J��9ϱ�Aϻ�G�$�o%�p8��z��L<<�(�4��q{�5�J�c{l�~�����k
�v��"d�rx��� ���)�~�����j!ɺN�*��~�C�x��N�Sa�ѩ������`�b�M��%�ܤ�7Rm�� ��[�|u`�����t���1����?�\i��	nc|�`v�6�2�[�
�����Oc:�ޤ�I�e���o�#�eM���C����<6Wkk��������9$>:�&O3���ߤYhI�T]�-�J���B���c!	z�#T��@�Ь@@�S�RQ~�M3����?u�n�Х�%<X�KH&!�`�_���f,:NT>�]��60��ːӂ��<9}�f���|[]g�.�֬��fJ��������K1��1oE�E��h�W�De}e��Oi쵝a�����Jp_r�������:��DMz��ȧ �Mi{�u�r~z)&�����UЪ+���Xw2h��);���B�U���:*��̺�ңsKRA2`�&	ݪW��~�C�݂�(�%@;Ov��2�Q�f	|R���D\�(�����v�y�>|n]������ҩ��i��:?�&���u���rK֪��\5�7a?N��R����xD)欒��Q��EEd�qL�87h� �{��;R�к��^���o���3��;�\�$+�Vc�P}���ۣ���ރ�@�C�.;��8�DO�!�_b�R����==����ƺ�YG��PO�ޏC�p�)��.Q�gl�����R��L4R�.i�"��@	�8v��wÏS���c2=�QU��
IM�X7I���+iV��*bc"LZ�و�������\hraOr ��EF���;�9����Ԥ�St:؄�}��H����
D7�fȆ81��O���S�:��C��ZŮ���ͦK��#4[nW�T��'\��_	�3-�Ҕ���d>�^����h�M���N�5���~�8�%�ڱ,��l
���0�����^�9��fm4tso)z.j�@����M
�գG"/���@agMm��`P�sL��4� p�v��;@+䥄�"�k2�k��,	��Z�>愹��w}N�s�0��V7����)�n��{4�~<�'x3ܗ�>���QVe��*�5Zj%$w��Nzju5��՞�I�G٨�J�-PݖmM��׎�7�=���W*�jz
�#�fb���+��b�Oh[k�«�F��h �^��D��Sk5�y��R�	ҿiHe_��� e@��wYY��x���[�3���C%Y���蜺*0C�<���g�\�@V�x��W�wgd�O�{���ԋ�S�u���#���%�����@ؙ��p+��(��اňv�@l3�
��K��C�O�9��l�Y0`<h"��0/�SJ,	�#a�%�Ǝ�����Ѩ+��?�����Tހp��i:�9Yبv���B��(��`��A �+�\����D>�Ee5%�@�Q��Ϲ����-���}�s�]|98y�=d�#�u����$�R���7��7���!uqk{2��@�_E/HA^|OEѱ^9�B.��,�mϭ=���أ�T����v���U�(��ZHV3K"vrQ�<��G�DT��a$9���|-�yxk�UL���O��Co�|�l>������/]_��@ΛԮ������W�U�{��y��ݯ�OtK�%K6F�c�}W@�@���"ۛ��]��t�w��ޢ7����}=,�H�j�፥���%���T�q��#���0/c�(U)��b�~y�:���(ܟ�ګo�9+f���}9�/C��yފnI��̦:��ΐ\�31,���0���y��f���|�i��jI�Xu+]�!��}����t$��3���;J[G�{Ul��Fce�ld�������~e���%0��e���8���=����Z�`���2����1�}*Dh��*4�#ۍF�̦Z��F�ln�ՉWc%A�䣄y�٩�0�x��%į���H&�z�}L�����b��ƹQn�J�Ҩ!�G�l�6�����)pҎl�e��~�e�su�v��6&ە|7�/Ԩe̴����v ��d(�%�褍�\W�l�|�&�W�1�^���L'75�v3�3��ш��w�������I����� ���3&��o�>��
	z2�E�������W��&s�2�8"��I9d�i1Y��؜�����$��>h,�	���v���>~B6���_��ɒ2������f���.�e+�f[�R�/� Q��T���~x�qI��;�~ �"����mcn[��\�w�NH�]$+yq�..(���U��Du�wb��_L[W��\��A�3�]����we�y�|��$��l��)�����]g�a�yۥ�2/n��vYn�u�� �h(t����럺������-��F4\�Ǿ���'1�@��z�W���3�IR�='}ܢ<�i5��ԧ�(d��`x�$-C>\��]���:�-��hr�Ӟ�3�w��I��U����&qZ��Z��n6'F��:Q]Փ��|ni	\22X���xݤ~��G��m��?3h|;���H=�!Z�|�/��>M�^x��F'��7&GP�;�(����e�*ɒ9��$:V%�_�,�Һ0?8v�t���U��j�����Tb6}��;�G�o�8;^Lh��S�j"��5,�1�A^��J������Z��-V/����gq*�74&��A�A��oj���X�r�C�
��m�6���Ȋ�SD�\B3����y( N	bJ���8ͯ�D 1K���h�p�/'W�9�~���R�цᲮ�/5�� ��� ��%��-�p��:O{��'p�@�)
�mUR£y0��5�þY��=�Z$����D�p�žZ���e[,U�vt	�'�J�&��������D͍���Ps>S<[)�))�#�=*��}�S~ 7�Ը��3�nO�����位���;���ev���B$g�$@}����_1�1���t�����\JD���"�cOO��=��
P �Y�ظ.��z�:��Z��bĉb\[2%�����% :�Mȿ�mP���҉�w�w��P4F����\���@[�c_��N ���ګ �[P���\���FR {n���i�VF407J�C)Ir]4���e��M�l?�'�F؊>���*�<">�td���1�;f��	]�G'Y�oq�.,��em�@�z�K����*���+*j�m[��FZ�xA���@��t����b�k���㟽_B��[��č�k�[�$13sTq��dԗ0Ϯ�8�[��M�n��`�Qh�����WM��zt��6̱�yl���� {o}���|��f��9��9�jBiW��[�Z�����zD��nm]�b����ɻwtk���i�C�կ����،���zl�߸�C�Q����A-��:/�P�;�n����r�?8ʛ-�ܭ���G�!GP��֣p�-�!�-�M�י���d��X?����/���-PH��z�4��OΌ�n|TgS	/�c"	2��pq�1����'��`�=� :�ƇL��V�����r�~��>�cfl�ũ��Me�1*�xm>�ujZ�\����������%�WPU�J�y�
f��:'L���}A�-{�h�&�#.
�M��y���!�qhvU�C�P`x���g�QţT����,�~x�ż_���^[�@�G��(�^��ӻ�+�Z[K5i��!�Ŭo� �.�0���� ���+�o�PV�c�ʇrw��je�;�%@���*�'�)�N��W���߿��ƇS��Ϻc�рAZ�rUO=k�MBH��llT[`֌��:X�g��7p��b,�I�c&}ƒ�Ш��HL�����;TRN����ܪ5o�JPB��3�,�ֺ{�����л�'�hHb&������A�$R0���m�PG�<Q��CLݮ�)��c������'�Q�AP�t�˗�{}��]vY����O/�M�����E��+��2�)�A/���J�&��6��dI�{��FE�3�ſ���|��r�9ϝ�<��F����!�w_�*��>�ml�B;��{1�J�C�ҟăGOa{,�D_N{HT�֯.��O��yt	��V/=��z�_fM�	��l^�힪 �(�U�c��o����G�bI�J�0G}��\��U*h�t����'L�Uk���TE^�M`�3�F��u�$%��M��=�Е�]�!y(m3Y���i�xӱȐ���M�C�>z��P�?�-E3�=����0�.m�Q�k���#E��!�L^cJv8�?a�\����=,�BK�W>�1���
bz�le�� `'�S�27x�f:(+OW��B5f�j��2#��ƅ�H���;�	v�W�b�4B_��η�D���m
�u$[r��h�YA4�ɾ8��lb�M��vr��}.���a���'�te��h�Y?ǆ$�sv��t�B���t�Q\O�z�͠n����
�ek��mnQ���i6n3mpk���h��=�]���[�ڪ�j�1#�X!�s��%oڀ�r���a5�uT�!|��Ʉ\�I��;",Q�3[�/��K6X[l��d^2>�oi��j~��֏�r��k��$0�7!Abֺ!(G�J�ժe�p���Wg!yCn� 
�N:_LA
u��#ɺ ��S�;�	�St� E�����j�zib1M���.�}�K����x����M� (����Rn ��>$�ŨF�h��"}�pƃv�vWqva}eW��MOY�N�9�ƞ�{n`̢�{�Cz�N�u�_��Cy�D@;y���qē#�X��f�^�l��~��Q�l����I�v��
g@k�P��~�"�vz�iT���TX��������-߹2�|}	�'��T=�D�`'_�!�K�| ��e����,g�� ��I�:�?U?-�hk�0"/�d�(O=�DV4a��Q1lp�|C�F�m=L�4��d�t;J�R.8v��旊E�@�+6NiE�q���h�~�`h��X��l��ez�l�W�e�^�vk���_�x��F��ve�%Q�ŤD�V���шa20�]=2}��e�o��H�yQ*jN���\������cw˹�Lyu���y �͒�
1�aTY
I�K�#Y�:�}�-�Z>���+�4%_ڒ��|�E�W����z�\" T�)�wӲ���_�	�N����8����Ź-b�M� �
�o�+>w �T���A�oz�/�߮n���={>㌶�(ɓI�`�I6&�U_�#h�9�%c��_��$M�쿚
-'�����?��t���{%ܶT��U��#��eHٴɂK"�q��g����@1ҟ�jX~'�"u�j*$FF���ez財��sh㲾F� 	�]��ކ"NcG�>G����Ok�6��d�Dt=1��{�Dp}w+�#�Y������Z�9�2x��G��KK��<��0c���l
]�`�fkn�-�����{�4�ɫ�^3e��97�y��i�������F��2�\"㲩��zl*i��孵)�%n�0�bg��sP�\k��z�>������zЇ�!��wQ��(�m�i��τeg�.�Qz��E�a��s�R8��)�NR��-r]�<.��P���I"<:�}��A�_T�M��R����۳�#S[�Q���2��l��>3}��6���"�R�2�_ �����k1�}1^�V�`?
�G�>W�b�m�����Nm�x�-߽_��U'sO�	Mg&��l���u�o���m�&#Ƹ}��Y�
=֞�*!4[j�y�?�ܶ!m��YԨ�+� e\�3(��@
�;�r������,��ѼV�ox���C�;�<q*�Ln�_��;az����qC5�aЙ[uH|kX�����/� �;t���m넜�1 a��f�J�=ۉ$���,�|�!c걦����۸��|3%1]�j��C]��?Қม����H+�EĠ�c�w�Q�u�����-�90&�n�!$Ղv���<V�<I��"2�WK�,�I7!{�}v��T�
�y�t����$ú ��������qB	���O�^���.K�6MO|T��J 2x�2�[˅�}
-�E�al����(:1��7�}��"��<�.Z�®��!қF��7/r��za2�S�����/UT";D�u�l�/��>��Y���~b��Ǔ^W�f	��rٰ�m,��?;�2�a��í��؛�`��8�	1�o� ��	��<���pi_vK 0�1yO���]F[5�X+\Wr�����|[�5��^��4#��&��k��~&V��؏2<�Glo��_�g&{�ΰ��ڎ�@���Σ1��e8μ\O�W�q��K�;��,K�͍���+%���⋆S��-�P4t�D.�X�7�������18S\�X�@ec�2�0A���l��J�A����e6.����a1(�9.6[Lm5mwA#z�V���к�	a�j���Z+{2��F �Ǡ@��u�~���d�T"����(ymk^�"G� uT��Uw�@~8yuA�1���g��ɦϨ�@�Lxj�I�_���ȅ����-ý��u��n����tz���U	�i�O��Χ5+�ї�B̽��>��9!��12z�A��f�b����Z�����ׁ���$�~}�{ԃ�d{���H�%k�����*U��ǏR��)���u�ƈ��I�́��Kg��]��`�H���{fb���g[�ʁi�b���n��i�ڟ��r:`�x<l�?��ߔ�^�aҭ켏$.�y�c������F��_���,�0�5�CnFY3O$��"��ġn	t�)�^ܠ^�)�gbuۥl�%�+��n?�cMz5 g��N'��_.+$h�nm9 �Ai��1�֛�P�nΥy0���>Ԋn�h%����3B���X=��C�dhcjW%�2g��.���]`C�����˲�!�����o��IY�)B`/n:QLwN�IeVn�v�ޯ��h���S�#�o K����Ƈ��_ｈmg&*c34�AS]= X ���-�Vy��3m��fV����o^~����؀�9�0�j�h$��©w���p	�@;DDԏ|����q���׊��!h�ˈ�*�O�Q���sZ�)�SI�h�l.|9��h"��ͤ�P���P���<_Lo�G��P�����d.�j�Gɂٴ�)��}���<�*В�HӯS�G|&�%*�6��T�:C�H�rt�8��
m{Hӵ������.5O��u�`���8�;_���g�>�g��l��kn
�K7�ts���^�
��v���v�K��m��Q��ҌIo��)���"��q"�-h�e	�{p�+�X����mo˙=�(�۬�1��?�1۳i,ȴ�A�ߍ>����?�t��_��<��!T��kހ�;�w�*d5�ˈ	F�N`w�ϊ%wϮ��{1נ�
�r���@��V�6�-_qMHkw�r��s4*�w#`�ڌq��mAP^zS	o�P����ZX2���h4��ܮ�Z�HQbɵơ�,%��>��i�-���U_[+!m��Y6,?�Ͻ����࿷�+�Y�a�O8D�=z@#h����t�ĺ
km�ʹ'̝HB�b���D�/���;�'�"D!�@���偲b�����9�5//����(㍤��|)���
|3��L�[�\��/]-e, ����ꑵp�fҲ��%�}�+J�5��'�������|V�}1�^�v
o�x���T1l���;q����=p�Jݩ:5���/2�����엧�=}�o%("o�� o-��d��=A���y��ĳ�:u�
����N��R��i��%�LȂl֌R_�Q�� �"+Z�hRR�������Zox�(2���w,���N�IY�&sn{P�j�ݧ�1^�YMx��0Շ��FQ��!��6Qk)�fDm�6���!��f�r���S�����Ln�bmz!�z�P6]d���Fh*�/p9�6��Pa�@�R�թ@s�R�19���>�4'�
��L�%�V+ߍU����K �$�I{|.�52���yVB�?F��v�8���w�9��t 7��I�#��>zK�K�N ��&T�{�Zu,���N��|~���y�35��y�1;k�S�����*�T�����F��Ԧ��������^s{a��W_�D�v��7a�>�XE�3��,�g���/Ð0G��L?h�% ���h�1�*��S�k��@�[��T��{�'۶l:��rn'o�zΡ�`gLg�Du*�U_�?�χ��r�l��ޅ���z��.�_`��HЌl���O,�EO#\m���� ���fs�%P�I{}c�N7�_�wQ�h�H-E��*�H8���;W��V���@	;��М�`�X�=�w�]��q�'����Xܬ�3��1j��ôg�y
��I�)X���r<q��qf8�,]�ϑ���d#*�,���_�5E�X����`�`>8��8Ǚ��]vC�M�H�	VKuTV��Ɋ�����~�'���lB?$��F��2D^�a˙��*l_�젫���7�+Nޡmm�_;+i����s%Ϋ�aq5.�͉u���e�6�'�R�p��73[I�e�	M~S:;ގm��ǌ��2��+Z�T�\���e!%�E;��,���xt���]�*��Ti�9"%�x�@�=-"��|�P)�j�d��z��(&�O��,�	 2Q�9m��+Ft~?��\\��m�Z�������Tz���3�l?V��*�s�ޙ�]cnd�:�Y|�wːUE;�ẫ��"��?X5"TL�'�ѣ�}u.;pi��'[�G=���*�l��T�[�i��t��B���g��4�/c�v��H�6d�%�ak.�h4pzXJ��+��J���b��7�.<�aJ��µ�&^#�������r�������y\
��������E�%���s{w�粡dfG$���i����E��%Isb���Y�=�պ3JB�؝��]�N}V���Q�!jao��l��A�L6��m��*��.�njs�#����9@��2b~o��u��]��ߐ�3���.�8iB�*w����`���*��C�W��W���h<̓�t�3��nE��o�F&���Ĝ�k;��0����H\ϙ�ZM��!C��%�q���W.[ј�5e�%�1��&==[E�ii�\�j�k��+�)���(Q����Cx�����ͬ�FF'3���"�qcZ��<���Kc:�kK��hg��w�}l\��-`�K�I��o�od	~'��*��z(��׫ka�����$��̭a�l���φ2�r#^��|���t����n4.x8˜�{e�i�%�N���>�ad��?��;I�� �����V�(�Fb��Ґ)Sj&�T^Ǎhx�x@�~6?��`�k>�w�_\� ���yr���^��n��A[h�eZ���[)U�#�ȵ�"���vp\��r��ԅ�A����
W�f�έ�Ӭ%���qg^g͕�Se�M��=�>��>.�Z[L�˶3��"������c�ͱs����I�F��h$+s�-~�]��n�+	F��
��wD����/��R��{��0���ڂ�2u��Z�ʾ�V��Z���O�0��_.kU|s�q����x}�%q�avU�&�� ��V\3�Yw��\��"�;�9Mu��ҥ.l�����G�e�Y,n+eXIr$Wwo����vcj�W��\[��G�H�%
̭.�с�a(��eCC��1*:=�Q\��]�*y�F����յ�y��<v�EF��إ����J�ò{�T�����g��ih�\���{gB!6��L�6�ˆ�Z�W^D��w�C'm�m8�-�Xa�s��4��)�(�=!�%����^�jCU�T�0����<Rք8��0�ލ��YB�c�>��PK�П�MM�|S ��l��q�-�]z3|<�$����9uj\r�T�WM�<G{�����e�8� l�8�B������yJ����
vu�k5��z-��Kh�R�Pp��������"E�1�:�f��N���M+%R	�&�\�Z�E/yQ�F}�;Uj�8{�&n[*i�W�C2��R��3��4�w$tߛI�g�=�I�s;�x`��e��M�,�p��
�l��_�{[0�>4O
�+���[4�y�&�E��k���v"ﱭb�x�]@� �|M�U�%5,���F3�g��uRY�-n�Бiwb*�(d��H�O�����e��C�j���f0����Kǧ%�{�;���	Y���mt@��dG�cd�i��_F9����/�v��!j����� �Y�s�+-T��܏��\���,��a�_�i�[PLSͽ)���Jι�ʦ���h�Z�C�2��Ŵn����Q=Vb�\I��֒�$}�WAZR��c����nөC9�v�cW��\N����p-���w^`|��	UTM��N�� \a .jM�E�hi]C�����Ր�ct�~�I���V����Gmfm��s���ծ���?���aR��~��mk���ʸ���/�T֕;Ă:W�-iV}�F���n��w����$�E	���u[��Iu;؉G@RoXKAΓ�D1j*�d4c���T����U�x�4��[�]c�$�g��D����O�D�����qD2�XBe�����KK������V�d��}�U�ytq4��Y{��$&C�*\(>��XgZ9�X��/]�;be1�箜�o��QU_}����C���Y+c�]��@����
	@�!�aY[���)�
{��M�D�A�M�b3� �g�p\���6�8���_��m�t`��9��}�'��t���<��1�$�f k\�D!��!�6����)�,� @��Q��`E����%+�I��ߩ���{!~	w,��e6��|W�ew^��R�kK����ª���]c�pfueH�@%ZB����S�̫6	��դF���{��b1�'�c;j��Z�Z/���|��187Z���*qd���M����8�������M�L~*��ixRU��6�D����$5������u�t}�|�e��,߼W�!��
,Bh)��Q~O }R���-��3�����P�X33pTd�����9/�E�n=͜�x��
��`e��|BUs���ǃ�϶����=��b��l��r���d�4�F!6�q��ڨ��箋Vt�&�^�TF�VEkŎ�'q��X}	N��~�?� nC�B�M�0��6�s�5������˨�,�"�)���hZ�2��Ϸ	�?���(Ӯ2|��t"��sh��d�u&S���y�٧0L����G�!	+�8j��r�\�InjxJ˒6�l��K��B�:x0wΔ�d_��睅���M�Ә1�*�ٝ�h�����[v����| Dō��Ҩ'������[Y�ʡT%�����s@
nF/%‖Ry�̯�	��\Ʃ�i�:.�S'�ӶC��«�*���z��s�AS���uH�:SU[���)q�����.����`)0�,��p/&5:₞���t[�s�6F4׀�r�{�c����U齤l�oX�h?3@��Ȧ��S�Q��ѐ�/����0��+�4;�-2\�~ά���	e��[ťzVK��HY�oۦc���g������	Eb'�$�|,6�ӌ����Û�K����- ����/{e�MV�W��Q��M~�{Z4>P�i����Y���N(&�԰sڲ�<@���� b���Y�.��y��퉁֖�k�='*��S�ϙj�k	�����+�x��\��Z�Z�	R�M*�a*��)�����-�I���r8��Uy�c�i�r?�u����nu�U��y���)�to�]�T�h���'�#�:�?Ro��w��3���_���:���^��č���>�o���i���GJ�������@�q���Y��V����m���������,���f2=MA2��J.�2��k�!�T�+�|�`|�����Ö{�,˗���Z��n�S�	�B&���wc%e�]�i���ͽ��7%��7F*��E|�v��P@���
[���ex��
���P��h�ہ�ߝ/�)b���sejⰋ�io��w������(�4�_�^*��L~
����11Ƅ?���eͷ��w9fC�-Ԧ��Kn�	V��A�����;`�Qݶ&5��AZz�k�^V���zY�U$��+�A��G�C)��}V���;�Fi;�
bR����[�����xa���A����N��k��ݺ˴��l�D�Ԋ:p�vQ�b�Q��ex��(��Z��vO��FL�YW�~3�ekjm�[�Ъ��HRy��N�>�����������4�;w��K�������%PA�1|��*I��`$���C�B��2�3C��Z<�/:�=:U�g�4�X�\�3<u�o����O�ZÔ��NL�n��OU��; �C��ӊ�姆�W^�轑��6�!�mHg��;s��!ڥc�q�t����|*D�bD���Z˺��� }�"���rN���=��$"їA�ф�{E�ԑ�$	���-3M�A�4�o�}J+�����/H�.b?�)����dj�a��}�!���p:�MՌՔ9�G+Hs��A��p�ȆQ��z�`�3����ޡvV��J߇mJ&@G�OW�8��X��̋MY�2��:�lB4J���^�l��J[JxG��!�y�U���&�����"0LFk�L��͊K�� �Fby�}'Vc�_��o�݄���N�!����[�A�b	���"&��Ϯ�G�d!9:"]}�?�4�����'�\�R �=��XB��[�#�0;���9_Y��of�����{��yay&��^�G��:y)�y1>��M|��v�,Zzi�����-�����Ҝ
�b"1�F�kǜ�z����a��=�MgOb\ť��ŭ�sT���%m�6t��2���?��W�eӈ�Ny@��!ZB�\4����6c���v�â%�O1*�;��Ǖ�f�0�� y%��r��2�I�/ꌢ�
C����.vh��_ 3렳���һ��jwp"�od��?�٨������$�[ӗ��b��J�u�w�ѓ�a�q�'	����џбA�d���(��Jq�@?2�#>�UZ7�ʚ܆���)��+��{D=<���g���r�0�T�Y�O�n��I���q�O �᱿!�Y�~I"d���`���tf������
�����+�T$"(�=3�`y�͖������a��~��K��iH:��	��)�D�v��F��\��:�|5Ym���@��&Gv�ɲbl���Hڄ�8�|�߶v�껚�+Ve�8Q��
L��E�E��cq����ht���c��Bf�\u�^Sr���2�zG��j�(�V�4K
�]V�Ha����Tuv���!������#�x�� �2i�c�1�S�3t����f+(��;��̨���R�AJ� Q�_��4(ke����O9�t�(8L��Ў��ݧ�@��p�ǳ�"|j�4��ju8�#��"㝼���+��v���j>X�8�Qw���kl2����4�XIP/Ñ#�1$Ltgo�QG�̱\��毎���nh�/ZB���#<�5s�o���c�bz� �l#�qh���:�U��7�
x$�����<�v\�e0�\�����Y���A��Z�9���y���7����yb�����������f� m�L�d]�Q��z���5v�Ƭ�N���5�h ��S2����(�&b�<,��[�[_O2F��Mv��L�N#(Z�N�g�Ԧ����N��;��)4�2`c�A��U����t�<�`/�����V�t\9��V�!#�v6�W�@�-E;E{�V쀹�,k=��{�f��ܳ��PB1ccM%%5��Q�WR������z�r�H����
]���j�� �3��;��,L!l�<`�k�`�'	��D�otf�cւ?����H���-F��af�VkTʙ��������ў�������]�6S���z�1��9o��ݞ�� �+��j�m؍�u�r�>͂	E���vW�����p<�vf?�vG�'*��w�3���$�@4	Út�	}IS��^�Q_J�^�2�Y.oыՖp�׽�H���u��d��G���ƪ¸���P��~���'�}D�5�-\��xZq>�����/	*+1��KӃiC�态I�0~���s�M��`Ot�1�¨�L���ē>4��4�4}���F�Մ��Ь>A�m\�kp�T2�6���8܇_LkQ�ɮ��f���d�i_��D8pO��|��<�zA�Oi�!e���Yfދ� ����Q*�C)�	�zw����V�|? 0��|].Y������/�=�����8/�bܘ���o�=�yZB��D��{R�:�$lQ?�a���t�A���f�!��n��~"��/�5�aZ+N`�}�4К'7���4��|�����\�}�/�Vm�_�f���en\H��_�1�.�Ehx�AC>���ե��䤕��2[��?�r�p�J��{  \z%�Yx�ԙ$�����؏CvCҏv�4��3�;��#X�
53f�_q�nL�|Т�rY�|�΢~�����ZB�T�q"1+0��"��C��n��G��XB`5��I�_����2�V����@'�l�oOʦ:�Cy��J[Y�R2o򠩒�t|nD���;D�V{�s���t�_�C2��
b�|�����5�\�y1�J��1h������~�q�$��mW|���K��f���lۥf�B0_�[���u�l-[7��m��X��V��OfW�V�7~�t��R�@�ƌ2PD�o����ՍV��
�pY��p�{`����@}�t�0l���X�]+'q�%��L��󆳗S]����x�7���3�}�lL�E������#"���R-a�=V���c���od��.ѭ�#
��XR��oy��G93b��"n�d2]ߥ��AXۗ�6zH���O(ю}S%��ؑ1N�ү��f>0�_.�qC�K���ۂ��ANy;U��ˏ����o�:�w�?�"Jl;� �*�l��d��R72O������R��s,��������}�M���,['��W���+1��f�|L
=ה2}�Τ�&MY�c�9(U;2,����svͩ��U���'S�CRVp��ז�P4��H���CCn�
g�>��P:�X�3���f�_n*���h�g�lu��o�(#&������@j�1��sa�&3�]�+�Y=��߭���Eڭ�V�Q.]�R�q58�-B�Za��a�nLf�[*0d�QJ\��o�GZ{�`�\�=�M1!�}$C�h��'aN89�:��u=�s(oJSs$��'TxR��eğB#N��j���S�PiS��U�\�be�ʔ4��d`x9"�5*��f_�2ry-6�q�B9�UЀ�6����`�5oPw�����J]<W'0;��G+�J`�bpF�O!��g��M�8������LG�֩	�Z�
���̧,��ۢf�Z��33��%����0b����O��V��f؉�	!'�1���uqi.i����t�3�;%�L�Y���i�V?�E�\��V�O�si���w��y���u�RVGY�,��Ҍ��SJc��N2´�h�K]������ϸ��q�5��*��2Ҧ��%��l�;s�h��i��CJ�s��+��ڿg�1ڱ>�#@pGσwP�tGz�U�����.иz�f�(F�#�����Nu�OU悢}��V���;x"�Y��h�ޅ������k6��b��FA|��_4��X�3N
��d�pLܽW���+?�?>F���?(F�|�6-�LK��О�u��o�.xʈM~��t�`�-5���%�-;����#[�ۊ"��^Ҳ�21�b���V��X���g�����(U��G#�u�-�Ƅ�� ���h?��+G#!�5����3L����trx���s�����A0�~}�J�&M���5�S���_���e��D���T�E*�#9�۞�H{��9/�O�a}�����a?v���ǁ�ŵ�x�yG��b6>HL�d̪'7��|��}*�����QG��yQt�tkj�*@��������z;��` H�%�O8���m�b�I�~n~l�:���ݿ��'��6X�k/^�n߄�j0�Y�N�>�q :Y�e�ӑ�n��t��01(�N=�y֡*�P���dhq�{+�s�=QJ<�{���x+�����
×��(�}�D��ZaG�;����Z.:�̞D�N�Z|��LH�kW�2�X`�/3�Q�L,�3��J�
�׊��4A���������|��'�_ԃ!d?��ʛ�@A<�$�p4�QZ��{3�ȹ��]���JV�cJ�W�s^�_�6y:1�e+?�~X0/���	|��<�p;��rRG���4�F�����;R����K4�����Lh��x�}&�33MNtA}�S���ף�P&8�*T*�T1�=�,FY����/9�vS��tZ���kw��*m�z�M��#u� � 94�Y�Ӿ4e6�I��4����m�:�9��<��7�Q@e�.�飛S�3f���Ԡ dƈ��S������@Ij�#gm4<+Y:b[3`*b/���Kp�^1�%�ڼ/d��B�-��� vҏ  ����^����L7T�FP�2 B��`��!��������w���XI��������@�"���U������Vc�m��l����`L�ζB}����{��8��5@��7/^��cN*�>��T���j!�O�y��vp�v&�.��'�'w������?	?ҦC������a�cB��耒9o��	h�x���qj�h��.)tA�(�^�;��\�~� {��Iw茆��
��¶�	�mp|';{+�m6v���`64%yM��nP![��q��������B�&�O��d��%�%6�8@�f	��iA�����cP���(~���� e�H%z�b,����C:I��Hh��Y��+�j(Þ�\2">n�RS�6_=��6�l�R?��i'�#���"Mc����/a�4�%�˻Z1Q<�RG&�$ن,H�����F��\�EJ������a�b�2�fV��O��Y�b1vN�L�m���SD��ց���#���� b�¾��\A#���<x�W+e:����o�5�5������ꢄ1b�IW��5��Kc��:���'��n
]���J�vrM��F>,r�6H���W��M��o�Yw��%Ja1ݝY������qp(}X����h :��I��Z����55�Xj0?|����_K�X�����9�8�E����\��&�L���}�X\��1�䮹kVl@ G)���KW+�صuZ��_d:������@���=Ү�8C�1�1�$fF��d��:	������9ҾU�fnH�ǘ�#| ��M0!���)�u���N,��d�Ⱦ��)$i��0�|u�A/U�2���#����A\.�;��eJ`�]e&����b��*�����1m���x�`n�X�����5'ǹ�;��?MeA{��:R��2�Ɩ� ɓ�M���i����s��]aO����q!9%�)4��a�s��Q��?�}�vf�^gvx��e+���5��x�ק"q���q���3v�yT�:o�Fg�o}��A���X`BnM�ҟe�*�z�jԫ)��kNZ� m�5���ۈ$R�k%�uN�@~�(�E�g���f�Ț������ ^�}K���H���Ӆe�^ztkwg�ݘ�|�+�����d��&�bu��XWj����i9,9�IB��O��:@�䶙�;u���l7�V��K~n��i��a�Yʸ�
� �6塹�UH`���4����2yj/yv��Ž�����Ͽ�u�nt�{������FD^b��T��& 3�5u��[�~�7���lWt��z�$��w8�/E�CC�'��C�o�_���od�(�$�v[�5/�ޔ��n�y�o[����t%EYm��J
�H2�}śv�c7�S�X�Ӯ��Gv�5�"C��p���81�Its��p�ۦ|L��7���"���*��$Ԛ�(�!p4��7�w�ұ�F��F��sQ�$]���uT����G���]%-"ڹ�u����ov�C���ql妢(P��T�SN�+΢���I�����3`�G�f�W����r�1�?	�� d�]a\�gy�J��U�"�d�[�ē̟E�ѯ;�0*�$�8��v-
� ��x���q���(������{|5�/��\+����H����w��5�ؤ�E�N��v���*%��u��	��%,�8�k`l�Y���r��.�_B��B��}�z&#Ɛ$w�::'d��) %����q�Sy"��=���q�M22:��Za�,N����(��beʥz)3֫:��\��N�]�G`=�-�A�R�E�X�"��84���!*�ǐ?mr�nX<�?���2m����{�7����Զg��S�?~�]Gl���HesU`�6�\��	.�{i�@]�<O�6��
?$W�%�0!�Pƪ$�I�٨�F��{�9T�\Lm4M7]�,�pG������;��Ē��,{�|��{Qh�[B,�H�9�f����3�\toR�W�Ì<ѿ��.^��JW�����Z�x���c�):NU�����fsF�-������ڼp���7��T�ݩ{�ΆN���YӁ4�t#��(
Ю�H�SH�]	�D����# �2����p�x�K�6-����M�\�w��k�O��m�1Lms�� Ym����MI�ܐ׈��s�؅f�BE��z�-NU>�1dݏ��q��]�\�vq�C�i��	x�yVg�js�M�A���Z&����g;dX�d�+��'qq<���աb$��*�e#�]@4�W��=v�e_:.�*�]�z���+������4����#��E��7�V���:�K�4?,QP��%dUH'���ZU?b���>?��5���G{7'�R�t|��2)/�P�[�._v�g��\���YVud'�I����cT�'�Mx��AA|U���}��g�b���� ցB��X���y/�A<#��{�[ZT4�#A9(�����I�k����nŴ��{bA���WP��;[�X���\�����d�0�ɰO�Z҉�Z�������ޟu���$;-��4C �U)77�8��/���������őWw,�Ȱ
���B>�I�EiU�E�EB�s�|au�ޥ�5�x���Y��h1kP��Jfs�5�fJz��}�3O��J�T�d���I��RzR%ڒ�Ni>��~�r���Z�ƪ5�J�����WA[ar��!�;AC᝺��B�4�D��s�φV�҃�o5�)D!��ӭ5����d�F��m7ݹ���z�D1�����Ƶ�)�S���S����Iu�f�H]&[^*o�=FMW+��v��k�#����'���~>��N�"�*ɘ&����\i�����QW����ds��Q�N[	K�ʛwzܻ�r�f��ᴴ�6�b�>��M��j��~�f|���&ֆ�gu�b��딐�g�����b?z��@��u�ƶ�io��g��^��Ϧ�6O%4տ0��9t1�����=� �B^֪Wy)���+l�)�Ԃ@����������ʫ+d����Ȁ��p2���S�p�/�׋z��¯�/��d0U��h�Z�e�D�	�(-a��������Y �V ���1�'����;��0����n`$S�}��t�b�y�����)\�e���묐p�i���1U��7m��H����S�֤�ڻ��(��:^,�K;G7�!���)9��rP����N掹�;$�V�,ŀ2څ�ͼ�
[������hck�ɓ��(����JvK�Tpw��J_�mL�p���*�9@S�'�B��A�� ����\6S�rKO9X+t�}\c��avl������O�@أ�V=�=��*j�3�œ̯� ˶q�n~o��?^��[�LY���[�;^>&����_�l���+ÐD�:�z0�'�;�O��f~��v|��j\�������6��"p����"�jW���&�M0�y�'S��4��DP
G�2�o�������GV�;�>��\�kxŜ?��=,v�.vG�h(��Vr�t�YL@f$��	�ކ턺\ͼ�IU��WY�$1�߽jҍ�P��Z�µ�٠9!��MZ�w����ȳ3�;6<�_�LY&e���K$�{�(�ݥ��c.jˤ����[ۖ���A%%�����!��r ����K��A�~�P�bYu7t�f�����Ǉ|���©�W/�V����𧗘�Nɳe�5H/{Ba�P[��&��Jp/�*�2�V��$���m�L�]9�8��}tŲZ��|����[�3�<Z���6���&�qd-�0z�i�/�@�ߠ�'.k���W��Ϊqȃz��:n�|7�쐓�yt��Y �����Q�2���|�Kpސ�=L��Wr~H���b�GGb���JD�\�/9f�
q�HF��i�BF��L@[���kuWq9= lӃp�u�e=g���%~��߃3X1x� X$�b���p�p�sC�]�����8�[O-�ޢ>���J�1�?�m]���$�w���?�ŗ��{�a���R�	^�(bS&,�
�}[��䤺�p��s��5FX����%G(�(�aUy� /�Y��yWۉfݡcO�}�*|qd?���f6��\n�����\�5��Fm;�Ųy��m�����!��� ;� �j�x�@��``Rf;Mb�Ү����c�/�U$QE9��X�v��X�9#"B��]9���D=!V�Ƴ9����jB)��̲\��\�V�6W�ӑ�1���o���*ŷ��@�h��F�21�꿂/9#W�ӿ5|WmC	#��jNzt�K�2���γ>K�]�>~gk��Ć��YS��1п^[dT�s�D)�'>P��$/t%�D�=#���xQ��M}��:�
#!�SH�(�j����� �p�x��=�i� l�=+w]�w����0���@�[;�d�F�f���1;��iu ��t�V��H��y��f� J�Y���8��	�#�=���`�o�l����x�B��ȋ���A����M��s����<����Xd��M6խ3חj>�PHН�s𑐎��<&�B;�Q�<8���ȘB�?l��:P�DK�v�dJ���av��/ǖY�R�ii�B�P�� �a|�o1+f��RG:2�-����Rx�._^e�c�̰�h�o��<oL4�n
иy�qr�v�ڇ��C�{t(�R�o����?��i��ݲ##c�'8��6wnS�܍��0�䠲u2�����2d ���K��Kȉ����蠹���Ba�q�®/='P칣��)�hO����Ao6���D�wU�᫏�VW�X�x�7�!0{��o���Ѽg@Lg���J��5Lk�P+U�]���$	z��9A�B��9����fg�6�M:��{o�ﹲ<�m�ha_�t��z����Bc/��X���1CA�c�t5Y"uX���^�&�*#��Z�� ?yf�����D<?+�@���hEV��c�[!���x7~�����g�=)��5m`/�vSٹ���M|f���j �Bֆj��	��U�Ks[���Ի+�Y����̥����`	7g&=�C��T��w	ܞOl:CRQi�����>��rV^ʖ�� g��~��#��]�"8cw��N�;`�j��W��"���!>
���s��`��=��?�x}-�w^�Y�č�E��!��{e�#}���%>�5�e�\�р��{=�	���6E����|J��pN�����D�_h�(�! {�Vܒ�ܔ��4Y�8���EV�Cİ�C����LP}fwc<)\~d���i[زګ�n���n�	v����^�G������{~:�Z��X:�o�H�R^��8��7���
@����l�ᨽ�
� E��(^C�s���A'ۤ�z Xa�Wx�䕒>�����p}p��!���2�*� ��Cm�R�a�O$��E�:�_�=����1mr7$ؐ̏N��@X�y;
P`�b��9�?f�gP�N�/W�y?��w��.�I���n
��a���"~�Uˁ�b�����ʪ+�\��L��;i�����Je�ґ��q{p���4����3��\�-�c����u�A�/�Ñ��n�4�:!xBæ�C�������I��Η�ziM��Ӭ�v� ��a�3�R�Z4	ϩ�CُlӉ���=ӹ>�n8Po�娘W!~	�FX��#�Z����lUj����}�GA���bp��kj$]�3���.>�6�cIԆ�+�پ�"~��j�ɛ�ok 2ay��f
���+��v�.c��W����=e<⛤��i�_
_�/�<���fV}Qd2ĪB��U�Q5�H��i��E8ٽ��v����
�x	���gH���\h����tl!��(C� ��5��=>[��[쏾n���"�#�.5M�MGܐ��ZD�}!!�EN{.U�;�<-T�+��d��U�ܑs2�����m�"�CV6%�h�$����,��m$wCX�J�)�������M	��=dmT������9/7��x����1G�B��:> �q� ��f�A'Q �N�ʽ24=�t�D[ڦ<���p���0�ox�m�B�I�ݑw���4Բ�%�İ��t���\H_\��cc	�J�\��y�0�!U�<e���� �Y�����V�(��D��<�7O�x�_�x�S�ޥ-P��yϛC����D-�2V)�����\J�5���֠6�^�-G�mM`� n��d�V����D�\[Đ��I�gV�0�(���&}x�nb{4E��2���R���0�j�	��/f� �L���d����Ã�82�P(.Sm�/�U-�f,�Ї3��aF�I�������3H���@OK�c8Im�=e�_��m`�؍�[���sQ�rz�E2�B��
窃���~]���4Y�|��;�[*�rF:7�I��z%�<9B
P:L{����)T�������ߌD�?��J��m��%�m����	᪹��y���/�W�����0̖F����r==������b���*���率>�c����骅�xrAPo�;��.��,�:r� ��ߊy�Bf)H��[��� l�P��-ƈ�D�:��Z�,mB��j�A���Rϡ71Nn�/�ϫ�Y[�'�E纻�T�+�����[�r�����G~�ǂ�>�TX*[G�kw�Ө!l��d<h�:�I�b�$�x�HH ڪ��#	z/���_�����"|v�-���R�E�,8�k���柁=U�~�5d��ͼ#7�V������8Y?]JR��C�Wo��Q�<7��Xp�_}�1d��AjT�}�.�1���58'�y��*���ց�C�؆���n��&ބ�n����ڀ�T�e��ג�ۧh��r��w��������v�y�	���X�W(��O�q�7��X�� 3Ƴw
S0���/d7s�dDe�1G�M���i
����&�9E�g���,Q�/���W�W��C�O��!��Ha�sY���?�|���w3�ino�+e}�������!~ a�	ٍ�*R�+`���uf4[�(�Zf��˄�GE�������8���Ͽ#�P�w�?V�sdxeQ�f��;�[�mt^�(��V�Y�|�*F�{��5P.g�P �~L���3��|և��2�;�b#A����o{�f�6.�G0ܒ��Ɍ����y.��"'�j���D���
G.�ƪ���((w�+ݘ*�<�����J�|���j��峭�r7g�X KV�̲S]�U=���Т�־I�UԽ�_��q���H`�7���U��DP��T5j>�.b�>�`���?�"aL�B�;�����`��r^����?�V��W����FS-d���lr�J;Ev�R�,��%����Wá��D�Z���EwS� �f�\���u�)飅�_�!?�ؿ����1�t�"���U���*��R�ѱ�FV��x�z�#q������eD�[�&��_AbT�s�3�GA@e���%��KD���8�~-JO�/_����M%ҥ��X�1إ��g1�V��:��9�E�A��O����aA���~��`���`�����8���׿	[�<ȄJ
/�r�tf�8+�����t��P}v��X�Z����z��R�ϡ�������6�z�E���g���9mJd���u"��z�2^^�{$7=����YK�f�h����h�*�Pέ(Afy�~��jd�։��)'��!b��q�s�UӊR�/��=��?���1���l���;0*��T���*���b/��(���
XV�J5�}�Ew���u} 9Y�?���$��%�c�ԭ��vRq���:��tW����iˬ��&�\S� �GH��C��]��T/��/���ȁmHb��r�Qr�3���9E
�l�'kr���*,�oQ7c�B̲[����>	j[k�|�7�M�_)��h�	�"1�}d��oZ�=8*���h	�$.�<yԵ���泀5M3AW�M���,6�����Ij��t��rϺ&������r�W��%a�O�H�~{��8���߯�3P��}�0�#�t��Bh�t!���qx��1J.�(Vf�"�t=Co�q����p8�s8�ߘ�Tu�9'>'!� .������|X��>�a�jl��so�":QZ�E���X=��1̲�0���F��m����1�J^�t|���<8�?����Q K%�#At���2��}L�K�E�ٹe� ٢��˩�6�*;Ӳ�������gS�C��R�8�n��ʭ���ѳ�*/x&��Ā#D4_�C��n
+	���������Q2c�� �!Mg��c߱~!�}����Yz�8�b�7���qd������ ��S�]��梟���ޅq�8n,3�r�=�e�=XT�̷x���r��z\�[8G|���1�Q���f�+z<0��'.I�y����d����2Yƚ���4�6�����lU�m���'�B���H��	�]f��*X3:�l(U���n��j��ui�=��Q�|��e��Q�d�9��#��E=�R�$Z�������Z�a�� ����!;epÉ$�Ro�����ć��U;_ٔ�2��+o3�z�DӉ��&gt��y꯫��<��H�x��)Y��4xi��_�ֱ=N��!L��cg�D֮�����
9��X��$�;>��{����2�x��M�2�~
��:�jnH��
x�H��o�|��v_�["]�O[�&�/,�ϑ�-!��B�II�-�УVx����ɱm�+��H�J "�'e��������P��!��exA���V��Y��rO��?1����d3�=�-����v���$l��᠍!yHX ư�$��r.U&��+p�xQ�XI3�J��|aV��uдꗏXye����S4L�����N2�Y�/=ZLР�n�d1E�r��~JWK��٭Cfuő�������{f�e�S �#���y\?xn'�n�� ������'~ٵ �O��9l�̓���kxq�[�X�}�j�S^Ag�WR��/MM�
�r��a����0��R�{J�KrIL(RH#� Y���B\�I���պ������~�r5y��3�2�b�Ĳ#��fX}�e߸��*������Bo�GGs}1�L�i���V�r�13�/0�!K�@�!��M1����U��Oз�Z[J�`t�S��V,Rdx�ns�;�5^&nor�j����^��4;�y�h�M���vQ�%��i��:�p��'I�~>�T��������L� �u������a�RL��b"� �wtF6: d������e��{����ЌIO�~�"n=1a�D����I�6ݲC��V�9τ�F�Ƴv�}��UT#�M8�[�H�8yg��<.���">W�.9��7V��\�A�������_8Bո��u�;MdC�������0�%���h��Ô���vc�=c�����"P*PU�A/���Qh�^I]���~�\;%�?�7ރ[�E�^>j���}#��o449W���G�?J�x�"�j����K���j0�7h&�0� E�M��y���M\�+�K0 ��p�0a%V]E~�m�i��L�}�԰���AK�;���c����0I��������G���a��p��|�|�ڥYi�r��\X���1��̛Q�z�o/`��h�!j_Kgm������Ȍ��ܷ��w��a9}�{���2�ܼ�f���jg�����"�6������UΦ��?6�� 9I�1l�=�3��ᛋ3kwwG���`�̶�<d��.�0rop��E<[��ۧ���+=��{���Eu��_�@�kڊ�N��Mɋ,7��5�M��o��dyqO�Ɵ�y�c�Y�į���Hؗ˰�|�.�"��aB�N=M�3z�c�k�n�RL�c?�/u�5p�B5]E��q�i1�$6� ?�Q�{3��WCi���G7_
�fA�;�G8>V��w�?@�>�[f(�ɧ1�bB���Fx,�P1�n7�)��"w*���I�'���_��~n�K�~@��]bf��Fu��.����)�-p�⋚0b�JA<�� g���*:�Y��\mF�J/8n�x(�ݶt'����C*h��@̀|�D����E��Z5�L�&4]��e���$���g�n1l��Y�<�?�����p���l�e�	����zČ}����=}�I���K�}�{�<zR�{���"��^�R�r�W�on ����K]��X�7-�4��XoW��k�o��S�D�����s�����9�r͕0Py-�Vk.%��XK����}�k��Yɠ�V�Vz^��9;7��n^n"Ρ/�'�#�CqI:Fr�M��xxS+�Z;��u}mH��Խ��҂u$���-7�s�D��~�T��-��(�<s��Pw=l;-���6Ey��[0���y��ɪ/���4]:�^�d��p-�-��Jr�-�d��3�� ��:b_�O�!�+��O���~���I�a�4�
5'���.�[{#�����0��ki���	~U�e�+(�~J�Wmg�B?6�)�)g�Z�3������u$y�Eٗ�N4��ӳ��kΗпN��&+ˈ#`Q�$f�c�+���L�w��3���R�X�h����&�EAn�J|͇x�ܷ��-��
[y�O0���)�;��Jb�|!��a�qѷ�|U�����`٢��XYn���#U��q�N�S���f���k�>r@c��>x���#�ǝQ�u�"�_/�(�ݚ-uQhu�v�I��})}kd�~�_�E�f��F�3�����J��qn҆�����x��=
\k�����I/�ed�>�Gb}�1ٞ�#w4��,Q��-(^4n���_�Ge�D�֫(Nq/��b,~ɺ�/�(�U#��z�ju�HӃ��e
��mj�gm(��\�<�N�F,N�wƱ�\ȰžP��_�=-�K�]0�a3�l��d�k]�e���|���XQ8;��������g�Hyl�������6���)���zx���#C���Zm�����"K�rݶ��	�.}����Y_;'WRֱ��΃�"M�כ�	a�\=S�+$d�p��^S�K��e ���V�9�_�E�2���U`���V�x;�-A��n�9	U�OWO��pUnȇ��ti.���0>C�S?��+��m1�W��9�p�Iaތ$�8hF-��1g�_d�J0D��J�ؽYA
+i�j}��vu���\a֔��^���>�@�Hzj&V�7�z��@�|�eɑ?�����K�J�c�D�B���v���\ַ����$1��l��ä�_�7!��܊�Xh6N�'#�����{���#�R�v^�;U�o%��'Y�o`��aQ�h\�/|Uh��=��?�m<�X����`�4�0���(�]֙������b{7U=��m43O�9��q6}��,�`��!7B��|����kx٬�YR���9���4[�ւ�[�]6W��!�8/
2d�[����Ž�����hP�������g��Ss\�jCU ����T@�â� ��f��>l��	yT'����X����^��F�9j��S6
x��@��K�Ww������U��$kE��Qsȉ~�)YO+0���:�
�T^��p�2)�h�YY��Wy������w��1��D.��umhU��~�k�� GL�7�@q�X��HV�PX�"�!�R��S�o!Nf�NW��x���E�X��=sێ�����`�k��"z?����T_�o�{��N�Z��
�z�uY9>X����H�n9�MS�Ur��<o�}C{�%�+� M��T���XtZP�b�^��⦀e?uV2~g�+7�n5�����ű��0c�j;��5}�O��%}uԏ�4/�0r<�f0�-�Sć]�hJ�`�+' ��i)�J�V(^�w��M# ;Uk�O&]]P�ռ�4��})�!���l� e��_V��&�~T���/��U�+��j"gEd����qzX$1��m����P���uu�^�����&0���sw��.fahhg��c����g&��jʈqNA.:�~�lU-$�v��)��c�tCy�6�!����dU��nm;��A�(v����%S��a�^ �I��{UiE^�t��g1}?R�TV&$��$Tt��u@����?A������>`����<�t%W$T�����Q�ڇ��?�7�ؚ*���yjF�@��j��\ג}Ʒ�x�;��#:���mj�r��"�g�lx5~�)�oRv�'�J�y\jHˌv���T�,|KSu����3��	����e�k��q�̧��p�b��}# �w�\��:I,��Pc�}�)?���SXg8#�f�J���l�S�%�����T�ॷl~id��i�c�e@���~�AV�v�$}�?sU�����E�@�IÓo����n[���*����nt�h�V��b#���UeөY4R�ؒ���?��a�
'cM��/�J� �ߊ���7��+�]�����*�K/�ڀ��R��V�6�z|�!C����J.��Y��C�βQ|���		�y�jׅ�#s�Q4w/�!y���B?n�T�z�� ��������)Ty�I��6%�@�v�<����
x�s�$X� �ձ6�O�_:�i/�9"��� �����Yb�����b�E?"w��/m�o6m��������承%���#��Kq��no|>�?3jt�ܹ�4�O�	�B�z(lé:UI�*N�D��=�qҤ�"~��)�j	�=/�1�t/_�ՈS2ɒ��Cɵt���W���|ކ(�
�iL�8�Ѵ!��UQ�H��pf���!l�+�9�`-?z��S"�䐠�m��2���9����V?)��Y_5���B�K���m^�N�H�W��4Y�;��beY�1;^@�)�M{��� 2�8m�������49!�t��p�+.}=m�-���؎";����V)��@A�^I'��!��@hL6t�v#��@�����vj�D�Y:8o�^!V���}:������t���_� u��a-�����Hܬ7}SױI����k�u�S�,� jD�F�[��6�=|��p";pЩ�{��wC��ź�f�#��7
I�u�_O�l*�e�F=e�Y33��&��@���Ֆ�1 ]|������5-�	�Z�C�|F�]��%�Ču�i	6��;����Ϲ"(�����[�NL��P�&�r5LzO��Q��
��"u�g<s�c��x5 8�Iuh�oRy�)��k�V�X��ƥN:>)���4�b>��}�c���za<�=�e�v��� ;|&ǳ�{*�k��-�V&~�s����%@��h�V�lz�g�������r憑;7�DZ}4?��_K�q|B�������]q�ь�qF��G�,=)�] �C�gw����/���kO���"��}��B��.��_��*����w;�� ȭ�b���i�3Q�����Q���U�va���; �:�Zv%�,d9�Q%$����x؅�B*n
!^�?��\w����@檩V�Y%rJ����r#�ʞxC!������ė�.����ת�`��F�� �����!Iv�c�R|16&8�<����>�JV����yK��&�4��QP��2/�D�|H�6������P�1o.U��h�M�y�����@�rh��1h����;���Y.clc����m���xSs�8�C��l�k?��I�Ւ�e|˟�vd��"%{�0p�놨6���_d ���1�4}ō^�y�C����:|P���H���6{�o8�P�,%?� :�Y�UDl��D.������lݸKތ}6�S_M;t���.�]��w.�8��X���߫+ۍWЩ��e��	���+Ҧ�y��zJ�����87ZD�q�R�
?i�C���|%��{��-(�`?�L|�m�8�XTH�/M�C��r�AtyzԜ�Z��i"���^���J�lH~P�3n1BHR����Jxz:a�^�G�`�?W��}�,.�-Y�TR�E*N��<듘<k��9������um����-��� )�N�Ӡ��N�#�
XtES��Y�z��w�u��0��֙�C'�:�C��sN��s�rQ��	�DU�I�=�$5������ޯ:苴eTh����)�B���0zלD��GjЄt�;M�kW(�ߩ8o�=4�����OSQi�18�%O��O��3c�<��neGQ�ɬ�|�K!�J��$��U�_%���΄�ʎO<W�����U�)�����~P��q�q�̦Q,�{3��1���%ƙ��qVQ��'��I9I�=�%�r0��˻�=�)��E�`�����Y����̔�<W��M�գPt��C��^��C|��dN/��6�\�L+�c�|��feI���. =�4P��W#4Z���F��]��[�����\��kN�B/�P�xU����8@a�L���g�*�����~��ON�� �u>е/�PWL��*ݻ#���E=H������;z�16�p��ۻ�0������f�x*XJ��DU� �I�,t��~�ޗ����o�7:2q�.��[�Hi=|�0f*�n>����m��`��D����CYӭB��8Μ4���^1���ӛ�����C�ǎ���Ʒ������p]>�~g͈k%�÷͢l�F�7��D���;�Ȗ������G�����J�Y9��g�;�`gm�ZS��Hv�!���e�4_A1�Z��-�\��{Q���1k�A�\�}��i�jR4~H?ҫ2Ce�}~Xߦ#E�®��d��Od�`%.|�D���&S�Hl{&p	V��Ӯ3Q>d寝�PH~7�/��֤sY5�_p���t��
딅������vukHؘ�Q"����BN6q��h'T������!���*KMx����o��)w�*��`���?�K^]&;����Yj�d<צ��P��<�
�-���_lZ��]I��nӑ%)��9�O媄�ܽ�Z0�B(؅)+?�K-'�i��'�3i��]��в�(b��)�1�S(�ВӃ���2"ݽ ݦ^]���� �CP���Cq�ԏVax���{v%4���1�'0�^`�A��ǽ��wq9��>0*�wаI#��e[���7�W�խ~Mޙ���+�������0��>q/�`i�ejf�oDO]���������;�kd[^��n���Mu���]i��h)�G3�1/k��P���w5QJΔ��a�_˧������L��o��[Gi���6�O���ݹ�֒ �h��p9������K�
���y�'��H�vP�"��H,imy*�n�y��Y� ����6~��L�����C,�6�nS+H-��(-��M�����lgf�W�uq/��� �^-?�q9t��?������*��n}�`U�H������N��ѢL ���*=v<b���c|�g�0d���r2�%Y�����N[�6��^��]~�a�E>��4�v� �c��R�l�Q?uS=�����T�Ib�*-o�~�:@`���b�&��d_�c�?�R�@��-��.�_&X|�l�������-��J��m��&����ǖ ~7��~�{�0޽@�J[�$��`9�Z��CPC�D?l��ջ>��bˁ<�G��=k5y����W^c�@m������h�8G��tj��e�#�El
\,&�S���x�ה��Z � wg�5P�v0���Q��
ddRC$Y���Z��W�a�w={�$�~��'<bm6K����h��4tg^����߅�F��j�=N'�˛��v�Z'�o�8Q�.���c~����������N]�@֑D�U�>��L�=P�5�p�{(�A�cj>�V��R���-r8$�};
���P����������؏���-*�$4��	�(����R�B=ʟ�����G(4�b���j+m���B�(K��1W��$/(O��?_p����H!��Ej�'R碇`r�@��0=���!��NDȦeI�\q��&�.w5���P9���d�>=�"�ӎj��%�1�KK~��U�?��&f���Qg��^�N�j�� �3n	�n1�@��	[�d͘���+�;���c��ͩ�wp�D%<u��O���i5:m�ǹ�H�/��"1�Z�St�h:�Íf�H �tƚo']�t$����Ѩ�>��,a�v��NwlF�Cm�V�d�)݌�C�����)g�>�Ԅ22A㰲G�T����/�����s��:[e67��?��ʕ�.<�V�GF�H��6s�6��8�骚��la���N�3��vR�ƏG�*�槴�>o�!_�,Q{4�v��K����ˮ��|�H���]W)B��һt�;-m�ri��,�����N�b��F�>1��)�����Oj| �G�S`���uջе6�卵��7���b0a�Нڑ�S2��mm/t��3*�-c S��E�eӢ���ɴ�e�D5�x�*�Sr���qy�;������A��"c�p:��v!Wl�i�������]�WUg��p��1�L�ψ8Cy��	�~����4S�kt�<Q喛DA��^j/�y�j����~a �H��w�0�8H��e�Q��7��P�:�^����*�u5O��>0��|s�}�8�[��г9�eSPw��we�� �2X08,��ռ�.��2�h����`�^�?���)x>���-A�%CZ�T@�v���1�B���-C H:�[(r�tw46��[����'��L����Q#�8����B�L�{�� \���þqa ���ۛN^0��*����i��k5����r2]J?�����6�����|� c߻G1?j��R����9�j� C]ӣ����4��7�y�>������ӌ�T��i�Q���3�����Sk�o����8cF�N�'-��@�d"��G}늖��üړ��[D(�S�~�A����1Ƽ�`�"��Fћ��8[�D���`�Ye���W� Pr?T���h\����h�6�x�I����/��譖aT���_-���p�b�.E$�d�1#O��T�IsZ��O`(1�T��6�!��˜hݹ�?��gIGD���QYG�{�اr�3Ŗ@�HQ=�h���x����������	��`�q��T5wPB�O���)�X�=�A���DK����r�	?H��{��>SVŔ˱0m�D��!��"ע��܂�a	n������fр��WX��*o��(#5X�Cx:�g�nRENO���� �<�p��?B��'�^g :ak*!�܄{O�G�һ:p�s-8���9���o�v<�oZ8zD��;�$"IC|܍����K�--����#9n�%H�2X|&�*�����;Cr��m��W�C׾�����ܑ�3�l� ���%�ޒ;AL����J!��@��@���ݶm��d�x���W��!v����{K��O��{Ч"�P���疃�C܎#I�`}�����d⧏o玟���?0��8��!��3n_�N���>0���P���,s���wCri`�/H��^�,.���Na,x�!�'�pt\L�R��0�� ���s�P���2,�9�-8�����D��!M,�g�W��`i��.�ߒ�'No|���g1AR��v5�nN�*�&ĵG����}б��4��
Vt�}���y/��\���c`�5~��kF
�
+<U�Z���;�|Q���W�4`º˧�_�2�M��W~u����+[ ���'�v!r�4����Mˍ*B��_��^�ƥ���c�g(�b�x��_k�h1m,���goc53V��*���Ye�J'�3x ���o"V��J�Q����t۪	P�X��w�<�F�߬�j)�:s�K�e+�Gb��F���n.�$Uj�'G��&��;�K��]d�y�w��Q��@��;X��1�H��,�e�n�ڸ ��#(V��{�wTB��U���@e�t!��.�c�m���QezށM}�	VQah>0�Uj�]%,I��$��vtW��`_���dٟW/v�.+��L�bps`����{�=/�Q�t�`���#�[��m�\K0}P�7n)&����<��G9�jňy��z�3DB�H��:3�����L0#X�E�1��!�X���-cЉ�+�Z�Ӌy��ޘ�٢���A�d��j��h^3/�[h���[}`ze�}�z�[�	��<�埮i\Hf��"�S���wW{��&�_/�0�<d�%� �6�ӷ<�3*%���Ԡ�)%��ƕXu��I��$WYiG<^�
	[[R�  �f�*Ҿ�s���&��z���Y^�%����Qb6t�Њ����������J�N��Ak�:�g�2����&�dג�����Y=��k�؞1��t��U�����D���a�<��!`��^{� fQOS���1!��MJ��Wm��J4��	�b���c&^��T'F0�P��ȋ�ٲ~��J 0��3�H�M���I��<�9��|k��]"��?����RO�@�T��}��{ŵ�/jI&�Y��� �����Xx-$$���8Ih:>�. j�	�P��}E)îNm�L�
n�u��P��3��f͐��X#�Qf,%�����E,���6�t��䝀L0��Z%��%oN��u��ƞ����AL��S��c�x5¥�5�z:O/Ć�Jz���^K"����*?�S,�Xc��kF�dHl����,9�g�VT��\9U��Ю�ߎ���n�)Π���ps�����l���Pr5%Τ��1��9��B��|8�/�(��86�+�����:re4d��oD=. \-�950,`�����)<��FxǙ�6�
f���w�����l������AecǢ����ķU�d��lE�$�9�ϯ��l���eE �$�k�xup���<=\�D;w�F�fp���G��I0�����/&��>�W�m���8� �> w�!�+t)1���L��_�J ���m�����O��Zg����vV��+�ͺHAI��in��]N Y��4��ڪ����':�{$�b�ʩ�$��J{�چ�x�=�5r0FM��n���A3\���n�׈Ϭ���̥��*����S2��J�`�����}@td�/��������j�.T�t��rR%9�/��j�QzY O�+mM��t�3���j,��։F�?KԩBvu���ښM��J�6۠�U��rBY����"�+�M B��IN1Td��+BX�oyO�V�
b:U������H�1�b�*����G��'��6�V!RALXMؽ��]L�^�j)�-�JUاL���f���%������$������3���]�G�P��H�
0���>�Bgo��*_��*&f���y�d$�yih�A=�R�Z(�5�O{�Xv��,Σ2�sE s�+�s�q"��[��B�BN5�Rwkq�%�6&L��E�҃pa�������ؿ��p���ݩ��Y�v�� �,9��)McSc�
+<�L%���t Bh��n�al�� ̹����P�öfY�7���_�V/q��H�ǉ�u^\/r]�MH�p�� :-3Q�U�蘻�����w�1>�QК�`_mR
�]���̦ҺM�G�+8�`�wg��x)6�hw�Rf�9�;�ο؄�k}��޲Uj��' ��q;mP�k�*6���)ɝ/�,1���U����?���'����x�VؐE���_��6�.C�h��~�8C���ɃM�BG;�5��j۶A��mp�-�'��Xu6}��1��ߺ�YCt�!�Raދ)�&��q����
��?�5_!��QBb�Z��n�Ǆ��`��/G3ޢ?u����O/ ��c~u�i��2�J��!��#9ɧ �q`T�Ժ�nL��	��XPQT[�?)�����%|6���C�
P��FլX;iͬ�q���h�"�_=@8�c`
	���Q|>̘^N?���x��Z<��\�����E�v���<��p{y��tD�F�	����M���q$�����hI��zf��Vke��Z��c�^�8:psb\�V��:�Tbbx�媶�ɟ������q�{ L}��c���	��D�4Jm��o˶���f^�]�)�y�YR�����a�N$D�WUjq�#V�$�Z�_w(�#~Vt��+��zȁ�[�� �?~��7A���w��m_���Dz��Y5ݭ${<����eK�k&�x(�Cޯ�x��`�Xu�n6����������SB�'�Jx;�I��R+�,�7� �2��!Ej��_ؚ�
WА��V�������8�+�[�质ٯ�ury��w�3����|���ǽ��%˜GZ)��@��́Kc�e)^5#�{���l�.��³�7�h4j���0c�ѹ}�&m�����Gh_Qct����8��4>9"�U�K�?V�h]6ԩڿ*2��`u�<Δ�U���k}��=�gù�9j+��I�1熭)ŊK�'o�ږ�ޚ^}�D!s��'��3�w�p�0]~�EC
����%Э$㰋+�ܷU�E�X�[RQ�+���y;���������l�q�K�G�Ŋ�A�X�xq�:jǕ��7I*ϡ�}�#��q���p+��T��?
�������6/��H���ȹG~����Ԓ��U�)���g���j|��#M�G���㞮�'A�}�h�T�]sh���1vB�R���S	��<65�V��ϖL�4�e��bw��a���f�ze��D�˒�'a7oy��G�p|�l���*��U�uZH�6CVF¾�C3�-��a=�R���A"���b@�Rס,O�f��v�H}�����z�|8h+k3�$5�4&�ૹ_��E��m��R-��YDm���N�ݙ��9�pk��sɫt����0���Δ$h�JZ��!g�0�d6>n�FW�U�e�a���uT&m�8�AP����oa5 �U�����UWg���d�\-�d���1��)���ծ']�7�����TmN�#[�Y>�[e�Or�8O�@�j�+����uOe�sv5���	(f�M����m�\F��CL�*�J���Z#QoSP�ѱ��{�۵�����X�����U��T�s~�f�IVHZc�<��4�[�t�>kX�&�,B�ȴk���n^3����+#}�r�e2���j�)���\Cr7�N ��:�2w�	�:���o��HD)
4���v��㦵9���>0�i��ڀ�A�N�*�^3?YOi��F���E;�WA�"��J�ݾ1�����p�OQ`���#UIm�g����R��nV2%
�L˭�2�����K�E����Ғ8?`RK �c�g��(��ri5P��X��"b�/<��~?����9��0F�,vO����o�JTF�r�!i*�i�=)ď0����d@�k���o��Q_|�R��%�E��ZK��*<ѿ̖�j3I2y~3�+�72����̕�� U��a�5���t@)����N)�w��#�����?-!�g�GV�����6��y�_
�2��ΊgG.��҅��/�kq�
��%z������6Ku���Z�D1���c����8�C��;���bb�f���fMC4�0�*7�s�}������L��HPn��9����|`�^�Y���!��M��H�x��*�1ʥ�֝���^��P�����/o~*˃G��	
���ۊ3��`�R �/�p>�o� �g8��HK͡-P{vz�[��'mY��
c�����ĸ�PXǪ��c�n�t�'F�qe:dF�HmI�S��
)^�:~�%�%pP�;��ؤ� ]���89�/��2�Nb�� @G�׺R���;
oP��?c�_�*��86z'���=�p�Mw�A���I�]eڲkT71��%�G~l[P�L-�/MҌ��qD��|�������JiRU�(s�]7đ\�@> �k��IB�'g�k����w6�rvi��4ʙ�Xf�Z��äp��h��/��� q*�|O�yBҩu�(���s�o��	���`��}\��E�f�����r���4��mb
�;b�_C��Z�ҒC�.}/b�4,�c�|�q��K� �ڵй5)��e�.���=l�6�=F^��*ע,cI���|���Z��ˈTQ
���B�&e�w�i�#w���~�@�ޱ��V��얮�М��yL@ܘf_A�gk⠻u���&9�4(DC%x��Q�ܰ��7]��cc!4�B�q�<�q��)
���'��(cSu1�&�H���v��D�	�4~���="��&=�����������ؙ�Zs��� ġ�mdQ�X_��-T^L���wt�i���7
��'�����͕H]fks��!Jȗ��P��Ps�QF�yuU��Io�[ɯH��-�D)�,�g����ɖ�>
:x�|x�A�V�Yf�;�5 p��e9����.�4�]|�j�r42����z�T����z�iv�
��8���,fyCع�1����Ϙ�Q �N��xL�ʘ�%��W�Q�s�MEj�L��BD�x�f��Eb������㟫?��=���=��_%+�/Fs}dl%Rzi]�$��N\(��s�)�R��<����zD% U���D��I�\M�"��2�~�3��z<E	cG>P�E�ܜ�֝����2:ε[7.%\����t�<��܉oCັ����O�{�u��.�crWO�F~����yy�X*��R(���˲a׸j��#X�b�;�k�I�C�<~�&U���@1�'��1�B
ч_�����i��3����M���b��vދ��%n����/)�)Y_y�?�c��Ȣ6���RP�de��I']�A�^EJ��_T^�0�s}�sҎ���0�١i^%�uӄ^�/E*(��.������/�3n�Y�>L&��h�-�����3��C{���p/s�Ӧ�x����>Z+ɣ��eU�.����.I�-��+�آ��Z�Tn��eB�"�A=O�9�8�=MA�� �5as݅�X[�h���E�理D�f�=���_��Rlֈb�d@M��z��L$�w��7��X�({D|\���`��ɺN?����yϲ�iZ>�L�bJh���E8���X6�㧻v��l��B烖�%h$+�Xr�iA�5��r��5�c�����"5����,*56�g����c���}�V��N�H���;� �68� �),Z��o� QG��&�i&�z���L\`Tt���`e{�z��@ׂ�sed� �q�Ys�������\I=��ܟ��F�0mr���0 �+W�U�.���W�vy�[�>�Rv����#B�I�E�v���}�(�w�뒢R�ż��K�uW�p���9\�E�c�t��"uH[����6�c\���BY�X)_hʙ���2�l�xU�@ t��sUs�)H�s]F��~
'�̎9+��#}��!Y6������j�W�Y
�r6x�UBa+u�V�E��u5�����&$B/� C2���̛$Î���Q�b��	��
K��x����h���*J?fY"3A��k���F���V�:��>{��'�Y�b`�� �P��J��C�o�TuP���9U�b���� R{��ޱ���E����&$�#�'p]p��;~�� ���H��')�k=��bD�������˔��Z��@f�jh�26�!!���!�u��ߵ�۔�����3�g9u$vʂY�Y
�Ș�, ߉���vw�.�:HM��ͭ���:��ң�=�C�%<W3_�ح����O!��Hen$q7@�I�u��lb~0Y�Gd��L���9&V�x#�K���T�����ma@D���z��Ē�x%� ꑘ��z�gm>O��x�/����t����R���|sX��f��L�o_�|�@h�a��c1�#��vC9��N}�=�4{����	>$�M�WP��c�.�gM�eX8r6���R�(r��R��F5|K�R��/�&��x����
"io..��h/��&f�T� �������p:�Ӏ��<����eH��y���4�l �S^�:+4�ۿF���0�$�g�������ÞK!%�o��Z@ї�%���MeP�HrH��y����!��:.��f����%�Y�ֹ4ގz2��C��;�Y�.�ĎЃ��1��!�;B�aƎ-��4�( �^H��:v��b	 �jB]��l0���F��oT#��b9��xF@���+7�B=�A�+�J��Q�m���g^�\i��lG}O$���|�3Se!�}�UC���2hq)������	O*[���~K���{(d6��
��Y���p=����i�Dͺ1�-�	S��-�X=��H3J!�Ձ�$I��7/7&G�h�����^-��>|�V�0��߿p{ʉ�$����_�0+�RW�ko/��9����.�7� �D���;8����i����pmw-=���(�;^>��詝��X�%��%��P�L����/!5�l�n_p��'�:my�:���ᾄ;�X��}�U"	P4F��̩�"�}����[5�"�`���u�������!�tw|�M���E��xC�9�4��HW}2jI�T7%�r���9�N9�*Rg��^����&�J���~&�Y���H5����V_4��h���3+�ta�Q�;y��)2KHJ��3�$o����^վ�R��?��M��@��@H�/p	T	�V|�	I*�ʰ������_Z��-uE��׃�������U?�ʦl\�1O����i��	@s���0�ݸ4��0|8����6��fא�h�)���q���{��J�k�]���Ը㧒):\�i`̄�}>�q<G.=��-R�����9��l095.ؤS6���H��菒Մ?�e}�">I�xO�����ەM��#�R� �żKPu�M��#��M�&�'��T�!l�^��Xf�zBeQ��S�;��O>��eL��a;����T�_Mi x��f�6�ߝ�D�ĕ�'f"$�[�Oyo��GT��:�CBi���T��d�3����On��{��d��>��f2��*�]�7:��SS0�W�(��謉�W!0r~ ��|��###Es;�ph=ÜWc;dl?���!�L7����9���k߯#�l�M�/%��1�4Sˁ��Cg?��q�9�]�Vz����
%�d ���0�.dǷ�\��N�����D ��7~� ���^�z8(9�F��I�����m]��HB/�V��)��ޘx�N���|h�=��~ŕ��֜�n��n�T��)hO�~��1���sap�kXE׮o��_�`�
I|8������A��~T�EVn�+�Е��=pY5ij���C�gNe�Q�@l��*B6� �Qs
�(Q�����W���I!nA���s��S�`���:�8���`ԯ�x��H�`Et<�e,B �礗������zR�@5=����A��D��
6�c�B\<������� �+��\���mM%����E�D�:kZ����S�g��]�xn\���3_��ϙ�C�}�W[[�!�u������(y_$���uZ`m/��z>��?U��8o�t�_=�'�3�B�_�ڡ�7r6:��;��~��9gO̸�cz��Ze���j������q��B��N�qi�O���7T<% cuo�d��G�.}��~+�+�G�J��aޮ�S`Xă��B@ /jI�L[/��kF��|���M"�ӄ�kH���P;|���g�h�!���b6� �W��Y�E�~�LL�zW��{镁���r�.fY�Pʹ:\��4�m�<J�
ىl���E�w���������E��vj��M�t�tF�NiMj���hBTח5��T�X;5�Jw����YAoѿ�,�M���j=wSE?��t���h�����%��p�K�}	~�����>>�]⭑�X�Q���T>��ʴ���x��He�դ�կ��/U;P�M�څ�����O���+����;��	�݅�ԝ,U�ͧ(�D||E�X�y�0+q���dA�;�ʕg���=��֗3��Akfcoy(���h������O����S�H�n�b����7�"�Dݗ;����>�5�z��T�,V�Ȓ�R2��%���5Z4NU����$�&l+x�HVaB������(�g����+���v�IP$yCq$�j�F�W5ݸ�̇��40�f�m�����^��E<�W�8�;W$����+���P�Rl�n�{])�'M�*Gj��B��K�}�wD�n˨}V1�N�uyEt�TM���j;1D��A�T��]J����D%�Ԕ�� 4wǢ�ٸ�
�qq�0���X�C	���,�	��F4�a��9,�|x�4Y���|�Cz���>�a"��#1�d)�u���c�_q��j�BM��\�r�+�����πa�'7ۣ}j���:����I�D���i�}k'�jy^cGP�{Sǅt&��L�zÁf�	榣_�^~w!�ֿG9�⽦�9�$��U��P�P�yUU�- Vx�@�S{��e��1���*�(��OD8����~6) \㜟|�4m���	n"�ǋ�%��t��~8�!_@Y�gr���v��M�*n��Q��@����seh4��́w*4�ըj���D��4v$�~�	%Ač�vCg����[���y2����l�1[� ,#�z���=?v��sP��y/K'�g�(�{�űE�yĩ��C�����Ň곲 (�V#3s;�Y���F���c��sq��&d+,	_{<���7�:�&���Y�PI��G��擦|��F�9�7'����{�� P��1��.��������m"Ia�y��>D������I�`3W����4��";����ơz�R�c.c�Jg��ZN�((�j�s�?L"u~kaf�9�X��GW���G������,�ln(%Q��=�p���O�@��8_Q0�C;�$3Ґʒ��F�]�c��ZS�5��˼�S��E.r�[pL�����Y!�����\���q��}�y����I���e���u�}�9I���At�*v5q�pr�$+P�w�	4m-Bヴj�;�U�(OF������f��Z&w��'Ofi� Mh:.2�,#�-#3vq�\�d��4��#���R!
�E?$�ƴ0�o��c�����օ��B��!4��tvTL⢏�i�����?+R2��9N�Lp�{��]@vm<��%8��,ϯ��]k�tL[��OE+������<q����vn��E��5|�RX]���V|�T��I�	�U��|;����R�ˎ
 J��+�3�s�]F~�p�����p@2�=���勇���aU�ʋ��~�9G�I,h�9��.50륽F��Gr�s�R�d��� �i 9d~��᪬����wS�ۿk�ߥe�R%�h���v�!�%p�Q�C�\���<f��H,6>a���H��&��P�tam�H���@�q^�;<��k��1N��I*ԡ�1fe[��q"`m{�@3�%f�Q�7�����~]S��ko�^@v,�R"	�Y�b�!3:^��{ª�S�S�0��R���;'��ym�_�&7\,"�t���K��Es�nfd��(K�c����m����V�LSU�I+&�q��kfr�;/[),bG���R$Ø�����ق�M�AJJ��M �a ����_{�6&���/��4��v`�h��a=�䷕�o����=�'��_��g�Ғ@�N""��#��aC��n���'�7W��ž��ÓD�"�rp� Y]�ƅK��3�I��4��w�`ĊZ�M�Mʗ�,i��O�}.��xL(2�%/P��$@=�.u>`<��W��w�����t�$j�����b����N��%��"5�j��4�x/Ն��yN" ��*pڲ�F����s���ġQ:�!��ﱩ��yaj�}�s�G8�g�D�w�P4��y�{�O�߾*�.#N
�0�mԹ��C7�)��P�u��F�0���K�(?vݹ���nܿ����� f��m�����-㏙O���_NH�� )�>�ݾ�@��������㢋?���1���?��7C���+H|��L��;�N�o,#(�
D�o�n{N}1"3M����
���v��m{�uC��m��f3�qT��?�j(�>�_)2�Xr�gc^�.���z��qr��¡,�F��_�G��	��BQ�blm��I�xf�˩���O��%-/������hp*Q@�{��K�T������ X���S�������_.��WP�R�h���DI�����P�G�A�F�~���.%���p���Gg������D��M8�C���F���U`R�d@��n�c��`�Fr�N�`9Faȩ烆A<����A_��;|>Z�¡�Xq2Y��#.��H��l�\����c�W;e���z��r�)%K���a�N������a��ts4E΃�W�\��*ݦK����D���~�;PD�6_�A/�pҙ��.�ҸhӴ�$r)zܛ�|
�swV�YK���N*�߶~���76�V��3FO����Y���,x<{`���*1V0d������=�b.��c�܀�P�Qu����\Ǔ�Y.!�WV�E��>��Ν�1��X��+��;5�ަ��V�jX}1�l�FU������K4�F/�B�Å�k%Z�k9q	�,g�������8G�}�7-ت����Ȣk�H覘�l�~�P(]C��]x������(��W��"��؀]=���M*,A-�|~8�XZNK���S肈��r�1�_��[>`L�̌�W��k+��Zt�Rj����X�7-��-\oo�)� ��aD ���s0���I�he�D<��}:e�T�*�TL�}��A��O8�F#G������ʿ2�H5l=���6�FנD<%0�������J�+� '��[�	��lJ/
��e�$�0�	�TV���uq%��Nf�=z�m��ȁ�7_E����hSUjA��Yk	v�0�?�ٟÔ�>�c{���K�|�}�	�P`TD���x/���M���v��V�e��_1ex�����������-�C����k�K��Le��r|�Ά7�/������|��
��\D�2����*:��s,A�:�4�r_�k��(Z�#��~�%���a6)ǾN�`����6]��W��U�c�/�I|����q�#t��s����_�;&�i�_K���f~��ЖA(2�K^��r�_\|�!��Ǳ��n �]�`��SH�U}�׼�.�7���ƪ\i*̩��De�ol
��WL��J��T����'��1o�A��%�1{�=��Aham�A����5ѯ�F�'����Ե�}6��6���=C�mO���h�~�*F�њ������Q�-�Q�2���@s���k޳6��a�c�B�˸-p}�}��G��[�p���@�����e5��+Y��?H���:�sd^��u�00��j�w'���GH�3�T������)I +���O�Z����A\5p��z�Fb`ń5P9��P�H0������\�s����`H�4�GȨ�����훢�s5˻C������V�%�Mo:Y�O{�(SFN`��fsr����O�UM��<�O����撢����5\n[�Q�3f)�?0�־�C���z��O��_�� wIi���OL�?~!��}�a%QC}� �G�$�&2=����� �xb�l47A,���4/�c/ �L1��'ĉ~R֍���J[�Pd��2X���}���aa���H�m���`6N0й��u(@����D̘`N`�Nhg�|d�OT[���0�=U�:I�jѤ���I�%�mTlx3��?C��
��f�ZX��p�!�KRe$�{���fx|�$���n����JE���7�v��Οi�%�m�+F0dz�׽Ϗ�;��5� ����@�\�[��.��fl!��A�P�-��C�^�׺�}��� �x�	���gιJR�o~��p���e��{����q���|cZ��D��E��xO≰׊m��-�K��(�+5oý��p��g��d ��@0�v�螵��y"���]_�B�d4 ���'D� ��^��QN���)�$�Z��񥎮UX�5��%N����} ڸ�����9�DG����:�/�
.p�l�+b�2��8��=[����J����F�;г�mk�Ij�>J�w����9P&��P�UM~Hd���	�+|�DU1tٞ�7�.����`x���#�=�E�1�u�I�,��_-1�}Ӛ���F�~�!�T���K�j%ߍخy�X�FӨߍ�N���=�B8:���X�Ue΃د�B
>ɲWOm̀�t�ꙫr0'�� 9�}D%#Pզ��v��;��@��Mr��zx<��%|��0yE&�W>��n~M��c;�O"�;��8�3�|�;F�ͼj��9{8�C�y����K�~j�;ƴ��[��<����~�&���Ӑ� �#�4�B"���R7c��>K�� L�)�	�l?��I:pѱ�j�Cc�U�?Q���P}E|m�/�5�W���}|�h_7DV"X�Y BN�A~���0-8yR��pv�s� K���6;9B�"␃=P<�h��f,[~��_ ��h��+�c/�xO��ݰo1��e �5>>�����R-糵vs�I;��i5S	�u�B�����{r�G���Ҳ��B80����_�����%���H��3��=���N�����������75}�6�_���W�������3ll=�gP|�\����)L/{Mw����,�� �~e��l}s������
z��=��TPN�R$�(�{�B����7	/�Us�2�G��5Dn$*�����.%m�-�$�T��<��D�sB�'PY���tQ��K�Н��Lm��3��[qC���c�/�nR;����U�$j"=�+	�f��Z٭�99,��'�1ؤ��f�A\�01nƢ���f0,�,# �ȁcE����<j\.�dP[�l�[��^����vʮS�-C�p����v�E�y.IL��|��}��@+����"B�n窍�P5x���/<)���Qg��4%�VH�����z�YȔ3�\���w*i{k�І�Ю�`��vZ[l2~�\�@�`'�M�����I@%��^+G�A���AA����a�$� Κ�Ff|Nb�cv�ɔ7U���E}�9���b.�C�^|A��xH���ڰk�[�w��T!�������*��"60;�	<���4����o���8Ӫ�X|e�ܸ����1a�k�}썧��F��nt��✡Lx��,���x������EZ�xګM��y�=A������k���-tnI������2���w2�,��έ�>�(�'����5�ڙ{H4Nu���~Y����P�͟��T���J��
ְJWk�RK ����.8֥���J�U�`�/TY(��e�θn��n3�|7��S`�+��v�ຒ��`�$��]�Ѕ�{Q���]0V�����L�m���r��jl���ō(&�59�%?�Xc��@����DB�]�j\��p*��+��^i�<�0��^��(7�	�e.�B��i�P�_�n��ê ��Po�xnǒ ��K��� ;�?H`Y[����3J�XZ?�{Y绻&:bY#;t�B�١}����4kaT-�Cj7�� ��B�Y0��nL��r%p��]�J�_�s	��S�	�ybkq��m���F��w���Q��8������.ᦣ�xF/�@��[��G�����	�;D��5׃]��}�	=�Lg0{�������3q�q�x[X͏���TCPl�����ơL�_h'P[������i��`�H�B� ��*�5�'��J%�D���ش�5j���j]�T�
~jbX+�l��G7�5ߦ��%=��x�~ ���R��4<:_��%�7�W?�h���$"F�%lѣQ�v	��ϊӢ��8+��E��0z\(��J��d��Yɍ�"8��`4��ǈ9Տٰ*Qؚ�8gϋcK�^�g��r`A��:�y W3�b�JFB����{���.�揟��{F�_ܭN�<	�3�={��Ӫ�X�m� z���w#t�9���|�S+9
�9�HӦ�{j�7O������wq�9a�
�MspCڣ���H���` 3Y'5>�}����̱/�aj�Q}�O�@�a&	F��n:"����L�"Tđ���g/aS�iqjڷ޲��u�y&�G���a�.YmB��b��A�XV��M�c�ZK.V�L��1�D��8[�/`}�6�z��˰�L�/�Z 4��k�hm�z�X.����ʴ��5��-��ҕ~��K���;R�.���uVB�I�
5S:�"KЫT��4�@�ԃ��3G��P&08�Ϟ���2�N��oCDz+e4�0��
N��ɸ�3^�V��Y)�EV�E%��t8��=|ݝ�Β3RG��%G17q��%��--p���ʉ������y�];E�K8J��d��t:)�K�6y{ɞR3�6Tf��d�)��������?�Uȱ#ԟH5��Iq;�1��w�OQ�a�hQ#]�N:"�KAO}�tڻ�M��q�G����jy��)�NWQ��ߐ�ۓ֗��T"�B]���֠D��E�N��Z1���L4���@�	n6��>d���M�1��u�V�C.�K�w�H�ao��z3�3��
�G����|G�����_n������,=c�c*�+�0}Xb��J�\��|�+fk�A���A�z�}T��R�!}^
\����=����%,�;��/.�y�#��X{Zօ�@%;bN�7�Ɔ;��R`�2lTZ{��:7�� {��>|l�����YO7bC��.������a1�"E���6�ࣼҲh�q�3 �eR��iY�w�H5�ﬅ�'�V�K��?�o!�#;O�>��$����U=����qN�N���A�_%<ZxK}GZ���o�Z(�@ݬی�<�K-D����5n����b�2�����E��1�Tq���"(�ɑ���9�:����j�'D�׺���y�x�u����1�� ��l�٩]]���W���ѕ3Z"�	�}���Fj�N��oXq�47G(y+?b_�{�����_��7��.��ՒW��	X��NJ��֖���)[
��C�Y"�Ww�?Zk�;FB����N�L���n�MdC@~����Y�[4k��
r�V��r<+j���_ L��5�s�D/#�+���f��S�M<T�.�4��Փ�	��E����}<�_�f�56�YGpN�NN��Ⓚ�Y]�����p�;pK_M��W�k�E)�����Gm�5�VU������-��p�&\Q�0t6�o����',m��I����qpS��ȗ��U��W���v�����f|�c� �,�����?�X�6���)gb���o��]!���e���e��L�;ӷ�:<UC��KK��j��Ո�X�n���C+T9g-�&2�36��ضTξ�8-��I"^�X�uY�^g���n׽�$�ὖ<�YE��c�p*����M4Ȟ��N�"tN+A�<�&-�#�t�Z�3��O�X�=���p�Z{�sw��%@
�DcFIv% Vu��jX���i
�H��Sç���P&V*`aw>�⤋�����6�F�fI׊����GEś	G��AJs��痂�ye�+�W`�YĨ�\�A���+����=���tP;դZH��ଂF�����	"�L��*([*�_{t	�\K�>�j���$ݩ�1��<���cy8ǡ�khG�<�$�j�I����8oۆ�cF��ޔ8�*|�w���o?��*��	Cэ��l�?����yp�Ɗ�:���ӗfί�2��<M���ѽ+��l��v�m^r4�3A�g#�Z���݁�s�WbYXۀWȲ��u�	-ؑZ�5,ޣ�h��c/՜�x�\ $U<�����Ҽ�^բ��E#@��X��+-ས�k��X�j&����$Q=i�ь����K�W}�,�9��8q�g$��A��Kڶ=>T�P5��8H�}�����>��X�7���&�$
����o�̖/H
S܍���4%.G�(}��uA;��.�ͶI�}��RA|Ps��=b�R�[Tz��2��kh��z+wy3���a�<K���$�H�VI2$����CT�>��Y�
���/�m9H����һ��[��z��HH�l��
��]V�]�^b����d�	�j�������2jM��-	�B�޼����,T`��Zj9ږ�`>;h�Dl�IZ��V�|�O)�Uq�,w��6 ?=T���������.&��bV�4	�N4�=
S�Z�>�bB�b�K����Y�<���r�q
r;g�5��O�TK��������p�Fs�vU��Yb�~9��Z·%�dO䓺���&�Fy(�/��8M�,�Z��J��Ҕ����>gb>6^��?�1��z�yx���~��.p'������A������;�20�+ۥ�𪐍i��\��U��F�(9�5�2q��p�z:�������#�,�~�-J����	��ۅ����6��_D�0��^�¾���h�h����Ij0�e�8^/M���`�Z0�k��lԳE��$�X�t ���h�,�'JJ��&�:ZɩA)ҦM��F�8���g������v~���sҩ���|�&������(����2C��-mֽSG:1L�]�,�O�T����F&W����Fȁ����B��e6�0���p�U�AΩ���>ұ$w�b�B��<�f��Τ��Z� �M5z�� `����W��ax����H�����l���6឵����ʾm�N@����\�d�$�Jf�j�Y5�U����>m����0=.��1`@q�玴��}پ�V�m�Ȯ�l �~%N_�i5�A���MİʹCZ*��߫�������6���0 �k.N��Qd09�}��-Kr����������`� $NxА1�6�� &.��I`خ}9��7�
��ًYGDI5�Гӡ��x�g�^���O{!�*~N RM�mr0��o���W֢��(��?�O�mv&���Ț�[��1Pq9)i�`&e;��	�öoQ��=�x[���K�M��L7T]��H\��vZ3��~��J�7�kة�Fz��6��:��4į�uz����;(�	&E�lp���~��@��C�y`�w\'7�[hG�$#؝
��,���:)n����9,E}7�[�&��-���iF�ſ��V�+:��v�:厚$:� �=��!ve:�$`�n�X���� ���X�ۢ��F�+c�B~��P��i�d�P��ċ<Q��-Ҩ���5����=l#���1�O�h[}@�Ao���%3_q�c��������=@gڛrN�;8	� ��du��XeE�]C��@�0Q"�Q�{ ,�+��"����I:]E�$%}(\PXN�cF�\k��Y��4g� �L��?�(>-�#�'�C*?�zĎ@�t�@r<�N+���V^����r��σSfOuR8���I��aR\�q/,w:7�����3s-+;����+n*�`[�n>7�s&��l9�x��3)�jGՍN�m)u*Vz8����{��4�:y=#/�;�"x>5�e�i��)����i
���Mu�N�L�Y�C�b�#����9�l���/��]J>�ϊ2r<�W�� �U珜6*�<I��r��U��l.�*���QU�3"b��hŕ�?��r*�`բ,�֓<n�;�)j�>h@#��r����	��a[dbg��-�#)3z���R�Z�x���E>l����wWv_��H�-1ʉF�t���ݺ�b"!���
d�@��}S���ρǫ;�S8��8{��5��N���U�c�܌]�Ԣao5�ܹ#Ș�Yj�?>a\����A.�/�ٯ`��g�+(ê��qf�]�?��ٲ	1�N�s���1�緱�Ղ6u�#�g0�`S��?�hːp�'O���楷p&n�;��.ls���_Q$�[Y;��I�G>&���6T�{����bR0���wU��H9�͏·e
�b+'rEҧ��d�W:h6���:��.����\�ʦ��xM����Ը�N�U���ܜ�9��&�I嵲��4=z��Q��X�U�L��{�}�8t+`��(�/e�)�B�?V��i���|3^R�Lؐ�<1t���>J���p�N*v*3%���r�_y��>�t���XRQ6��E�pخև�Q��x�?�V�yi��O��ؘ�$�b���W�6��4��c�B��L�`eb�w���9é�|g�Za;���"&�_ӯ�Sl*&�gP�����jDT�7d<4�Z!b�oZ<�lə�/�����KP !Z�M�6�Ï{rS��z�K'��P���ǷBp��	��п�LQf�9��$g�����c>��v�r�r�� ������ ����16l�P��r�AF��K��Tmĉ4GD��B���p3�I��}<�*1�!�{�~z̥�ܠ��~p�$�?u|ٌ�d(C�Wo�����e�0�C(�jk)�|����n�!�G|`v��ϓ"��c��l]A��Ywٜ�["��٤j�g�]�����c�#�j����	���@8�XYɺ�Tέ�&�7���ZT}�&�?r�lPbs����8�.ڮ?}�h��c��\���T��O��ɲ
�C\�h����֒G���|�!XUs�=p��3s]1��C_o `�o6E}[nM���0+1	}m�AԷ O�'��il��
�~){�K�Aз��p�$�U�/^��l6*���zn/s���|�ʻ;7��Pnr���аӺEZgu��]��G'.>�6*"�P���U�{��R3�zA��|��FR8��(B|��Yh�J��FG�o?YB�ɭ����!�C�ҏ�& <��^�@gq��6y�y�#�O�>��51B�^%a2Rr_���'d�y���n�0g��'5&�=E7r�i�K� ��Q���(���iE����o��&�rR���5�L1�..��E��h���'��B����P��zT�rj�=Ц<�k@�b|���#�Nʴ)��b�:	kJ�q�
��Vu]i������K��:U�뭮ь�9L��w��5x�,fC0"|2����f�p`�H��8�1*gn�����E8�,���(��P�7�� �8�x�]VZ�l�UK���aj��G�������0G�XN��3�
��lt̀�iG�u��������Y�vP:�����q������������C�U�����J���;Q��>� VDr�]$,�����EV�h�yd�K�I}e�����X��¦l��S�$�D��k��а��g����T���|-'<}�����V�֔����	:���)�뛚=�L,�X����]���֛ �ؕ���#<�ɩN���j�����_�H߶��R�����`AX+p$����rO�R�#���x�W���0Ydc���6d������X��2���)uk!�#_v�_h��1 ����$��bZ9������qì�ן�a@�P@V���Ԕ�9��W�*����Ϥ*r0@��C��t�eb���������<.d�_��P�Y[�Q�{�z�e�+���`Zi�.JlkL��z4���9-UJ�/za��v�ջ���Ĳ�1��5#¾\�,r�W#a��Wn��\d�I��8�.�N���>ß�Z�#�ƛ.s�6�L/�t)�����G)_TZ��i�>��~��`�Ҁ����[*�O@{�m<̞vu�<4�.���k�)�"|bQ��[�$q���j[�C0U��<���Q4@�W�q��� ��Y�E�|������4��=��X3c���/��1E���QE��M,�m6%^`rGV?��W%N#�ٔD:y�R�ʕ�X�3�x]����9�3�V��EQ�C'Y!����g�{�N.�*-OɫUB����["ε��t�g4'��~�K�b�*h-��/���w:,�ri��TӾ��_�m�_XcQV���ݭ9҉��n ��ߓ4��W1\�z;:.zԁg۞�����,YF�׽j1�aU��S`�[�BF�Ni��`8P��%�����5  c<�y{�'��o������5o{�R
��ˡy�kvy� ���@M��S��z�T���T�mA�c=h)����yAб{:��� ӭ�X�JW���,��mx�Z�M��mC �Q���x�/-X E�~�	S��II���q��&n����/���l�R��1�������"f�8�)3�J��}~B�}ڰ/6�N����&;s���������h[;m�GMaMe�� ��V6��*���j�3�����	M�j%4g�hZ=�y��a[zT���Q\{㳓"���^�;m. d���Š�Vy�����xp��C�@�B`q�1h(��;F!�S	+�O���P�G�#�L%LM��&��G�^x��J�|&ZNca��ڂ>l��v�t�/zBG1,X/�y�<���
)�W�2JX��<�����=9!K�h���X��$��TH�{d0E�If�+�W��UPp\2y�&P�]�]˾4��3������i8,�43�vy",�/�8�:eP`uBdg����C,�L�.^��u��CJ`fu2��3��-og�0���
a���\=7�꒢֬���ʅ��Z��B������/�WpS�L��.F��o�Ӗ��N�ߓ#�4� "�j���8Ҭb /t���ml��^ڶ�����{�U<r|8b�$��鳻�ǻ2�0�������eOV	����;?�b�cqT�꒣.�>����@t��D.�h��˝w��{2G��p��)�J+
�b���ܷ(yD��Ϋ�SA�����j ��EH�$:-U����B��*��X	�Ǿ�0���_�4����bZ&y����:23�!�1l:R����s��+
��w�k x2��H�3F`�Ycif�Z���C}J��ga!jf�IE�@Ӏ+��1�D�aF��x�H���J��'=e/��6I�xOQ�]#��@I_��r�]J�+4���ც�x�v�mZ`1�:|pl;p��CA��#�б"}�`^ �yӸGh���(�fz���obz)$~X�)����Թ�i����sE�����a���[[@�~�P&BZ��4��ۘ�����"<�|�m7�j�_r5{C�w��[ ��A~:�=�Me�����Rt�t���]΃��)���d
a�9��Q�]eH���B�[�9����+�)Z7s0bR��^�^x�0ʫu�8n�U�	���D'2Y����͌�Zv(�y4\XP\U۰`�U�0>pm�	<��ve����4����X�O_��g̅e�£�z�s[D����Q�%F�6�D��qԜ�x��L��[G�� >A�&PqH#?���z%���'������������^\�g)w���.�f���32�|��u��F��3O��m��?G�L;>��3����:O��$Nh
�8w%l�*ܰ(pQ�k4O��[/惓0��:�N:�"���
;O�qu�V2@	��x��$W�w�/z��)�%T�[�,C��K6�Ck����CvY��#/w;	
MƲ<��˯f��d��Vd��s�0������I;$�:���R��xj�z�~ᓍ���)΋�±�Xo�m'���iF_�8���v8�k!�9˂��|\$��xi	�h^#K3�JT�Yj�㶟s�B�S�N��2���xn¿AxW��E�Fzڱ\�����~�O���A��c	a׊g�~���6_`�j�<
ml�e���6���9��VZ7�I��ϋځI�ܸ���"U���ܭZW�x�60%K�R*��kC�=�t�&�,�xsK�>�Z7�:;[0C[@6�A�w;�~��� �=��)�@-�����vd��\0,d	f���͖��3T�G��X���->ly���6�^�JPfWrv��)�7W/�/JGm'*X���WPaY�����u���l���u�� ��pT�h��:�Pm���+i�g����i1���\<���ձ�hx���.�@6�SJ����C��&%WE�G����/~�IL�P�ň�����������uxuZW�U�f�GSy`8��>\H��`7�6��D�����=����܊�)�9���l=��"*��8���po���>��Ч�vom��u{��7����(�>���v�RC}}�������T�Hdą�|�r��{����BZ�.�:k(M���61�E���4Q�^�wB��sHH")7X)��g�I����ى6vT�g�P��{Jq�wg�FcI:U��_�~ͮl{�1�� m(_�T���e������Y#%��>�r�cx�� �a���D�Qs8Xh+����W���,�����9#�7�G2P���ė%W	y�~�OH�a��;��{e��rr���4ˣ��w�ʄ�
[�A�d3�8�k����4V^�WĢ��g)Z<Q���w�&���=]�`��NO�QA��*ɫR�ED��^�O�:qa�C�M��Dth���".����l��I�� �0�Y��n��v�ԕ���M�<.�<���o�q@MY����� [�ы��	T���%c[,�v��KM�
��l&oh�P;-��V���*�
���K��]�Xlyt��"ׁ�0���F��yO���Wp;�T�wS9��	�A#��e���[�O����2��*JYFD����ۼM�9��P�������>$�0f����2XMo�<����5Ҏ����k�1T�L%�_	� �S�9/yo�����ބ����t��74�[	� ���ޖPG�W$U��:�����]�X"���kғ��ftٺ���V~����:�R�Qc���g�݋u��؊�u�Œ=s��w7FȊ�D�	��'_9~�cŮ�0!��&�Q��⧵�.��fB��_li���5��L���%�8T(�����E׍�Ź�������Ʋ{ߏ���wŻ6� ����N�W��e�����\KL�eR� ����8>�*�Z���8�ڭ�ȁ8p��~z'�i�,��i�Y�����a���mae6�ʍ�;D�1
���Q������\J�> ����J�u@�;�ϻ�V7g��a��_>ڕ=�[�l?��\>��Sr3�s�O�NV��ŭ�=G����!-he�[KP�k�^2�{���t׾�Tg<��b���R�8t��32-��1!�z��w{�07]rX;���N���������)�h���)�����P|l⍥l�T��-=�%'�7?uɉ0�'d.���e�I�S��/䥿��u=G�4eI�6��?{%��c��΄M'4vqQ	�R�Kn�D���k�A��xU�������W�|𻅠\�m5�FݘR]T�VS�	��1�q�nn/����2O�〸D��m�4-��M?Ѻͦ�i����x>Mj��I_��~�3�:Ul�$C�.2{����Ur4h�7��?��[�˓`%\j�!U䐘j��n�D��a��W�Kt�C(1*LM���Iů8 ��kgfJ�g"�Y�ذe"y=��� �heY|QX �:�t��9�N���*�̾O�[�}�.bI��ءR}�������a��������z��.���/̓ʝ�@Q��r�%�[1OܦM8#��xi�	�RXY�7 Gk+�C���u��Y8�=�~�!�0 ������7G�K�/?�Tt�6[��9C�Ҵ
�q�]q����-M���rl�{j�e��>�
締\M{R3ؾF_�+�k�IZ@W������I�o��v�m�Y�������vmݰ�T����c9���`�)�I4,}r���8o�À6�Ha:�A�m�Z1H7.�4~�l���J[/m�g��T���s��#��p��������Oۡ}��~���m�=�ɼQ�V`	���e���c�獕���!�D0��@#\-LZnE��y��طQ�3u�w��HO����P)g��n�bU;�e��Y����i�܋2�Hw��m+J7kA��7����6�"��+��)1��,��ҳm��>�/f��?�Ҩ��K���U[ym�)Ώ������I���Yc�X�cb�$�k)$<�0x�&\`�k_|�91R��	z��i�2<N��i�U����)�Th{��?GNU�|\�u��F�jTG
�9��L����#�p�&O�.�z0i���k�	���7�kZ�U�%q\��t���j �}�+�v6%���m��������j�P%�Y��2 �S|k�N/����������K*����Z�0�S2�y�	���&�GVHX�\Q���������n@V+�y^b�Sn�y����y��F��/�3��5���.�~��.m��C�E9�Q�?OU�͑��0/��JǑ��U�����0!J����j�c�Ol~_r�?��,�ƅL�\9��ȧ*�M�� ���c�����l���f��$_T
�~�n=���@m���M�E�#�e�t͛���6ښ�%u�K�$�{0�9�T�i��J������¯xe�*�sw�����A��V0��h�J/n׊�J*�H�٩�}�b�n�oV`�XA�����[��5����?A��v�p�OwY¹�0j>��u#F���֫5��R,����C�0@T��y�x��c�&\��:p� ��NY�HZ�v�K%ay��-7}��%J�x.8_?
�(�.NqY�/�_m���|��^�|-"4�Mf=�c�!z3j�X�����Mh�d0f@�X[J�<��E����#�w�\p��P�l�z�tYmm�kNNXX����D �@��%���*'��cp|f���;�%U�n.z��~jj�����Ya��	�3��<��5��h>�9�C"����rv|z5�1I��WA:�02�W3w��c?����0]���>�˧*&>3}[�c�2�`$}P^�bt{��<�$�!��������+r=�dJ��f)�f�����no�8 4� �+iָh�[��� h�F�$�{	�%�ϴ����@P���}[��/��SzؤHj����N�wQr/v��n�����z��Ҽ((�lC��'a�!xz��fe��q�=v��X�{#�Qx��Z�J=d���#ɽŀ=�K��gU����xP@�?���ߧ=<���5!�P �\�sp$���z�����d��9�j�0o�s04H�D��� '���'�Nzaߗ'�ٞ�S���2J�?U��K�0%`��E�V��,Z#�|O�k�ju�Ѷz�����l�|]@@��PΦ�mp��/����úT�v;�s��Mb�ko����p�����Տ���cy���w���0X	�͔#�%T�[N�}�oFU�L�ݫ@�
�+ԟ��/΋�O�q�<���`y�X��(A��L`{ԚY[%�$W�Dl�JxY�y3*Ey,AK]�!/�x�nh�!���q�h9����j�,�����68x��50�fܕ�OUn��і׮_��U"��6˾2�WI�b8���ga�D��՛b݌ַۚ��c"��thԸ!����!t�+$�x3�;��U���+HS��ҋV�Q��ݑ����p���Nb�T�X<�IF�������u�+T*�F�*��C�g�9��P+�"<�Y}s���x��l��(ޕ��0H_ת�N��_���2��0B�T�B0�a�<Iz�cAV����!���|�ɲv�6���o\>2�I�	�w�_��G�/�5���|`����"��^��&=UЭ�[����y�w�REZa,K�9c:�k�@����&+#���b�J7-�j�:W"�m��T�	ΧQ�c2j� `"��(�j-��A�˧�/�i��W4�&��OC�C��S��=U~��7��͇�������y̨�əq\�uonY�6G�'��͟�P+�W��1J�)W�[_�t���۴-��z�z�q���rH4��8ȕ�x�.�gtB���WOR��� =�y��m1�[�6�)7:U�/����m��Ecg�E�K�ɰ�}�7b�����Lg[n��	��\N��9C7�#9Gߘ�rJ�l�a�<|�"��t�p��G��&U��O�
��u��J��O��%�Z���_`@(��|��1������T��v�,ˋ*YsH���%�4�Ч�O�=S���J�"�M��Z���j1�k��֠��}�]�����stN������\�p�a�p��0f!Y�?��0ib�sq�D-��/�hm	JP��EOq�r$b�M���e���zܚ`��^OG��iO��ug��w�<�:�_(�IfKK[�f��Ǯ�k:^{��y�	iMWh䖰��f�V�&g$��^%(�I�v�G8-Q����Z���cI�V���ؼ ��i|��-⍖�qDe�1S�&�R�E��9>`�6�{h�����ׄ��̄EU�sCb��q��'��+�]�u����|��`"p��,!�B���LE>�ęGom����9AB5���ʹ��guAj�.0=�tL��p�O���I/9�� �Gi�	:m��z�k��2��uX>̭�;\�һ���3r�t���pHw���Q�B<\��p����]2��Y��9R�Љ-<K�aQ��h6���_a���IA.eA�ϓC�9'���k�4@u��Ep�+��͂C~ЛV#��uz�^�'����g+�ÜpP76�~	�e^F��h�H#�ճ��o9���x5��S�R�����w��<&�L	�<�)}�Pi\�1
��K!�}ME�{�)м���z[�K��N�����o�K4�)�4!��t��|㑅��H!}���w�ɢ���LV��CC��#Vp���cd�p]-��Ɍ�"~u��VԮ(�����3���џ~!��;�$
��K�6����0�S���
ѭ�lR]s�/0E�¹�&�G�`0V�a@��90!~�7
#�GA�Ԥw��Bȝ�&�����8�a~EZ�� �#�yc��U�KPpL�����l���_n3�����CD�ܣ㥾BO��x����
{����C�_5ؔ�|�N�8���=���hF�RsތX���}#\ʛ���yk[V˩�5���D/���^���Y�0h�jȦ�!��iFθ�< �UUd��ٴ����	�l�ʹG�5���XU��ф�b"ߔ:����v|��Ao����C�\KR<E�WRjTb̑�ON��ƶF�g:*QT��=�����d+C�rT��1��|js'¡���KW�i�����{'G�%�Ap�os�)�y��5����A�!r0���/�[C �}���)���2��B�>�m3�S��LX��-g2�|��~�;	E���~�)4��1-��wh�Aԟ�����-�ƙ�ƨW�
���z� �����
�	�j��ލh"���4-���K�z��+�ˈN��RuC����Zy|�K���gm����s
�q�<��*K�n��&/�~BY��3������x!v�k'_Ы�=�K�W02(u�]<�I0���02��y�̐�U8��C4'���y4�:r�����>81`�����K�������f�����|���ާ�0j�R��T�m�=�{��4�h�5nuI�V�7H�޼�p2��8 R)�SD���8�=޼���50��m�[|���f��( "Н�2�޺1{M'�P�*0��R�;3lGg'�fU٠��wnP�¶:�N���W��!#�Ϗ�Ze,�Z��2 <V����|C�=�� z�!ވ�#�	s\s@�+ѣq1�2ܘ�P��RX&ޮ]�*�/�-䣻����fe��m
�tz�;�E�pR�s�d�^W�������������a�@�Ň W���
�L��zPF�	f����� "_�Of�e�r4x\>ɏoţӴ,}��U�H8h�lNt��vA�\��[N��W�5ɶ/U!���5C���u�`���i=[��I؜[���p���5�g�/��=I!)�Ý�ٟdψ�陸��ڷDÅ{瘣\*�w���3��y�Q�O�F�v�zGzN� |HsӠ��������KJGM��7}��j��_�,�m���E��dJ�25�,~�5�
5���G��SL��c;P�aϯ�J�䳝�%/j�����������6� 9�.#IH��6��ޡ���פ�\5���@i�KR��P�9�����'�C,�gz���6�.a���ur��0퉣�#��i��6�Jܨh���h���i ���^�Z�F��T�Hh���I�ɿ�H�-�b�tB�TՆ��_��]��S�����mvέ�r��1I{ �nB�"+y1fokh��S�O�Ӿ!�K������p�Q�U%��viNiAO���T���Hk���S��ؙ��:�����Zs0���'��o4 �Yn�	w��P��p 9�g������7�4�nDڠ v�8�E�������R����7(̮�0���HȜ�Ȇ�"֥V��V1�A�Ņ<����"�]m1V��,N�U�ۡ�����ͱf���w�c�N�~FӬ!��3l���z�(�>EK�Hw0�`�m�����|L�l���q��~̑u5����(�f%l�Ml��^z)�_P�ROF�,;���	O���8U"��f|�K��Af�_3����Ż�ב;y霏�!7ܝ$��E6��_�e��,N�I�\_��ް)G]��[��\,�=ca4�k�y��2_�[��>�,i��ta�Ŷ4p
0a+gM��A�[���sByԉ�<�'\dt;zP �V��KS��5� ��]�	z�fdx.G�TEO|�X�R��P���@�]esVkX������ig���i19r�� ���x�NB�%PF	IӰolU���������{��q��[��� El����L�<�A��a�tA��?"�~�����������i(	ɬo� -9��2�pr�=,L���� Fw�<��5����fmC]m6{ĺ�k�ie�+�F�.�̳(J3�c�M85,
���)�H5=R�MsL��_��
dq�>&8�G�O���[�%�ڲ$�<$�+�ʖ�hj�����)����x���"�&8m�;;Q�Z�@��ͥ�2տme�L�w��`������Z¯���K�<ʓdF���ح��"�`�A�kz���D�yϹC/���.d�Q�>����c�%�\g�� e��$�� �18��i-���"Id.��/�ZWI;��"�Qa��n<0�+*� ��|\�󗦑��3][4�U�C8C�~T#�����?)���a{���Rb�R�f��J�s�V���jrDC` �+����p*����ӈ�\
�I�9�j� �1h���g.�T9�:ph��T����"� xJ���wڢ��O���2�.�&����GP��,f�ͧd���*fk������@�����]���hD�7������R��~e�	0v&ǰ�PH�Z�p�[���1eD�W2|,��+�x:9�^�	
X�1t�1\�R	R�(�O�Gja�v�h���ٳwәN��
��/��MQ��]@��ᱽ�t�JRjE�C�(1�8�a�Ͳ��i��6y˵����	2wsʛ���.Mݑ�o&�l��N9YŐ��������?=uJ��)mJF�X�'���)�NJk�/":���i̞ʥ�bJ-���U��*.�Nk��+�v�u	�JY����?5������gA����wQz�t���(��LU��DuW�X��@!��"�XR��ѡ�mD9����O�� K����T�.RS��2*��������l��/�דl��r�"Mn��4R���R-~��0u�1S߸,�B��C�$��f?��#�����X`h����s4휲��x1�n����aӏ����U�M�?���4S�8���N�k�kG��=#�E�4�؞�hp񐓭޷�v��2;] �����ߙn��PS�+���rb&��t������9R�o��3�p@a�����FG��%���=FD�0\�h�6-[�`e������Y��7�j��GҰc���Z���l��A6����HULz?(3~����µU6��W��C��2��G�$B� ם���F(=���0��� ��Nϫ����1c,-W�X�zj\1��9I��oT�?"�`��3�}u�����4�&��=��w�R(T��P�qY'g� ����*w��nW�5��	.�07��&1��F��׊��pa��2��}c�-���&'_-���O�)���O_J��A��6=��竬Ʌn��`���/e�]M )a����핯j���F�Q����%��];��tT,ڟ]�f����_���X-z�瑰���3]g}���j��l*W?�q�w��:��Q8Ӓ>=��5���]Cs<W��K�u(�֠�̜֫�鄒ka7 �}�P�������9�^Ue@�ys�X��T_���D�CE�X��W�k\ճ��K�x��t,�8G�`��E��޷�wGJ��N{b��zOm�f�ڡ�g]:�@������Mʶ������s�m ?����,��C�n'jbX�p=pI�č� �� ��>�S
Vio
�l���qa��9��Q�]�bst�S�NA�_�[��F#��{�)���2����2Q%��x�	�����>�w��A�c�ᰶ-��h��RB�2�>�~�tB���j�v��a�耂�گ��Vs/qs�4c��MaLݝ��P3���M�S�sH�XL�4�cp͔�-&�lx���W�w!{��Jz���չ����|�IIe�bu�ƝF?�^F�c[E	kX]T7g�Ke�1G�-"�pe�Ȕ>�U�A���3��.�!�����Wl�?�-�U�ɘ����e�X	�L/�V@�8G�^������Ơr-4������'�75o�Uʍ��Λ�8��? +���y{��:�z�5N��4C,jv����+�Y%�D�B�+�>�2���6:�k��x��'�&Ƃ�.L�ӵ"����R۵@�<��<h�1�����́��xچ��G��}Ol��&iB�)<��c���K����"�~jĻ"�S-A$�'"���<��L���~[�� Y��-�+�gK�Z`�j���U�v�xp�z\��TI�<{�Le�+��/q����7�q�r57C���ߘ�E���ę�5�Ưٹ�ǈe��bW�Z�ɸX�*��ھ��O�y���=�H[�m\�o-"-����������F+����D�p
|����Vyi63R����c���&�;>|���3�{>c&Z+�	�Htcu�S���i��^�7��� ����T��c[;�z��;xr��wr g�9�S��5uv�~IR��O�3����m�:Hn��,�$��L�y�%r��D��Dh����;� xǟN/�~�G��|x��$����97�Wg^�-��Q���|a����"�Sk���)�^�8ۓR��!3nX��DrlJF������@Ѫ!U�@�B��1�sn6�c9�	?Z�T:�����DbD�Y1�;O|zb�J�âc�D�N���0at�L��ۈ�$������؏�T"El?�~�*ᢕ�5Q�UT�ى��A��[U�?�����rQ�v�v���H��+��י�*��`�&��$�F�6��P7r}�����'�P��T��쀜x���
��<�?�l�YY�zI	� 2�6!���fG�,H!&�-6����Ό�I5U~FM�Y�o�E������	�r5�@�\��2�O���Ԑv�s�G�����h_�B�-b��ԥ�o5��D$)��!����� [#�jۿ;��m�2�G��7��"� �U�T=��Ƥ+��jO��A7��+���e3A(b:""����O��jK��)�U���(�W��]OR��bD�?��
Ί�V�Ec,P�4����m�� Nh�YDJ�A!{VnTg<��t��1?��f�-������'�r�SA#z���¡@,\%�
�  �!� ͑ f��x{2�]�#'�>�x.�5w�����#���z�~(qi�^�M�|�m���T�\#�~���9�����pc��;)� &�=4uD3`���:�cB����j�n�@R�
��G?lL&��vG�������q��N!Lzz+��#'w��{(_�+��I�H^�X ����.	�y̑?��Vbܥd� �s���$y�Ra��Np�F�����ҙ�W�aѩi��5F��.Z��®r����#�A��nBC��]98��~���o�;�Q5���v�m,�.�
kY'�s��c���1b��)r�����{���v�(aJ:A}�]�>���βH�Gܲ4��a��F���B����?X	�M���M҅?ꬱ���@b���m��cb�2�Q�>���/ʗ�eL����r���4�q� �fgk[�
����1&\����u��ܽLS��镠��;��0�O�q�a>h�t���N%�(pb{�����ַ'EX�Z�pe��s���	�h-����178���ϳ|��^EL��I7�(G��"F3�Bė����	ty�����,���E��c>��NCHX��>�ۊ��/�t�q d�o����O�)}A��'��ۜ�a�g:Q��s�'U�<�居K�Ղ��K�@�g�g��S���!�N���NW�A>&�%W������i
�{Dj	�)�l�\[������o�`�Zl��*��RC�x�ox�^�kT�q��l�f �D�S�4Y��s��|�H��j�;��/ޅ���6W)m� ��Sc��������L�jL�.J������'7�s���2�0g�q�]J��Z_^����W�j�c��tBl���l�mP����COS2qߋTY��������@������6�k�*9'���F� ���m�` u6s���@g"�2+���ʈ�D+��%�҂�
�!:h9��ΞM���l�>��$�'6H�M�5AuU�P
zY���V,��8:mTD�!�Fx��h����O�Ҷ_�����#ƽ���u�$�Br��j�e�`S���{ȉXF�s5P���gu�r�0~�+`0__Z]�CT�'~D�㯦�:4l�%&��=
�O�X�����h�٫p�P�)=0�P��-|��́��eHo;*
[���?�g��얥�u�x���ܺS���։U�+���H䀹)"u$v����]����Jd��I�ř*��W�'�'�֡��o>+��\�"z������x��)3�� \��u�G�-я]b���m|��xc3�F	�1-_t�Z��2.��S~o�,���2�K k�ilh>���p�����?E�Pxj�T�1�,�,E��(^��6@�f���db��5�4�"�� <"Rn��ddyL:ȅ^�r'�7A�JżBw���P��)�2� ��۬Đ Fh$	��ı����N�ffXU��7r�h�S<'���z-YX��k���:�J��"z԰�@�{���[��
�t��K�v��i?@�Ҡ� ��^�-3-ݣYD4���|�����x��!��X�$���V�ϡIe0<F��,7� &��	����?��CƄۧ��r��:����������3�",��i�)2��>��q	��W���8���S�g�����ΐ{Cx�Z$�Tg�x����Z��5�Ə��ZX�T��0��r��iP7b�ʇ�c<�S��Bu�4�6�F�ҙ-��ݖ�Z�FvS�x��ڥc�T���i�
J�C dԬf<��� �h�qD(�����Jf� )T^[\%eaұ��ă�O�7��/�$g*Lf�j��=���}���Ӑ�kҿ̘QݷN��𵴌��;�5��0��h�ov��ۼ{h��l��	�x��=!n[Õ9��s	O����%�Z���y�%ް�<��>cX|_n�;�u���l/��>_ɚ��y�/�$��Pbq��ռ���;2~W��3ׯ �:�%@�(OY��HS��g�9�J�U�����gV5p�-�2Lf�+y�m�^��ԑ�ӈiv����P^��|��=�VH:׌<�N���N������d0�ElZ���S�ܟː2�6븏j�-;�C�l	�U�X>�(~��zwk.�����=uq� �d�`Mn�E�n�=:�S5�)�������� Ա��txc�h0�_V�f4+�=�4�dlJ��������񈔾�
���Ѥ�E��g��$�.d����C���Ǫ3R���Y�\��skU��U����-����ro��KW�:k��՘-[��Z*����EУ��=�[(3�9d�f�{���<�Ż�Q��d�i*���?�U� �CȄ�9��BX/��x��P��K`��bg��
�j����!�?��M��I��*��C���DRvZڶ����N��/���PO2 ����D�}t��r"Ɲ��Rːֲ�#(b��+��4c穎���bc��s5�W�6��G9c�s���V��������Y8\���4#Ti��[��Ìf�#ƞ��&�¸y"^���\�}�>7X_P�w�ēf�#9�dР{�O6Bǅ�Yd~���iQ�Zy�G���W�������@3ܙ��x
��`���#��·�VO ��̺�N�{�8]���O��1RoǿTMs��E�{��Ss��X2����viɅ�(#�;s泀�0� ��gix�����!zZ�::g8�,�B�5#=U�itq"�ҧ���3��Gč�baH9�c��P�q�i{�Yê�$M�'d����M�& ������>�;���2��FW��{?I����Ӹf u�B�E�^��a��Of�*0<��ɷ3�6�[�t���[�P�栨��8�*X��g�ɔ��T��	#=�4 ^�}Z�9��-���+�;�Jd2���@�m�|�����kP���(���%U�AXI��8�ٴ�#-�5j�A���)��c���CE����q�����ѻ�(5�Ђ'F�:������� ��}���I5���`�N���������婑P���ʌح�C��AP�ec���~���#]�S	S�f�l��^\gĹ,�G�����Q��������8~�F٤!hD��]�y���,o[/)�5��Y��
�tU�|�;�|�N���ZG�h�T������|���.�3t��`v@�9�pP�*9MoT+��I�m!$mؤld�ߞJ�ء��ߒ]�)�v���V��rZ�H��o���ʄ48|��b�ʞ�nZ��#�����;���X �6kkO��Js*��J�"�	&�j]fHт&�Mƒ]럥)� ����reL��C�BQ���*�6�]�W���!6^Y�U��<�VDT�PY�Z?��oA�xɷ�Ǜk~B͒�k���������V��*���i.B�.���7u]���CR�V���iQc*\�CiV.h5%ބU� �/�ϛ���m]v�������.��Iz��fH��]^�G�׺�5f<�nW�����.U�抴ə6�$��4��^<����y>f�jt��]^��8��ؗ�;��3��>I��+7H�zP�}Hl�P	7h����=��\�f���b�֒A'T>*B�4$����[@������+W^<����&6�|t�)�`�)a%�>���q�9y�BQ~򷴢����6��d�������8Y�U�S���ê�l�BqD�;�*6^��{���YX�3)G���Q����e�h�iMn B�zz�E�G'���	������Q�F�w�򤕻4�"�o��1Jj߁�y���;$�D��ٕ�ĭ�X5I{�.��������\c�$NlWyC�["{Y��P'�u��u*�Iܮ��k1��Ch�\�܁!���y��T$^{
y�f%=x�)fjG�/���N�4�aɁ
q=�2��0q����,C=�Hg
`�Ц�"��a��fo7ǄTj���֯[O�v��l����@9��f;���Z����Š�Qx��>���$��~�e�*$i���Ls�瓺��r櫘Ǳz	[(v@~AA�7�>��(}��^Ӓ��9M��~�x��T�t/�X6x0�R�~�l8��LU�v�u/q�� )�X*�3SGZ��UaY�u��;.��fۤ�N;6�AWq�����Oڀ��%�kh�'�!������<=scE�ؾe���i͸�<�w���p<l�����"(�3M���GW������̊E�[n�[X:���O���GJ�zG~��H?HQDY�) uc�E���d�F�Ľ�.?�X�9c��wӋ����}��=��<�n�}��ʴ&�X�_�[�fo��^��|rr)7�L����?�Z���}\i�4C��F���-�!��.[ɼ�w ~���7<dk�F=��SA+a.4 �ҝ��f�I�	��]�w��	���C��$A�Z{U/���*��_jE�l�����z3W4[���2[]���2�H��k�G0�����_\)f~:D*�v��n����uS�C��"y.����n5C9���䖤ST�of`�H�M�@x�]M�y�e�,�.m.�i�i��$Dy"�Y݁�V�Y,S����"sr�*g6Ka9��Q[�4�� R�i_}�F��0_@+CX���{J��6lm�7f�B�y�FX"q�,h�+沬c&,p蕇l|�ֶ��+�p��@FO?��;�ԥ�/�������J�wg���R��NZԒ�k5�c�JЮ5v�1�!�On��C�v�28�&��Y=%3��{���Yu�H���W|}�#d�G�<��!-X�.��'A���5�&���Rg�vw�m�
=�ɷ�� �z8i����t��j�J���-�����\�j4��'��S�J�J#�tin�X��5�F��m��M��Q��5ܚf�4*���\n�%+���M�܋�&�.��,�K�q4V~�{5�E�S� ���`�k�6c��v-����Tp�s�i�b��ϓ���J��L����,���H�Bgw�3W�%�=�nƜ]&�
��U"��;z 3f�L��iV�����/"_�,�@R�"��z=�,���е?=�n!��i��Zp���?&���m�mG�C/97.�b�T!�����r�3��EJ%[�*����f���Й4dFJF^�m-�$����/� �e�kW	���	�.��Ka����/�d_�u����s
5���;� �a������%����
��Q��oha�:�M�:�w���F�桫��,�BKW���2<���D|+��x�Q��G�6[]�l��|v�C@���汀�6褹ȑ��q�,�3�Ì�ve󄇥��Dg��]D�rL�I���s���tm�U)9�����ؔ�t��G�<�^4��{A8���숛i_N�l���lNZ:g��C�2�y��:�w'��T���]ǄHz#uC;7���Qي���W����.Q�M�:z2�u�����;����W>���a$�b����FYP�M};��M��N�K�æ	���D�';A�%Q@K�.�


{d�K��@����~sq;�fbP��s�N��.�8eTt�a����d����%t-Mia}T���������d��Ŷ�%ő�|�fj�mY���o�]p����a;����B,S8�d�����p��l�6�X��̟"h y(i�^�4�����2�|K���1$����!o9��~���s��o[%[�5�{̿�D&s���+Ԭ�{��bZ4#��IM�}��܍�_�L\IW��ڿp^[��D�[��d'Btux�L�Pa���s��o� :�E�5�*Se*9���@g �d��=bM��;jlȮ������>Q	m��K����7y�� 
�A�"K&�uy��~�I���j�CvĿ���|a��g=S�nA���f�Dz�ٓ-�RJ4�҆h��F���2ЈS��?X�|���
��ʵ��$;1�0g0%�V�05B��u���y�d�OXey�1�l+�/�}F�3#�������Ҕd������P�Iؒ�yH�;�LڴN
�Ŭ������IHJYg1��d?=�Y��2�>*�Uc{�E] aI+�5	�c5��t�=�\���� WѺ���`R��p%՗��h -���.%�c��G؋� �\a�Vr4��uu!�k/N��k�ӫ�b�sE���h8���5k9K���҄'P�c�c^��w��/.�c���`W��=_ ������@��G]!$0_=��N"�:��)>��/��l#� ]��%�rh�2��B��8�J{Q�Hc�}fΰ!��ު� �S�9���<UB��uBgD��B2ˮ��6�,���|�y%t��DG�oe��s����<�C@Xy��0��
�t��Bh>�o�F`��f���T�K�O���7^�k��u(>(�sp�I�����6��x�-���iݺ�Iۡ�`N���	��ކ��4`%Juh���o�S�0:�;��)���O7�����%$8�D�Xcɾ�Uܮ����Z��U{6�3�1����Ù���QZ���Efy�H8�����u'si
������E��e�F�'�o��}R#.J�?M�-w[L�v3ݑ�2:/��9����?��lHn,��	��q��0Yxr��Y�?���k�oZ�{r�}��3��ax���1݈�6�C�<�P溟����~�Ob�ϐ��1�M����B3�ʇ��m�=��[���tO[ze�X)y��BL�,�7��@7��lt�x��W������w�;�o�����SCC�C�*�('!2;�'����2j"\�M���gC�ZO,[E{�r~l�ܴ@=�]����G�ݍ�7 x�oJ�����������I<��4���Y^����>>�Ãq�ɒ/)�^�v��xY��t���2BKL+UFH���dC�i��!���΍LV]��冪�k3D�:������Ov煋xB�����SL�e�ZC�=TĆÑ�����x�j�~����~ǻ�N���/v��5���Qs�V}.��
47@ɶr	���wx�S=i~N��Д��|�Jߍ��]���%���޳�U�wy/.�Н!�E�m���bT�Dju^�l�y@�ܽUS����2��F.tŖ��JO�dA,x������X���^!X~=�X���L;�y�\��&}���+!䝱K���1B�N!����t�t#�giO��ԅ��Uk@G��a56�%%{����M�j{�'�Ŵ)��i����U�@�c)�+�c��j^�����%��u�4���̏T�2�M�w/��Ƌ�כzv��сݞ�c�����V�m�d�"~��S��<�X���8Hi^��?C�S.%����������-�䍿�+�����S���T�.ul&4~8��Azq�E��Fѡ�/HzY�}��� ��G�WqYv�|�rIE\�`�!b1�bH`��#5$�����{w´��ڒ!�T&��x0�`<:o��� 
�r��S�=��F��{�z��lգ�QP�M�,h�A��+[&��@[���p��HF�Nb�pȩq��/��Lc���a�<^�-�����T�;�R��h�����J��v�Q�w6k������F������&�1q_�T>+ ��<�����'Y珓w%�p�������L�]�$�������5�l�Y�X<�e<F�3԰�Z�{X�;
*�	��>�Ű���>���]�%E>1�����Jw�ze�N'pjײk���*�)V1RΤ�y�[��C�������+�#��:���G6��oy ��P����ѿK���0�q��&���1�q�Pd�ޘK�Ӂ�>��+�q^5�4��"�ζ��hUY�G�ޣ��{;c��	�`���*��<�&猁�o^ȣ�ը u���A4B���'��%�޼��7rR'PNI�<s4
���2�3��9��_�|�F�c+��5%�I�@���j(V�� J���4 ��t:�P1,���ҡ� 7�g�ƒ�˺c��$G?���t.A��%�ZR#�U��k�²��E#���v���T��� �D�8�ݧ!M���Pgۅ���?�V���nı%L/��p�S+`�ǆv��D���0�򠖖���2�n����Ƹi�[i=�q�!:LoY2f=�,+���?�*W���ʶeJێ�rL&�g����F����ꉘH��9��۟� �Z4�6�'��vΧ_}D����3|�C�o�9q��r��6�˼u�[�-w�uA����*n��G�~�6'	0���З;�A���=�&W�|��k��5�c�a�NSJ��b���8H�t�W!)�n�M�2��ܺ�޻q�]��n=��c�,����!&�פ����*X��Pg��쇞�T��Wp�a�ˑR��I3Ĺ�qL��$K����;6���Q9�;�H8><�C�K�	L�<Z�@� !����p����e����]��g�F�-m�H)AI��(�Y��٨kj����Ix�lD���E��@���M�&$����_$�hC(p�3�up�8H>c�ɍ�Nq+��Mr��Sr�h�KW����2��^�T(���#�f�e�8��qsBE�f���rDS�2�s'Y��+O��J���$��b+s���A�/�SW��=�:�:��x��$�F��sk@k3��^@Ͻ�x��cgs����j�d�W�D�
�����|imj3�e�n�n=G�M͐@��Z۹���4�6ԐNA� ���m���1�D�CdI�A�ldS0=p��t�J���>��������ɯ���sa�^�����<(Y�C$��w���c0B�#��xB�*^C��>��/?#�}�>����U�!�*���{�uE[:�����`��\�	�
��N"�c�$���9 �����o+�7=��!K��#��gn��n,��]�{���|�9�J5�_RQ�n���_-��(x\��i���� ��
��.ٿ��������FB�;��b^s"��d�!�K'ġ�
^`'��r.DА�Z��9\(����� ����L|�*%ז(Ec���'�����*H�X�w���
������5,	Ь�1 �F�F��#��.������9�pOI���FœEV��E����d�M:����!�6�+#�XX��FQ
��Ϡ!�BbMP�Dd:.�'�h-�XL�SwQ�o���U'˾;�}+{q��P@��g��>+}�x͢�i��"����7/��;���ѣW�� ���ME%I������	��.s����7���g�)���L	�#�`Y�8':yI���U�{.��2J�	��G�z�/��Kp���`ݷUW�p���*u�Bk�J��	b7�7{A��H�=�ĺ�uۇۖ�������� ��{���q�U��)�糝�2�x����6&z��%��9�[�2��b�2�z�ڶ���c--M�<|2SP��^��*[V��jx���À�}��ks��q��0���5.�ń���߮c�_`�U�Tک����j9k�/]Znu�wQW!D�<����"�����F�)Al��Ժ�$!Mi@����D���^�95潱R�b�+y�g�b�ݱ���X�t��UaF�� &���U�ʸ_�1d��{���	z�.�>��x7 �P17������M�Hq��]��Wb�R��> ��.��)ھ����W,�@y����7�A��<&S�2!�����8^�녉��P����(�k1�7I�j$|���'Q��ŖRAA�N	y����hPoʻ�j4�F4��S���U"��.�k=�����lc��n�c�SvZ�m=0��(4���CQ���B�!6�<�VmZ5�����0v����U	�n�՗�}�I��Բ"S�3�Ȫ�o���_1X!,.<C>��1c�ztY =y(b�W�/���[4�Ѳv3Iǵ�;��'�:�W��˱&[��}��7#bU������N`v�*�j�<�;|�M��pI�G�?6�]7Z��l<\�,�l�����!,S�*���~o�ԏ��R'7����L���j���aE���c�w���L	��#E��9DW-+#A�q�R���(|�Iٺ~6�>�% ��}�˗�%?�g�nF�o 4m�!H�n��a��N��uT�(Q�@���9�-v�)�mh���U���悰����4[пP(4H!�1�E�P�w��r�%q�&ayV��`��g$x�1?�N���+���4)}�̎�ҝx34+����a��� ݤML��D�JU��� �
���p�j=:��r��}��)>|�^�T���+&;K%�%4����W'��q.�hfP;t&�_\@tf�n���>f������e}O����"��~�O�.�J����V<hj�ʗ�'z�l�'-��xd�O6F� ���s��F�1���ڥQ/�5Y���x:"7��
w� �n�N琗����":#����=9�0T��D�"�!��`�����u1�]"�d#�[�"Fp���!��sb�(��������爸o�1�R�A0�_/v|�U�����C���m��|:w���sQ,�K�FY�"��\�<L	Ax��� �#�����  ��$�FAЪ�)Sg?JV�a=�q�pU���&�O�[�Qd��(��֒D�=��d�{�-�ǉvw<ٿ�^=���h RW��ҙ8��6�N�y/ڔ��A��1!�,`�O��Qq����	&�O%��i�B�����U�ob �	 2y����D�N�pNc���JMm���PcE��]dן�b��R7��[�%"�!0�jb�x.���#�5�D�07���!�*w�v�~<�C���'E$Bħ�1�����2�e^G%6��������8캪,���l�-�asD��y�8�s���`�{ϛ���D1���-X)�j�{g ��Q���H���gZ@:���_e���݌Q	b�4Ä����'��"�uT�;=���؄e���T!,�]<U� �;X�US�<b˚e#_J� #^�\���/�(���N����p�b�9�a�]+K�����x@圴F.R-���
�����a{0�f̠��=3Uxg�e��|��������`�3�6�p92V���,w�~X�:�XA�.���h�iK�f��FA�W��骊�uwe"|����Ė$���T���30ZGS>��b�������+�oOq�.�S�>V�%Ԅ�f�B9R��,%0���EY��a�7~�YE��̖|.՘�]�),�7�����nr����\�m4V
j��У�׮Mʩ(ȭ����J��_#m����m70+�y�2�TFl0z?2��<'!� 1M�������~*/GS"�U,P��PB'�����CZ0	u��O\�D�� ّ����`����R�D��'r�Ŭ}̵�(�J�+rfk�T�<��A��W����i�rA��K*�<c��wr�83�F�Т[�;
,�|��. Hd�I
o Ut���gQ��
,'f�֞@aM���7>ۣE�����dL��`�3n���'��Tg"�2� 윯l��:le�S���/��l��f���.�1����Zj���\pؙ3(��p��;��� 4vB2^��y��з��\��!���ɸ�\R�䵦X.���E����o�0�����J�Z 7�2x�j�Z+����#^�����H�3�NJ%�'�@i�{\�5tf���!|��1_a��P��gOP��q�8{g�+�ᐧ �(�.�^��z��:�L[X�� k�VQ�t�[mUШmN)·3�Q����Q]|K������Vi�ie��<?����!�8��A>�>���sOj���+�����x�M����4�/�Ӛ�����595��^�v!n-�y;i�8�
��9���
��h�������j�b�,�>��~���$�����[?�\f�o+��X�4{%3d�64�@]"�/<���$%���,0�o} ����>^���g�u0l���)�M��CK�i�����FP�7�qU��~1�$ܬ��m���l��҂Ε���?C<=�2�rhEƺ�2��on<̭*;��mG���-�(�H��W����ђ1џL;���d�! 'OkC9;;�p��g��z��+���~�4[�h0 i^p�yK$/9��L]��1�W���.�s�Q8�<H�Uu�a)`���3�C3_�":E�)  >����wJ#�X���&^�!���������G��v=yI�E��L�;��	n��SI����s|Qd�ƚ��4)���Ѩ>�]���,?��X�;���3\�>&�B���e���;n�����=���5���S�ǯݝ�(�/d 3�Xsj��i��v�b���+��L6� ��Ĭ2�[S�4�4[B�޻��1ӿ�zxQt�Z�g������9Q�tW`H�%b��	+�i�Q%��$��c]�=�2s�^#4�-B�X��!O�~8*7*U��""�x49����:���j���М�'A�\�_���t/;odiPI�:�x�b��0�d(_'5�oK��ńxH^��#Ҋ�.�%�\�u�}�r�(34���CcF~,[�*〥�K�~�'	�g��� ԫ�/i|y=ԉ���� ��6 ��C֝��l���lb{[�Drӡ2����-ح��ES>*��g� ��D���gXh����A�`-d�b9wcl�X�G�NJ��ڲ�-P�k�(t+���-Ērs�V��l�AS<+��M���e����^�F'<����a[�s#��>x�pfH��cZ�+&쀰�eޠ�O*WVlxO���48�w�җ�.�6�������^���`�����|%���w����56Ryi{����5��rj�QC����~^��,���?+Bw2��E�粉���� 5��ӓ;�+S`��1T.���;�Ke/QO)~��q:����Q_[flO��j����C�D���JieB|`�}p�?��S]��%���ȶ�1*�"�����G������YX������ר�k�vGi�AY���W��}\�_�dF�+�����/gQ��l�,{:�o�@��$㵂�y\a��%7}�����A��+	��Yq�(���J�q7��,�UX$�-3@��`*B��Z�-u?q�Y��,b�qVI�`���&$�)fC&�v���စ�����ڈby��;�ϟ_BN%���*�(���{d�UY>��9��������o��?��N������@�.���C�_� *Hn�)��Տ?����~��q6e�6�1��Y%����X4+�#xÁ��؉_�9]񤶝�&�l�==ɿSSm�>���T��]xګ�:�ԍ�Q=L7��<d���p�WG���0 c�
��cZ�e:g��R� �X���n;	�H��(u��N,T$[�=Zk�	�E¡�.��1�aRP�:���F���`̃��J2Rnz�q��0r.-�.i�򂏪#6rȱ��n�ވ"�����W��v��|�����aлkkw�G�O�U�,.��0�5	��xdh�ۯ��/�݇a��� ]rnp�_?A�౏o�yn�1�^=j�Ŗ�n*`����}��m�?%ay�]WK!@R[�O�Wv�.@SX�и�����f�]���ϱ+�t���7�������jקo�����YJ-�=��:����/sq����sZH�1q��u�I�F��i��	c�G%�
�S��!uh�+��<E<����{�����蒗P�5T��I����/46�x�1/��l���ei�.̥���X���1��eKBq���/��jDaX�~\V��M;�+�;P�g�@�r�%�Հ{Ŏ�(��'J�a�4ne({!�>6���O`��A�]]�ي4ԩ���Y��aS��FgR��"i��	Y��uW� t��pS�WV�1��cE�S����Rb	l&,pV#��=s�D>�������+�)a���G*�o���`l;�w�����@�rF���z�ʘ��g#�`��˧\1)�$�B�����)�=�V7�ل>
zQl��`�A|�ʝU�ia�R�t�����D^��y���q�Lc@��}M>w[�+L��h<J�!{�V�[+��KQP{�_�I!��'!��O�p����O�)t�.���Z��9����n�3��'��]����#����&2]�)�t)(�����Ś�y+�D�q\�;�$7��v�n2׺)���I�|ss�ol��Wo+$wτJq�Z5#�W�y�	����aw�@w��w� B`vGv"]#�ݘ��B��$l���2?�K���W�"�S�Bd-��[N��H=+�C�+?�z����X�;aweҐA=���yW�^��t%>���ގCj��Z����ȓ�Ib�ݫDL�g4�vp���k ѕf<�=;
��gY���)��?�Aչ����A��W��gpl-W��bX���b���,�p�����q� }E�n����4#��qg�ʩ54LD�
�NI�/�Y�[isU�5qB���8�*f��{ֽ�
��[\�D�����e�����Bco���V���ɝzgR��L�����4��� l��4S�U'��ʇ��pҷU�M���b�Y �1͙��9AvQǄ���jUj��V�x8�e_�үȹ�� ^l��9���{>+�`k=hsU���Cj`έy��,R�J�.��c��!��J��#��ˆ�R�h�ڹC{�H�ZI�e��Z���2����%}���lc��멼�����X����jcc�:Yi���X� ��j����f�����[����A�����2��o�]�'b_`���k�`�V̫�+N��jt��s��hZS2m�C#���~f�@�H��J_`I��z�ܷϥJ�K���~�v��mEт��i���C۴��9�-
^9�4��{��)
)�H���<ɭ�ZE��*G-y���u��e��96�f�&��*]����D�B��!YK��	8�1jWcϿ���T�؅V�of�4~6{D����Q�Z��~2 ݪ�隃��m�>�s��_���*��Z5�\ư��su���I�]�e,W�Y�l�`�̢^�&.�9�O��z��� �ٷ7�%Gm�!�����;�
5���x�-�pj�����wÝ�Z�xX���m~��X���14J�RH>H[7ː�ϛ�;�n�&OLb+Q�U�1;��� ���3DF}�7<Hh�qI�)ht���t~V&m�2a ��[P ;jZ�NOd{����v�lN�[;�k�}�g���E�y��bE������8���.�ݛK��;�1@�Hݪ-�Qq��Q����se�qtC���!Jq{���T:�9��rzm����N"5A��;:�6���:�@�8�R3��>��2�� �`З�b�����ԓ�-�8����^�z4����q��+Ɨ3�*���+��D�s0�#��莰�Rֿ��2�<�k��h��Qz4zF���~/C�������%�-�Ue
�X��U"K���)�l��\w�V�vv
�cV��vB}S����)�O�53��v��,�)��X��C��V�m�=��y��h�t�΄;�^V#���8���<]��=
�!�F�V�Be3n�$w���Y��7��~�|,�|KMJUbJ���:VKm�K*��!cȲ�V_g���G)�)rV��MS�vk��_!�ѡt!���Bm;�y�M8�wbC`�cv�J�$����yn�a�ڸ�F��%�h7Z`Ղ�e��A���W~V�frK��E/�m!�8�]��^�-?sz��%N�kbd*��?g<7��Z�jW�6t�O��(�2zcty^xD(f���]>�V�/���]eKfܩ�G���wY��k�6Y����s��o�A$�>���/ �O;��=&N�/zC2�l��6��n%���<��{,�(��{2L��[�M@(K��,����B��_	~��eE"Eͽ��ͼ6�ڀר,��ZNPH�'�Qo�BU�B#d���6D{��1X|2A9���|��E��6WbL�G]��_!�b��G팿�,n�T�Up���͕�O:�k�]��226��h2Z�?v�al�H~𻚁|̗/%��!��#xF@�+42%�}�4�x��)���z�z�!�$�4���� L����%����7VP���\ҏ�G"q�z��5���ړ�o{R)l�5�R�ޅ�'��3/ר�O�/B�џF��r��
�}���1�@�f��~bխ��1�K��%��ʞ˦,s�Ϧ6�el��Ō\<�~b��^�>���'g�%���QmҸ#i5^��Jl44��Q��:#6r/\9�KU�̀MV�u��)kf���xl�@���z#���s]�<s!v���C0�G�?<��@<���B�h,��0셷��$(�w�oc�e&T��D���)� �� ���.��Y[��]O<�A����u�hƩ4^� c�N͜��LV'��ܬ%E�*�t�q��X,�@Gk�J۰�64�3�޷�֩4����N�6��h�0�0u�\J�����#Q��_�a�L�ԳRA���G&�"]Ϣ(��7�.")�+�1���<��V�B�6�i�f�
�BJ'^�F.�t�ۺ�8t�9NC�����0#�f�Y(��Z >�H��~�
��k��mg9d���c�(�gg�mqp�@V��!�}QU<�������l�(w�*=(�yRxKaw���@��h�B�M\���������� ����.ᤒ%��| �U贶��P#r��P�����A�2T�:��%�/��2#�N�z�I�慁yO�������M9��V�Z�Z=3�plV_�\�K)�3���D�� �r�:���z�&�m��,r]c+�DT��x�,�g�
 
��b/��ȰPv^��ϖ�ߗ%�.\:O�
�_&�~�.���Ԫj�m�0*A��=�2�`;��aN[Z�}7h+O����0�pur0�N��B?�q��b�КK�k�tTo3H�fu�70K������Uk���%Uqު�߹��;��X �H{%����¼�(k�I*W�ߤ��-���ȇ�v���N[�wIz�&�����"ݤ�DV�%%̚r���EFf4�IR�(���>��|����g\���8�<��QNT����h���p���o�,�{[|��eZ���}�K-Sv�7F(8��
���'�Ra2"�p��po$�;�E:r��TO2��Fz.�}&9T@�8_ �o�ͬH�w��"yD�`�6���5_���;�����Vi��u����${�`��x�7��z��bp�?���0�>gbl�bC�a3�$��c���ߙ����^ц�D͜��:�~D�W��|:$��N�M���:>�s�]hBo?�k�t|�Y4��&��4�B���6Cx���+Mfj"�a��0������O���W�#f�K�����~�P!٥[u���r�wa�K,�2E��Iچ�������k��E���1#�u������a<�"=��b*`�]M�(
����@l�2t�Ũ.�u��3У���h9��+���O�e��S�r_|"e�^!����emQۼ �X4nS�Ί4��5�P�4W$4�w77c~����󮧝WG�bn�'Ǯ-� %%�0d��M2��۞Mx���)���8�jjv�;e�E�ϣ�(����WO�zJ-���0V�΋z�;�V4�~o�x�h��:�[$FQ�-sЗ�l۞�"6h�U0 �䋃�$��Iϱq;5u�l��͕ő�cK����P�o���@D��0��խ,̚k�I�t1�w���S���cWPq��Ƅؤ�[~��X�84_�~L��5�8KSU@-�BxUant��C]6��n/�����uP7��u������=�CXh�Rd˒WoE^������Y'�meO-\�I����\Id�-����)�����b�_��p�Wv�2�����q��'FC+C��9��;x`�_���9��]�Ƽ�m`'��ԓl/daa�K��k �R��#̎�ȿ;c����n![�h���7DbW�<[|�4ûz1$felI�����b��ݟ4�������t�eoK^����宒ʶ�P�/7J��^6�YW�3�'^>�"U�|:�A�(�z}!{S������ _-Xk�>��A���~e���q�X9w��a��7���O�G�$���w�7��]�_�l��Щ2���d�қ��� �X���u�w),ke�q���e��Dg�`DF"a� �JOLzD=��^H0Tu]c��i��r�`9�8�&�4�PPR4��(,��$��X�'�;�!E$�~�I�<�5 d4wఀ��<��(�c�h��҄q��RH��T��m�c\tG�s�wn/1Q��<��"�p@2M`JG��� �&Mx���<
�/��֧��:�	�7"���2����� ��x65��H�j@�piyN2�7UmO�ظQ�Z�-ʯI�������
�"���=���h$��}V�x���gx�k�wLp��n%K_-�2��S<��vnu�m��d�����������qg��5�.��.IRw�$�K��*�Y+��>?�����&C7Zi�{ٸd� �H��(�h�7��֑W��ZR����uQ!���2^2~Pe'��g���6�!$�\Ư*�3f�б�f����C&��ܵcbl��mHȘ���y��1bBF�U �lO\TgM�KW�.����h^��F���S	�N�>{[��;�
1WmXq�Q�]����-c�(A]X���sI����Y`gbW�Ќ�궈]A�°,��I$=�jَ�$`���LyT�*n���/�
�7u<܊d�	@h����{�v�\lo&��a]rlX��*)����i�G��7_��}�\E����@�cL��1O?�13��$4�̈���\���W��q~?���@���Pxt�O4.Y�'7IhФ'��]"��M�ѣ�C��Wu�@�5Hߤ���>�P�*@����/|SX��`�=(����`�N�̡J�U�䔑�
Z�^��&�z����կ*�q0�MN&�D�/���I���3�N�5��g�ن�j���ۂk�|L��m���(�6�6�,2n���#�e��A�2XFM����d�~'�S��d�֓#�W9pU�f:�����2�{�G'�A�� `���0�\�hj�X�?r���{���UY�v��+}��[���;%n�@\�zz�+��S)�3+��li-�W���Ͼ�|]�)�;��[�Ps�jc-JZZ2xD'�kE#��� �_���	���06
%``W'򊚸؞E1ԩ�yq}�j���B��O��:��E�X���Ȕ�~�u��Hoï�e�u\����%V���[���{�u%�������*��� u��/�F�fMt1&�{L��8=�oa�6!�� f��1�9>���f�f�~ʊN�O?o����]/�W��%X�:BI���٨"�	��/:��f�Q�_`J�Ή*Q��t�/��2������!n@e�vi䀺f�e��Np�*k�l�B}R����s��=��8wn-�`���!�s�RL��O�HXݵ�?
aY˽���~��|}���L5�����_(.�T�Pu�hb<��f38g�1^��?'���T�8dQr���]+l_l��Hdű�@E�q�Y-3�z_��l�}�\���ũ:��S�ӨB��	Ȏ�JC=ox~V�<�m�!��j�=3֝����ʓ,��ҝ�Nh����u�)̌@}�� �V����-�<�b�@lP����U�2�w�gLT�SG��w�B���~�v��;��F���]
�l���l^q�5:3t^����wt���0��h�y������hCl�uk��HS�A?���y����* �t����,R��ߋ��"�Ay@n2�m��H������ʜ��Sn*�j������Ip"ʶ<��h�;�ߞ���k��ժ������[X��!l��n^���u�'�+��L����M�x�^��O�Tm��D�à��ah�^��W~I�`�Yģ�K���8t��V[_-^�Tgѕ�k[�D'��|���ߩ\?;�(���7,cCy�S��"�bl�;!C�HmW|����+���v�����D��-�pYX�P����e�yaDO~M�_�i�?e]Q�y.N\��z�|:�xJ��à�>q����Č���EF.L+&�M�ɚ�#�s����M�6�T��aC`uH-��^�J���`�	}&���
�3o$];�?'Z�_b�%E�=��8�Nr���Lk;�����4�G1J��̈́{ŋ�Q^���u�&���瀙��.?,[�ָZPQ,CB��/�)�a�B�D�T�H����v �d8�(P=s�ҫ�v>����f�Z.B�����̄���]}�N&���w��u��8-���B5�7�&&��Ld�S���_�=
��@{���q�k#4�9�k|8!C�)>�<#�83��FX1�Za4�a~fz~ᇼ^Ɗ�}kVF�D� qQ�5�?˿b�t#~�G�aoI���1���_k�n|\�,91��]#	� �mqX;�V�b&��Ft���o,��N@Z�mG���>�J�i�#�V�V�sܪdM��?ŃU6��6)S�\�5ʤ�#p�!�O��Oi�0�q(��d��k"\ ���>���m���:Z�j�V}�O\R�粊�C�`�8o�*ؤ��X�k��+ǈA�~p)���Uaf�i���"vL�m�"�E�	T���..�X�ݬ�����W�af���o�D��_TՆ�s-u3���޳�8C�RG�@[��
4���`�\��׏������/e���}{��QDՂT�:CoJ���% ��Мo����8�-�x����=)���FF��Wm���̓����/!Ul��d��д8�Ή~�F���# �<��Xe�̟6�hܙ1���jFհ*/���˔<�sP��a�-�l�b�[t"���?s������@�����ͤ��_�{7�k�u
u�҅���Nl'��`���P�_�OT���	J8��	�S��N�:���{xS�}.���4_4�z)�>�S��u�{�����%S�>E�Gr�#�~m�k=�ħ�&b1c�(��&�r��ɴ��:�M�=}#Z��-hެ��i�Ո�Tv�L�|L��(u��S+xr$sp�D�}*u��@9���u��t��l_f����EГ�2�+�/;ΑִaQ�9���,խx{�f8zc0��mT��`���8K6@�%(#�h�2�}�Y�	�k��Q������Z�̹A2{�B|BY��s�9z]�k�$���3��V�3+p�9N-��<���?���J'G�~w��o��p�_A:g����.�ٲM�ew�йr�����\/9o��ֽt/�;�Iuwn�[2c�Ǽʠ���ʩ����_C�#ٽQ/<��h���Q�v�^$/�e^ϭ��ܢ�\+����Oױ"��iZ�Q�&9�����S2#Z��DZV��x�y��Bu��ơ�"�Y�Ch?��]���I)��ϙ��Sz�����}׉��{T	[B�(�N�&H�(9s�äue{84���i�)b��� b��z�ѕ��%=j ��T�O�o�y|���M%D�*�0pP��2�%K{UX�u�O�	�Z.�1w�ET���:Ep�Dՠv#�(-�U��r�M@���!=��_9�h!I���Jt�\���횥��&���o�P^�N�QIW�嘆O(�����Vj�����QL����E�WIT}Qۗ--"�
��6���n ��vO@�'���2�Yh��e��몬���ڑ�zf^r�w�#m`��1��A�8aA�'�]�ǿ�n3�$�����G�Ev)F��e���
H���T����J��q9��W����QS��Ȁw/�OHd��SIT%� �uaE2j�-�j*���IbM_�W��=_�~����x�$���Ӆ�'��� ���|E֛Wz�M�j�q53���5�Vl{-�y�3ap�澭�l���<,y�^������g��:�b����L��4�{����>'���׮�Tj �s}6&@�w��	�-}+�%�б.=ۏ��u$1ƎW��r��p�������:���6���wG
z�@�Lql�Z��e��� U٥.�R]�F�;���z��n�k�t#��_B,���!�7$�e���Xu�%y9��/<\��up����G�&��<���%�ͥ�0|�~�0	)����|>����v�����b]5�|=���r�+.}����!��z[q�5
܋�/�ͯ�'��&C�
�`��N��L�A�dYZ5~��h�{$�򴦽��涘��9�W��!��7���� Yi��d{uu"};+[yn��ñOm�r(�^��q�Gt2xc�c�5"���fQ��j�$��(�a	Y�3�G.������F}|�&`��R{���rm%ML�OL��'H��/�Ig��ץ\P�nF�X)�(f5K�\ް	�4ݹH!�6����J&�_v㓀�S�[X������1#E
�쳲;-α%��A��C�EP�֝�������z�/l
�K��^��ɛy<��?���#���H�EaVA}+������w�f���Y��
!���mG���/�_z�����7B#����-�߶��V����'�#�fn���[���I%����a�':���+8��x� Omu��������:Q�-O�1���Y����	Ʉ2П�q��X������~�E�����J�W]�M?��2�9�����7�N�1)��f��� �������
k������;왨�dkQ9�<�dZ�d���4�@�'���O�(��Y�ŵ����%_���$��$I��/�0��Xr�O����r��k\ۡ�,Z��Z��O!�7�r�X�5V8�J�qd_���}��x��"RX��}I����x#��ߗ��������X��9��r�}¥V�&�JFy�ɧĶ�c�6�<�O�?_�����>>+t�c�I(p��P�ab��4�N����,Ж�;`�"��=�
}S�E����V?_nc!�"��������Tf1�^aN�ej-e?��'4_�-�9���D��Ch���4Q�?���w%Z1-YkN��tM�����lm���j��{,���E��_��3���Af5qiw�8�'���>�.�����:��Mb[dH����Yi�v��{$�C}�Ts3� ��u6Ț"�UǇNk �~��U�8g�m���^�_jPSD*�7�!�������ꊘ��S��5LY.\��Gd'�#3�v��w`���n���o*��mÌ��a���w�E�@�L�|&	[�Hg�ͤ��\_?|��!����C�-&�kN�m�� �h��T�J�Z]�i@b��/rx<�ڭHvh�ЪT��pɨ�^
L0���A�Y�o�O3#k:�|��Y���l��1�� @sN��}����qi�ib��0��P $�E6�V>�ЛL���.fُh�7?�w��u#΍e�;UjHheq��`���l~Dy�w%�m/nv�Z{"KB�.H�d�΅��FS��ZQ��6%P�wznx���p��D�H� kX5L�'���,���V�}$��ޱj��
U�ۼP	L�p(�`��Z�w�{t!#��j�w^)�|'�ku�6\��i00�w"M�+��R��o�0�@�(oB�1}�F�����?M��j�&1ܤ���o����x���?H��n�xN#�3��,a8�ZM��(�ww�,e��}F9�)�����sY��n�z�KnK��a�
-�?����]�D�� bK[-���d��{�ħ��M����oގJ�x�@@[�5r����턆��Y=�C���Ѡ��a|7������z�Z߾�t�8��xP��x����"��NY�&���j���e���R�;yq;�e�D@��q���Z�� ���W�'h�]Dx�(@=�_5<�S\�|�lQ4ɞSXi�\�.t�;I�H`}�7Q�?\��N-Sr��������vj���7�}�;!��X�:x�(]%��q�=�����H�(:�;?�pǵ�h����Q�N�Y�1����G��,���J}�E��	���6ޡ�Uqwˊ��܎�49�?��"�i��bR��.��A;�x�\���`�=��o\, �/e��ҕ�i;�f_�{t����!�+�?}��2�޿�cS��mL�����UK����$��!��6F�<�0�Aqو��Z���l���;��v�l�JS�F������JEl]6=�2���c��m_@N���:0��@RAG���P���/O����0~ �#����r,�1y2�����4h=�Y�/�C�&�G�&t�y�t�
t��F�Y_b��S_m���d�F���@-��0�]Y�1h���00��!s�0$��Bk�3Ƅs�$dK�V��3Gt������x��c��$l�T�)/��RP�p�$�	�9�\��=k��̱K�!���-ӭjע�2�*%���]�^cdmjt�sRSv6���T+�l�!�۔L�����%x�s?�q.�����QruB9Ӓ7�֡���:b��;X�E��F�J��(��blB��X}٩1�W���FY����2Eh�ne\R��-$#u�#[�V��W�v}M
�6f����_�)j���k�Fŭ\�a�K��X�� \���r����|����C�ދ,h5=�:̬�7r>�Ϟz�M��t)��o�^���װ�w�[�٫^���{��q R�4�V�b�;i���۝�nN�%�G/D��JXJwmMd,��4j#V�<4Y������J���N7p��x��C��"����/�nyMV���z�3f�Ej����l����a��[ζ~B8�������?���eh��]B�&7�.B;���hxb����j={�,��M�-�΢dl�D[v9]{���|�<���mCx�X*݄rS�2�\ ���Ǐ��L�UzR���;�����r��{4�D	.��a$�TAb�Vv/<kX �l>C������R믢v�Q�<�L�<��'��1�Mv����&�`k�e
��B��a�'V\ܼh�l�������s��.������>m8�����D�X��Qp���ԁBz�Xwh#D1�}������Z�6�ꀡ�kz򴂿�
��\u"q�NJqeO?^+J�h�C�\G%쬘)��p��T��Sn�YFajӐu�rj;�~p�uȄ+��\��z>��eR�=Ys>�o��8�G�g|/��� �Ud�SK�0S�$�E�pգ]�7=�p	H��}��[p�Vjy�y�=���eO�c񊼠�hGT�Vm���8�FG��%���;--�~�B��)��b���)�ĸұ��&��Ѫ�O.��Xްa�f`$-����\&�(s-���"`C��]�����b�:&X��_�^���������-����V��#�l�5�����к4V�$K�:ss�%ټ����0m��v�,�!�
?/c�Lq��Cn�!��js��qb;��+��.a��or��K���kn��o����Y~�G{Hq��<�L�e�O[�ꍮ�χ\�b_d�V%��9�4��3��)B;��k����aM_uGf��-��W�إ~{�R�a��Љb�����./����A����z�`�Z����?ͷ�u�Bv$0f賙s�����,8���C�����M�C�~l���%I���.��D)��5iV�������ᘢtӮ��z��E1K�z�C������,fQ��ɨA_�D�Lp�w��<$
��C�C��&@��3`��d��?Y�\z�+�>�� w���3m8�a�aί�U��Y����$�iGl����%o� 1u�-%2ބ�-1'�Q,���iNzc�l#أ��@C���QS��ѫ@�<1 ����.�8׽�a���Φ��2~A؈B�b[5
v�_p�\W>�u[
��[�����>����`^r�STq��̈߅�yU��*��T������e��⛈���U%/����rv���̨޽j)v�� �1J�׫�T��dT�m@(��)l9	��~�ی�D�0[7T���q����ƈN����n�P9��:B�ɏ�di�v#%۾FSk�v�Y��>@��/4���-V����EU[��7>�W�J���V��֋Y 5�E
�Eɍ#�� ��r���K��Kb�]w���;ק�����/xf�e���V��o�wmKbӕhs��|P���hy�1o>V��0�O��ʫG���D��f�j�Ɇ����upp"r��̘��I7
�%m�vd�==y(���C���	֚?��.Vn�X��t5��[��WU����\���.�`v�OG�PW����k�[Z��Oʞ�yi~|��2B�v܋��!m��w�$Z�Y��%	�8�Mfr������~�{��A�T+K��.�����b>|J�����$�G�XE�L��N��3����������W��Þ�l��	�`���cA�c�͡��]䢰蹴�C�5���ÖuM_�YHeޗ�Td��?��}�W>~�!`��y�]��-�?��QIZ�A9Zg��pҟM$ �����|��0=���F��cޱ�'h�:�<c�;��G�\,�+1���&S�LY��[��;yʛ~�/i�4+c��.�Bi�S���*ON��Ɣ��ü��9TC�;��c*���j�!Ջd�&���@��&mL���72�$d�䮭�X~E������to��s)�U'ĸq�;B��OV$cU�E��GSR��|G� ꑂʖT��K#i���J�V�@�'"��d����b%�@���?>�f��?.�6&�L̗yd.�����G�!�h�q3���yZ�Eڅ��E$�_�!v"���ΰԳJ�Ub珂 ���B�t�4�)5�4�9�O�烍� ��,�2�-%�"H�<��b
!o�u����p1��1.$�I�`� �5�k~qq1༑��M�jo�{{��B����B�&�g��;J�,�_J�OD(�T�T
k�n��b���Z��~��Ii�Z �*V~�5�ӣ��r���t��<�Z�F��=�0~�5��p�:Ҿzfv�������u�慩�-䀇�B�x���Б\��1Y`�+���E \���E�D}��$ژ9yX9��m.�vg��J�?y��hԙ�d8�[�9��p�W�яye�5����m��g�o�*�߉�6	6w4��W��P��|��KŁ���UNѺ�`��:�5�j5,�d�V<�z�4��xP�/�V����4�m��3~E�v4�������_��!X�A�֟�q#Wd �Ҷ�F���K���=�v�ơD-�w�ݿ���36?dÛ�q�h�ن��"R����!Tu7쓺m�0C�%XB���:hѪ���FIj���|�T3��~"�<ʊL�dHeZ�R佊1rx Jg1��P�R0�tJ��p��d 9�'b(��,U�!��x�i�Ҷ2�K�e�@mY��ɔׯ�w�����;q���j
�1�a5��]+D&Y����B�b���`T�#�?�b}[{�`��q�5WЦ�>��"�8����<�f��O�)�F	�u�8O�8�Ţ��p��nŀE�O�ŭEt��Ígwӯ���]Y��� �R�G���zYb�
��39n���/��L劙I���Jr�e6 �j&�:�����'��@p��^˅_�T?}�4GxXV�{r�\�.�d6��w�5O�$�{׹c!���Þ��#��b8'�X�X�B��p��Np�04w%"��Ko<tG�$�!���h�X��F$%i�]����L��em�b.ms�x��М�a*Z�SD�'�OŚP¼H�����`ѹ%珂_<�B�K3H}�N4�?m#�ɳz�8v��RN�r�;c��`��-3?R%�^!�t`͙	��S�Me�!Uo[3�����l7��A9J��X�0�X��|�ㅬ�'їf�ujy����B���(.�P�=��`)H.�3)��-D���]sc�Ӟ��PM=S��y%�|���X{=�(���Ms�漈�̭";���CV��܅���^��g��� ���\+��1����F�0��]���%Ky-��E�>,7ŕ�n��d`Ą�=1�o���3s�M������j~G
��Y�%a��Z�b#��ՊA��#É�J��so���L-�#!�n�Iu�(|��(Kܕ�͇��,~ї;#v8v��Nݒ����ׇo�ߚa���2=��������� H���J<v7�tt|��/���.�$�%¨{)u�غ��* (���c���al�b8�L�\�x�M����w�o��ХJ�F�$�^��
�%H��Rց�->�E=�5B�?>�z�����.0kh��.����Y^;3QǇx �@D�?�M������ǭ����pOx��`;�T�����=�``�I�K�T н�V��5���u�������a�'�H1�s�Ӗ�=�6x�x]����̄;�r�����	��`����j�
wO�$��$�긡�,�0�ڮ&�g�o�)�;��(��	^x���YDy���m:t�.@���ȶ���{��ԟ�%�R�Z��37!�<#\q@���[��C�>�h��ﵙC�䢐�_%����q]�uh����~��]e%�������BshH��K�YqSHi�P�gz�.>F����|7�U��P�m�n�����M�W��Wԭ����Pa�t�,%�}�lk�L���N�_����sѭnL�xs�!d��I�!��J�,�醤{��T!-6	ⲍ�̶�Z�����:;�}���.��lߝL�`=�}nȒt�e?�*k�����u��ԡ�82��o�G���-0�8�{蟅t�.邴�oQ�;�h�c��<)�/X�H�6��@�f}�����M�	���`2����}VVM{�7����b�Up��f^���2.Ր�;�y6��F��Z�~�j�,�9�^�5�!�)61��ۢE�7����1,��^������ذs�=�蟞���el�p��l"t���Ʋ+����<9��D�O�{�ƈ��ܻ'L\l,���ڥ������}e���2�Φ7���x��e
u��H�<�ٿ����f�֝��S�t�I�a�Y��^t����5�56S5��E7� HC�x��+c���[U�	����f�&7��U��"J��{���?�]@���vﻦ�$��r�.���OgLE�����0p%��3�,)(dS\���h�ln����ϡG��y���"���kzo�Ge4��P��(�%䘍{��\a� {uG^��Vc���J2n�.R6�V�?���mć$ͦ2��>��:�Y��	/
fE�W�ĭ����H�E�eI��8f��͈���ZTw%M�@��1�N�|C� �6� �g3`ew5��Ɖ�fek�>�m�}k��04����Y���/4��� @���7H �xU!5�D�)��+4��n��G����R���r�Y�IYx!���ep���I�b�D��dl������S
�~U�G�;_�GI�E*���O����u�)���6�p����*�Nb���b�DFi�B�x����o�6�M�_`W5���J0F��ђe`�w�7֥S�cJ&{�Ӝ�^�-��&Ӧ8�W�ihI�fa�e�5lq���� '�/#��L ��>��!ѽ,���}�R�a�~���,�<�PU�Z�0lA��k7uj>���W˙%�">���1��E"�k#W=vL���W)�O૮��&���8
����H�&j��Gb���'4f؇�z��^m���D���@gk1�Y���j�*��t3R[s�.T��Z/�}�]i������`����س��LgQ[��oI��M��On}������l����A�JY%�A�ɓ� ��]����b�(��pSi�ZOI��-ݭ��M�nK��|E؊{����vDDl*�褌�-��S(�-Ć� �>z����*S�M@%0����AxSq�Q��1z>�Q�լ
x����դܾ:���ag�6��^q��%��	��N�|�����,�oD�����O&�a�H�P���^�J�y����!����&Yb� *p�CQ.����9�������<
>��p��M�E���{Mf�h���^{i@�𪮟��4�wGd����2�I�m��+������pO��]c�q�F �a��Nv���q�J�c	�O������1{�A�[��:�����~����6�n %���E�{ܸ*�۝2�����rQ��14#p���X#'67⊘� ��{X�̓(
�=�)G�s�Ҡ��D�����ԯ�1��ڤ�g�F�Z��*�n�	��+�_��,�	wĻ����d+2�`��,ͬ�@ ��n����-�y r�rB�i��Z��7Ԃ
�o�f02{m�G��g"��hE\��=�Y�R��?a�̞��R����c(�Y���)�p!�U�W�(�5���|��[mL�P?����%�?n�q�xH������P<�9Rg�
f(y �p�`�fq,�	�xP�V�3�@u�E�/C��X���m��/|_�l��>d>2�v�;�?�y�<LՋ߳X�s	��CHV�J����xHM0��ٔ��5���D�����2���MV�TY�Zh�Il�hl`��è:,y�e�r�s[�P�/S�fY� ���N*~���k�*�p�_,��I6�H�T��W�F۬Oi�~�UnU�'3�@�s�R]!('�%��L�I;�gn�l��o8�-���*S�L'"�Yv��3\��k������T�8�
���9����׫lo9:H. �^��|a�:m�7����9��о�n��ҙ70,= �	����%�2D�>��Ke4�9j��(�!\-i^��jH�����a�5��e4;�.a�[QOChwꔆ�u�]W��?V�x�
�R��(*&S~��ԿU2�" Ƚ��eKs�Ӹ���|�n|6Z��Sr~��+%z���U觼�=�6=��C1�Au�)���;x��0���0�2����i���4�w���+��h�f��A�o3�R��ÿ�~Bp)\1I~��E��Gr� 3�%� ��K�&�D,d�%��^�����؏TG4^z�~��t��S���:�������d� g��q?�9�	�9��i�`G�q�c������4'z��� �Ep�ٵ��{����/�`�(�e�t���!��3�� �����-z��bHҝA����䁊k.s��0��-�����N���N�Q9�ދ{|�ݰ$�6�PH�L��I��B6�ز�o�w@�2����y���Sui�e��z��J���S,#7p:o��u��O�b�\_z�F�A���L�T�ko����>|ݍ�������������'�c&P�����~%�,xH���1</ʢ#ĠC]�C�"O&��[(i���K@@`�1I�K_a'��s�� ��B�+��ˈ��а72� Pi�,��mݴ��ʐ;�U���ʖ�@b�J������^�7x�\�z��ϓ�����'~wsM���I�]��&_�ʤ���b�Qm̈���p�����n��lk��%Km����^ن{�^����1��b�+'$/{��m�P�Q�,T �*Ụ�HQ��U^/�{�����v�~w��V�~�O\*����,�_�?&'�l^�%�'O�z�ؐc�����Cz���i(K��x���f�q̯j�K7a��=�-����-e�n�$oI����5�7����й��� ��\�f���>#�J(����(��h�����b�qP)�l��D'�7�f9��9fT�W����2AJ��m��*��8T�{�
�<��xA&����^��_�/�[�"�;�vq���OWB+�������U?>����S�@�����@����J�d�����H���π��,�G.�@��1#�Z����x|��B�,/u��`�$��_��]5A߰2_�BĶ�ڨ��r�TE��RK�l�J�$}4�G�V(��FQJ�&`&��ߞ�/l>��'� u��&�L@t���J;g_��E��: û���ً�_4L�����^��� �Q C�(�3(U�1,U=m�B9���D��[{�ô#���.�ՙK����T�6�Q�ϙ�ۆL������5|��_Y�:ᐸ�E�(2���Hymݱ��)�zPT������f���� ����Yh�:�;Z�Y;���b���l�
��)�Յ켛>�0ե��$�g�1�$*+���<���p/��[�Ï�LY�i��x�{e�D�������F���<ο�5�e���WQ�*���S�A�f�#�����;E�!�&�����mY�mA�uƟS�<�Aز��X�0�ӯ���y�/2�[����(g|\�vD���D�t)�k��Ax1m�ou�u�2x�� �6��K�ݶܾF��͍���QJ����Z��z15����?�A� �q�іtz^�*� �~�i�#����goeu��!N����1�T�������[+�AA�X��㝩��Dt����_`>��8��j!$Ӏ�* �%xx�#U�W�^)��oc=��S�z��/h`�ݗ
@�1�i����H��ኈ@�ݿ� �H��ɀ�q�(#�^aܔ4	Qi�Ȋ4�q��|���8��%0d���� n<�c8��|��F�[�^��̇� �
�u�;I,b�ڠY�K��ʳ�����!٫��hњ��蹎�Ms'n�ˤL�����n�)E�Ua��,�!�C�����Q�¬��N�@���7�5�=���a��n�D�^��4�S1���d�KU������a~��@�P�Zi�a�J��)kD�}�p��5�1ɭٓ�yka$A�"�wڎwN%eDD��
CN�2V�	/!���m7��cQ��0I�k<�#��O�f(��������
���^�l�
�#Z+݄�A2�)s&ܺx�s�4)9���kR�jɶ1�KO-5R�k����~��+�0d�Y�C�R2)5��Cרv���Ϧ��Y����ɡ�&{M5}w��W��"�'w�ɽ��^���;�li��c�H9yu�=���8H�s�QCW����hk���{�m���H01�o��r�0�h���J�
�&���bY��>v�a�A_��� ��!��� pua�Wg�"*G���)f�S覞�����mYA�h��R�u)e��نcc&>������}�x���NT�����ǁ�k�Utm�Ҹ6�'7Mr��+O�䤳�נq �z�T�%��1�DH3�6�}쇾�o��a�A����]��a�ܢMg�;*<�#.���s�"�_�$��1,��y���-24�t��M��t��B*��p�N�1�����;8\������%���R����<ڽ�����y���Jb[���5����2�`>��1�x%4�lw ���M��O�H�m&6�r��K16���<����Ǣ�����9N�+�,�`���|�x�U��Q��O��f�q��غ�rڴ��L���YH!��尪�\�(�2ǉָ~T���/%}:p�a.|�o�W8G��,P���Ƭ@�Sԍ]��@4����>�Q�9T��F7,�0a����M�������2!9�	�ia	4�J9�$O�4��>V�,��0M��'}�:�|U�OT3�BH,,�ΪM��w��D�1�Any^�q�1�
�g�7�43��LJ�FG7QU�y6����������|i{�]N	��>S�)�k<$���U����}��+5BΦ4��Z���+0"����#��Re/{��(iP���5�c����۲�6�Mu
�$�d9��}MB�^���XE�5{Apv�5|�Z��Ɏ*������0Qk�B���.�A���N�O�/���r������~S�����+�'%�5@��!����xX��۽f�w5QIgBN;��E5��j'GQ������#ޢ8���	���Sz�a�4��8�j�z8�
ѿ���c���[C�����o��g���'M�ݶ,���&�`L6)��������	Rp���35c���.�23�Y'���1��
��7��q��������c�]���FfH{�l��5|N8�P�(w�Z� K �x���a��.��3U�n�>n����Y]��WF�v^(��H|�0	���l�ː�{nR'�[��9�^�o������k0�
$H�$���PM�n"�ښ�U��$�E]�]۵�j�E?��&F�$G��,�5]���+�[W��^�:�%�E��9��Ւ�W��.'���zGeu���BU�[�u5�T^�z�𬠰冑����-���h̛���=��b@�8Y��Z�5E���qb�=�-�z%6m'8-f$`}?ѧ`�P�7�0�5���X[��)�[ʇ	-�%��g�F���b���޻D�o<yɱ�1��4,�	 -�8��8���m!$q�*��ɫE�w��>��������(�K��Ǹ�����3 ���.O�hg����Ot��=	6�K�Qo��*�."W�n��T�qI���΋Lg:?��?p��Wߤe)g�-@-+fO5�5�W§�W��b�Y?�=#�qߡ�޿�V�PF��l�c�qE���7����u�u�%?J��&���o�"�Tq��ʐ��Y_\�j����ZO���G"qi�IGL(Gss�o('�� �����H��s�$l0�x�#!�5���Z��$��"}���&�r��<����B����I�>��t�J�0�R2��SY�\���d�w�ˍ����r+�.�
yo϶���H�tFt��L�����0s�A#l���Y��.1%9i~F��Z�k���b�
N��9�4�2��6��p����fw�Y΃o�ي�<�$!'@�|'���d�EZ�/��O�����@��%�U� ���_r�+�J�c=��m�Z�I8eb��ݿm�u���J�h�ϓ�3M��4'?[�k�a,i��6�/��E
`ʇW��7Q+8�4�h��ncbQĭ�N�w�|�.��e(N6w�b���0MC�c�"�-<�p G����a�鿯�I]�j��a8��)�; P�q]���e���B����3VélfQ���5S�T;a�D":9!\�������d� �5o��?�1�^L��^ �_�uJ5��+�
��ih�!V
��W�"1t9��e������s�y�ʯ��[��y,5 ���yb~-��"����.���$��tcW���C�mƳhvI���U����h[�욶y�w���:,����;5�e�ɥ�"A:]mz�lnmtQ�|��JQפs��*��V_�+@�6C���w8�y���9T�F��݂�55�4۴��y
E��SA8��g<`ԛg9w��se���32����0�������/�!��6^�c�&E���1Q!D��YE�4���gw�%؋�Mǽ��3_~�x~GA.��u����@��kM�%h|`�P��w:�u����І�@7Gm��'R.bv>b�?�KN�_������j0���i���G�`�,��P�)��x"5��֙<����K�{hq!W��n�4;����]"�M�'��IG/���V�7�ڍ��Z:���Uau�y��]=�.L,]«1YI��P����p��T&�8��
���=sޒM��(!6K����-�W�"���L�`��C��#6���e������y%�I�S�\&O������<��)��ձR�37M���N[\��~�RW�h�N�~/<q�N�[s����?m�k���, �eU��n7��e�i�����ٰߟ��;Ysh����F8��vЩ�Ǆ�ִ%p[	N;³���@}?	H��J���&l���wG�-�D��:-,��%���8��X���X�ECckh�D�F�98�?r
�d�x�*@Fr��'�Ӕp�Ú�a�S������3�4z��U�a>�A��\[_��x�:�>ר�$T.����ӃD"hǞ���f]�R%�����i��2y�v�w�!P�][U��U�њr.L�+��T37����k�.xh��s�A7�]��3�w�w��?c�\�\?vA%�s��d�j��@Z�/�i^fM�k��9u�m�V�5_1T46枫�l�)^1��(W�A�5���.�?iI�%�ژ$��)g�H7�?�=�ro4�8L*����
fr%�9�"_,�m�<̴�?35��w����ۑ�)����@s?����
���r,;�al+%U9�)�\���ݠF�
�38C��s��3�p���rP���2ȗ$E�����������9�r6��A�5���g��1͊��I����H�|�.�sKs��)K>�m��5���wM8;��u��&@�aj^ъ\*>���c>Rkiq`�83(�<���NM)����{f�_��nw)H��B��a�XIO'�Pw�H�>q��c �κ���D3�2��@M-b5�譋H�,b(��yi�	�wU�Li�I��{x����)�x�ԑ��ņЁWq�4�{���3)�?�����1C�jYʈ�bG����Y��f���%Ϳ���X�IM�~��Tz_���k�?�4(~�('Dt�tэHd�O��5���͞�Z��z�kj9yZx�4m����T��d�8]U�OK���F���YE��k���|�[���e0���ַ�[����U���p�A$���E�����n*_yb�k�I�UJ0:N���
41�p>a���4�B��w�~�q3`QE�8[l�A1!���@�(�g��վ�v�s���6=q�(����p�+z�%�g��G�>���o)�nt6vaw��!�\9�IO
�o^�k��6�Q��d9�%��ֽ���E�%�
�4���ҫ}��߯�r@M�m|D좳	Ӟ=���Q�?v#sk�l�n�lTsHI�	���3�:8,�����}걿��ָB�6���(W���IM���ĀBmт���6և�h�O�=9�lBh��GD9��p�`MX�7��ۦ9Ɗ��t���n�QP�'s�Qb�*;�5����5�:�;k"%V�2���)�.��%vBE	���
,^��D;u�P���5����u�P��� +�w{����m��j�Ņr�?Zs5�z�46���6� &j!;a��ǂy���e���l����Q�f�"�*-=}��pI-��-�w�J��o1�lK�~p��Qqdd��JTĩx�������.(gi��ʽ�̿�kA�`t�.W`�T`�����Knb�� �g�uA����I<���7�JR�Z��`�[Jpn�՜��ɭlU���j����=����<r�����6������HF	�y�^��kc,ͅ2�A��/�:��`o�H�I���h����LC�x�Xl���������c_-q?z7����,Qp
}&�����M�Y����%��� 0�P�aq����u>��ï�|�����`��=�?�I�_��v3��|�,�|p"��3_p��n���Lw>]�[�j֑��{�l�Y��fa����t,�����o�N^S���<�����j�f�	?e�$λH�üD8!�$2r��ԫ&A F)qYA�<R��Y�]���Ym�=�|�I]��:��`2�\��~&�I�Ւ���|�.8
�:&���xX����)�[��15����P�l���8���@dD�EK*xX?�����>MOL�$wS�����)8S]�A�p��3f%�p�wV� B�Ơ�;��O,_8�f�Q���~cLУ��nt�!����ciX�����SIx��Vh� 5����^�g����M�7��ۉb[J�5威!y�{��tR`m&� ��� 4�d(���{ l�G2U��c9-�e���^�4ᕫ����A���I`�&�7�F�u-X���2�Dj��mKU��itoU KWG�7��i���^�ޙr��K�ἫS���g�r~W�Q�	C0�/�ج�]�<Siiq��#x��q�����)]�x�)�a�e?���E�L� ���̵�Z�6;[m|L�u՟��u�w���T6���vߺU�2Q}������8/���캀�z����O����;g3a|~
�/Fc`_�#��s��Zv�G���,�tbw+!e�ѥo������d����p�^�g�d�@�Y5E��@iw� 6K�J[`�?eZ��k���&�~���mg��<H7h&�[s�DsO*�}Baq���g+����_;|���w\�z�������4xP�_�"g���`��[�%jh&?�p�A�\}������}%����'>.�.�Մ�˛�Zӓ�bp��l'fZc��@[]��b�N�L��4Ѣ����!��T�CO
ܤ�`lNf���YN��X2��R�l.�0Z��-�}/x�#"q|���<��5+5���D��{�(}��(�S��*�CB�]��z,�ކ�sƻ�w�"5n#�	�~1Ҳ����F��~�ii4��k���he�ӚI0�ؤ�Zm?�u�AH�2@�>��ؕ�S��Z��3��/o8����2�
Lm�u�g;Jw,��7A7Mq�w��G��0$K��i�u�ҁ����k�����W�(+) 鴓@4z��TZm���⦲�T��	��{=�na��!����x_��N��,�ǻ����&෻1eø��]��x
| 6q�����!��Ն�f*B��A�.��u��͢nK��7�k��~~��/��^��r����6�$:�=յ��YVd	R1+j���ϫ3����_�(7��Y8���{v�a���PSb.T�5�F=h���o����ܮy#���EM��g� �֫	r�?�t��쵛�CU��,�rq��,\���ov���i�s�W��l�2v\����X6)��A��t@�ҭ4��0��qj�Ԟ�"38��t����wX&�D����%{e؎g_�]X�T�]�%߅|��^;�?��{��w��t�n3���r�2��IV?*(*���78,!_�e��f<=O��][�p�:Vu�� �@�mɁ�S����>,eʽ�W�M:� �CO�L�����OĲ�%�z�wx�XaĴ+g�ct����suu2�@���4T�[%N�'B���@�����d$j`\>��[$O^�s9T�7����x��ǻ�-$r�����%V��G�!�
�k6D�ce�MrY���bU�G��c�8�!�UY,�@�o��Dɦ��>p
��-3�FcH!;��>�d#��ԓ���\v�Oߙ�Nƭ�gd1)�Hc�����Um��`s������&)�����l�����&IZ# 7��� Ğ=�w�l����/�L��^�R��49��0�W�xw5?�I��y�&v�j-|;�S����-6�P. 6�E�z��hSӽ�
�` �ֻs%����~�z�h��u������Ny�0�3��i1p��䈥0ƨ]'�n� z�qF��0+\����3��-}�y�_����O�	x�56���Nhg�#�$��Vvʡ/�Y�d^�0���5�7�>��V(+���O���L���&w�?e�  X��
��	E%�������E[��.ڰ����H��{��(���K�/66p�XS�#a��4�՛�qz˫���`@(#ăח�P"��χr�n��C�j�[�T�N2�Q.�U�a�ekW�	T�g�d���!�)�M��b�}�ɺ�#0jP/���QH�E��cd��Y��?���ƶ�
k
��_PT�����q��Hɯ6z��(w�!� �����݊tz����zal��N	}�F���7�Tsc�G!�z7C�G=6"�}�S�ʁ�����������"6�3:p��C��y�
M�3�Q��~��I��Ǎ�6�5��"I���@�I�HCN*�[ʦ�~�!�[���S�!l�,]�Z�,g��$�3��#�(?P�� =:D��,��_�����ϻ�����s�ej+�ct�k�W��
�q:T�����w(U��B�y�̣.� J�/	�Q�)r$��
�	)�V1/A�*=oc��<K�*(�U;�Ã���𲭓���#Q�Kp<����6�ϣw��f��R[�s\6%�c���x�.2��Y�9,��V��y|v;ve��-�'cF�տ��R��@�Y����^Zx��������μ7�Z�1���"U�k=�~����?�Ĉ ����̓�)�%�Eu.����]ѹ�令�5�LC��ZقS�G��q���n����.�U��Q�ODi]�R�:xƫ����n�-XV��(i�j�������1itnY�'d.��q���n�8� 5�Ŀ?G�a!�egj�e�g�U���. =��ĸ�+9{s/���{L��G��ƞ�y%�G�0�a��rF���0�̏(	��B�P:)HP�)DJp�	���&�ң����>y7䂄��.�,���6EQ�����t��l]4��I�����{C�.7���� ހi�l7BK�C=��O�q��g�fֽ]\����37�d��V�ޝ�Rp���<[At>#�7�d���X!�9���(��ȥ�d6�eK�aؐϼ��Ct�RPN�{+/�D� �c�Zޜ/��H����b0�I��G����^�5b��kS�K eޅY��Γ�	�K�h�!��:;%�6∆)�݌���S���Ⱦ1k���vM��f����r-��q�a}��kňy���/h�,����
���?��9�
�kr\as�=��"����CCyL�����*y]k�#W�L���!3 }S��1X���z}ͅ���5
a��<Xm�E*����/A��F �(�c~A!�f�=W�#�����@S���ךy����	 ��3ûC�����!��z*0?�y��Ya�T�&R�0j����h�#�.��0�wp�'�p�\�7T� Z�k������OR�XP(�w��m���󁋏��g+����u�@����|T�FA�I�9�e7�e�F~gA�ZW*g��F�?�P_���jk�}�3��{��%*��@Ǖ�7�'��{͑y���� e�9�sq1DA�au����r��A{@�<�y�{59���r����cә맄�|�͚��u֘�WǴb�7`�t�]�#�G�4 -;��|U��\�FT�#����9CtQ+G��7����I�9'_Sp�i+Zx�ĜE�-pO&��+�@����g�L)H;�h\�棫-G�c��)�z%����&�M2�w'�;΁8]��BN�J���I�U��U�n�X��]l�S]%xz�n����Y�Ƽ}�+����-�<(�x�\���=x����T64��x�����$�s��B�,�7��=C��g�3�({�K:�͍i �}\��+^k I����|x��鄔�h��p� ������Ni����R!����8�D�mܚRO���)R[j�r�O��i��?&cb��_��v�aJ�cY�4��ڣ��Ȋ6���!FG�o��M���Ǩ�=��]��v�(}ڇ^�829�����7Ḯe��JJ��5\���#QN��! �,��G��5���;Wˆ��%�������&_vkb*����}ߒ�ܔ��6C=�u�.�pj5;f�Z�����a@�N>8�5&�w���U���]8zQ n5)�~��'bz���5�;Z��m���PRZ�o�6��(�����&�@��;� s��S����#��ƞ�r����0U��7:"�!WG�#�A�ll��G �� N��'�F�^�9a����_�`�s0�)������q�Q�Վܙ�����ŧY��d�jѹ����<�@��w:mr8����,�% J�>���+�D���D�	ypUx",y;I��ֳc����qx y"�$ѓ�U�I�.�e�ANٯ�\UY�Og<[b�൨�Ѷ<=��G�\Y��~�'©*�>�U��{���ܖ~IW����.�$Dƹ�Q� X%���B�tTj�nSa�����u�b�8q�n�dA�g���WKNft~��m��������Ƚ����ގ8�{�����v�[���D][r���7��ټ-�<�Ҡp�m'JYc�W ژ{m5�n�j�����By��p�v�s��5A��AB���∃k
�f�m�x�6�Ɛ9�i;�U�Tq��=2S���Ε���~��E���Rl��*ͼ8&N:���z^ψ���X��˳X_K�m4:�P���;�>���|"됕<�8��v��/��,��4O	�`q1.K�Ow�Y��{U��'T=�(m�� 8�|Hϓ�$Tǳ3��c�S�FU0�ӂPqQ=m�f
��3�Yof�j�%��Tϑ1E��K��h7�60^� ?$��\-����\��rj�F����<��8]
����`����G�Ђ>`����~!�g�c�+�IH�8���_�:5(t�'�ovv�������U��^8��f��c����^�p�0P܇V�L�4VJ"������0�']�(��^��mf#	�C�Km��aڠBX�Ž3�40�L2�rN���/���G7��w��gڷXG���y������X���t�r?.W'���#9�h�`� ���Z��;9Z\�����t�hql���e&1;U�G��C٦�π((<�?R5��Aa�$�dm:�kt�����;cop���^Uk12����A �Q�<u�`��;�[ݯ_���/ǞD�عd�Jwܟ���"tmg䆨�ݦ���!WU�Ք`? �`ԖA��d��f��D�%LˤQGum��4(r���}wF_����RJ`x��	�A(�~�^�ô#C�`N=s�+{�P򏟔��	���%7f+a�<�n����.�݌6=��ww����R�]E@g������-�_����4A������{�lK�[M�~#�F���bT�m�����&�c>���N���ao�CU��M|w����\G"���3�v`��79��C{�M�/Ł�יw�@#-	]��,5���x���[ַ'�$��̓�<z�JŅoF,_އ��VN (���Gˢ�F�Z��:��bl�ؓ��+�%��fǏ�`t�����pI��}CZKEN��Z��ۍet(19:��/��4}9�R`��]��@k��������k:��0#e��Ժ�^�+/��A];oan�QYZ��XCF�N�X;�P��s!�`�8��I�[���ZTa�i���^�0��S���
�����. ,ex�m�ۑ�Es����o#��E�WU�H�Wt���f��x�AŚg#�I+7����-�=äc�����#��qxf�gIKC��8��K��Ԋ*���G[9��2��h7S�&���=�Ú��(%2�u+eMȽ��ю;N�{�8JO��WT�G�뿎����OɲUkt�W��Vǯ�(�I��	�+�t�B`X{Y�cp2f�Q��0ٯ��Tӟ��D�bay����]��`�L_����`6����TdÇ 8���7Ts܌�m𘕺�����}�s	[6�F^Rf�y���y��KA ��C� n
���p�l�ŦNv!!=����tɺ�0���`�YS�DyĂ�~츋�0|�p�� �@��)v��ҿ�X�~��+����#� tUy��xz-փL���=��7��H=T�c�n�n\�
��Abg��)���;���D����%s]8��N<ܱ�ts��V���z��B����H�.���I�GZ{�W�}i���u��I�'�r�(뢜�>H[�kE�H|=e�_w���'��T�M���v�����UCzʘ/8��^h�Dn'��_֐#����.�����y����շ
����u��.3$�w�T3F�n^ޫH���ϰ�S�NA�M	�,�Q���O)����0��4�����0���2'�Z�fe��f����"�}�l�gF���ǩ��U%5��&`�.[o� M���8��R�]P��e��>�f��V��bj�o��;f@�xAa���Lb6�7�O�lA�U:�chn����R˲iMm�u�����rH�����V}�����BGb����d�5n{m���0�3�e���X�螛�w�u�/���|�����&o�zT��Y�ZJt�r_�oo�1r����}�8辝�'���O5f���ֺ�~'���W-8�t�O�n�^lge�|�?�;�υLUŖa���$�N�Y0�r}�(2���)�ZH]��X� ������r���W��bY�9�/�/���"�D�i`���Ny࠮�N��gB��:��Q9��'9"#n�A,k���D#��E�5`�%q��r�sG�g�2R�B����~R2_��X��Eph��;{��j����a�fL5��b�{�%)#J9��s������+�s�� �հC�V�}����]�G��6�9�w�}��"���Xr�#5��#[�{s����?H���*h��Z8����;K��+Vi*����n�����[G�^g�9(1�"��P�����hKR��∽aAk�s����~RUܸ�
��k�u�:�>��H[�zB���'�w�R�f2%���[�<sFs1lP9f?��H�6+�V��?O�<�L�<=��Q#���_���J�މ��1D�⩟��l`�	#V��V WoM<���J jb"�ֆ��1���!�T@���˫�;��nѣ�|nDbsa�W�ɷjLf�u"Pr�l�N1�؅�.�6I�oF�j̘�/��wO��C��������O�������c
�l}�^����yLfJ���VmQ�R[a�w�\���	 ɛn�m%��+��2c��[�ϩeK���̈6	�WV!��OJePV��!>g�gT>���V\*f1�
�,�>��ʭg���?�_s���z���^����Q^Yd���o2U�Z��2h�Y&����#FE��1��,�V�S_C)fA-�$)����� �fZ�{ɠ^x���-y=)�����\u�ow���[�>���6/�]�W�Nf�]��",�����=!��ֺ�V�?x�1qX?��b�1ʲ�M��48wޤ�V��ʎ�F��N�#����
�P+�k1��Bebs1�J�P�Q�ɑ��I���!�6~z~�\,���P.���)��`R�,z��ғ �{wf$�0�ѻux�q���^�/:O(y���Y�>#���6���C��H�wgn�A���1�������-v�jh_P��*�¹�������H�l:W	-�xm�3^�WC��qъ��0��ӫ�d7c����3���yxg�C�	B�=��H�3���*���Ջy���K]����]^����	!}��&Y2N����� �-y���C�̑Ð�l�Z��C�ro����TS�h��eW@I��Iz�QQ�*�~�_ON�������fxg�`�\|�_Pܛ̍[�����p@p2���bsz�<��\�XΨc�F{�v�a(J�<p�
�*��W/���8����B+�L�[�"K���H����f�KZ0E�#���ո���^)�sP`�
S��@�s䓴�z��$@��I�e�=������ի���6�&��@"������]Y�~ع�T��W����Y@�f���b"�P̳'�� �Of}3�}��7�_�wT�kcXU� :sg[)<V#�`Z��������:u�
�A�@.?�Zٱ�r�8f�F+�,&ކdi�`��2+�@}���1��������%��7r�bXW�q���6-� ��^5�y�r���NW�S����OY�zn�䅹�����}y�&M�j�Tb���	��Ü��e�{�5p�Tn�
v|3���P�x�,0�=��qF��U��`��=�TX������B$C^�R3龭F@W��
�)�2b��:�I����f��C�qz��TL�/Әg5���ڷ'�W�;�������Äտ��	zD���E���e��͞�e��
����-���ʌ�>M��'#��v5�H��&oߣ�<��)p�0d�Zo�j�B��|aV����MS��X�c��.w�T�;H_s}Т`�&�q�0�k�цa�@.bG�ͦ]; k�iໃ$6�������<��w)��������?�ѭFO$g�>5���Ark�'�φaz�)us��U��5	bd�M�H�B�J��I�8O�R+
ݮ�K�r_� ��8��c�<���e�Q�gm�@5E� SNFQ�y�~�9��e������kz����I�d�6�)Z�l!�/G��L�LR�ъ��Z.�s�h�05�[�UH*���v�WpNp�.�$������,�3֪��3�c��رKN�~1ڗ��BJ-�#,/��M�TI�DvA~�!�:p����ޱ����"G���i<�LK��Ū��ŧ�����չׯ�{�&�Kɯj^�a��[r���-� �\��)2[���^��j��@��ݎw _�`��
We��4L�y���j��ҧl��_r���:g%(WwgAlNt���������lú���Ί�^_�N�AU�J�ɸ���^:f��F��(Z���K:#��M4�=~�?D�����Χᤨ���!�.���*B��!&Ӗ�3� ����L�Q i� �hmհV�s��=O�+��sn�����q|�5J��+=q�9-�.T�&���J �nE��@���"�~Y�=�5?�:j}���qJ�O�>�D��X�Kxk��z�G�XAir�� �5�Ǜ�Z��gn�#QY��A��ym��>��ӒJT)��9��A���d1z#+�h���1젒A����bu�T�"T&
8����Ȫ� �,���D+���=��5���Y�6隸X0�7�#�������+���`����UsU_<�/�_l`��N�����x �ѡ��kf�j�ƃe�%J	���0��"̋l>�z��ǒm�2�[!�]{'7�R��S+$��d<�:�=�c0��/n�x��хPq�25٪�}/x/Q��.��^���������A:��z��o9���5�a8������]����,��Y:xb�%phP.��q�/L֩�ڡ��o��w��� aR�4ܧVm�� ځh�_��Vܮںls�L�Y����\L��S"�'=���ذq���.hn:x��:BTI*)�9j���'�.\�Q>~{f�M#�(�B�sz�
K�7���3TD���濡���Q��P��zh8�[W�u��e�ځ'���N,�rف}�^��}�B$NX�߲۞~���
��j���-[m��dкJ�O@2��������n��T�}2�y0��a)�bޫl�)�oֽ��%c��@2 �{·ղ2X�?����82MqE-]�|?  ���͛�i�����WP4S�K�/dҸ�+�<ŷ�~�VnE�yA�^�\���y'STԌ2�g�ooC�q*��[�o�Ԙ(f/E��LHe��yT(��*�d��k��Í��Y]<ߩ�O�0]P���ແ��o�9(�Qe�?4�tF^�]xj�0L6��y�����*�d�iꬵh��r��h��{L�"h+g tz����A�b�����~���_CA`��������݉T���δIetD�Ρ�>�s9�67����kV��	]����d����=v�
O	�V���\��x�19�I K�� z���"����Jvuh� F����	�?'Z,}�!R��]92k����wH#q�i���������~[��U8����Xc� ����bL��c,ï"�q���"'���oV�x���\� e�o(�"l�f�\IR�qk��A�.�
���Is�B@f�C�N��#,���M�Pck��-zO��Ѿ�Y�ƞw&��rQ嬞Cea��+8[}l��Lz.�:�s�:a�v7��4\�˹A�3Z��ζ�������_%��~��}�;��ΡP�"۪��}_n"�Cwm��L}{ω���ٓ������=A4�r�k�.�}�3����-8�	�J�t�$���`I#b�8�_���8�0E���+m�+���1g6���Օٰ 87ggS���;�I���ܘ�[�"���*]Їbx��#c� ]�_�%�g�R���%��<.��f�����uܶA^-Pj���:Kxx]�����/m�
	�@�TT(f9"��G�)�n�H�e%:`�}���D�r���f��oL(F"W���¼�%��´�z6_���v���c&=��Zl0Ϥ�y���.SƊb�GMO����6b-wV���A�0ڕ��M
|$�iˈ�D8���.��,�A��LJ��8�U>U��͜�S�{��\]���΀��k�8��I_~Ϲ8�䕉 �J�'���NH�����ρ����XWctp�)5�����ܴ�7Iiٻ���Q24ѽ�{�k���ұ��.��w6#d�&�4j/^[��!�0�R,���e�7l�-0�h�q������,���u��̓D9T,�նC෍~*TK�0ȓǷ����i뚙E�z�Xoe�Ԉ�7�v����h��99[�&�%�����z��V�9�bJ
�LQ��_3"�G�r�ꛆ~T�~4���8��Ľ��C%e�Zy2�i�P�����U��Ǯ�����d�7꼬$��m����>���G<��=�v���s�њ�F��(��e�5O	�ǚB��m�2�-����R��S5:��<z�8cXe�������ffӄ>��撬���q&�����"��\-��6��Aʌ5�Ay�A���A�C�7K\�|�O������Z�06#a�(P�.�� �p4��&&�q����]g�o�7H�E�7�/|�s��7M���!�_��s(� ��?y�^�}`\���s<��Et���!�?I�(��
��5\,q9P�V�7�QI�x�k竏�p�3���#�뮣�<[�T�G���+��� _;AjQ�i�:���M,��	���@�xY�<�\Sqf�R��mwkO�-�qS#R��`��Z9�FU��(B���:�j���z�MI]�\��鵟	�8o&>Ũ/�$)��qyoOD}�'(k�����9�X�� ?�+�}+�;��������a����u�}e����0�=�/�#T�u�o�H¡��n�O�z"p��0�����Uڎ�4�C �dT:��d�q�9�j*�s��ՒL��'��E�3�%��j�;��
jJB����F���6�eu��4��y�p&f�C����Ư���:�\J�K�W@$	F���/�&�R�O��͵r��pZ��׃~���[m��̊�1�n�K0�U�w�;�ή�wg�>�N<^�Q��4����/�;��T"��yM�#�WLD	A���
<d�.2��N���9����I��{)���oְ#�����z�>�V���� l��,�]����uS�O�Q�rYbJ9��Ц�P$�4$׉P�Z;����ŏ����5���W��q`��A�+tm������Ȅi�Fcy�ͼH,%��ۉ���-\� �5�zW )���.!B��5R-����v���4
Ա^�~�,�_rin����OL����V͠=�9R�}��{g�]"<��;�Wq[��6��i_;��ŕ�x���P��k�E²lS�{�a���]�Y�y6t䷞e�<�5��^���V�R�N��,�ß8�{b5r	3� �Np����ʭ��5�Rbv�*� C�ɕ��>���$>�$֮c��]B�id����&�j��8b�����N�Օ��^N׺����GS��ާ�]��R����'L䷯P�6��9{i����sL�Չ�!�N�	F��Dl+u'��zz\}��K��՘��#�Io�(��ߩc��������:k8s��#�U#F��@��;��D\��lz��ta x)��OV$k�j���/��7c�|+�[,�RI`Y6&0�|1�ս(��g����Л戣f):�Mh`��ɸ�
.����O4��W˾WYA�Y_um�O�t
���\ �����%��t˒b$�AMu�Nh��D_�S�bU<2���}��Nﰎ��>n֭r!7-#��tb7�~�?�h�(C�U'����ƺPn�؛4>x���R�<G���y�_���O=biԢ��J�M��M���)�U���Ϡ8sS�O��{�o��� u�1Y�1Z�寕%�2Cʹ����.�"��W����r�i:i�b�
w�N'S���;�Cv�Os�[rb-��JY�B����D1׹Z�=���jl�_Ε�(%u	��+k�a/>O��N��/� p�,Gm����9�	�zV��
�.���p��K<�y�c�����S��봼�@h������V�c��Q��sG̓q#�3�1��A�̀]��B�L*>��EC8.��R#B�ؘ!�h6]�@aT��˗�p�+��тt�Q��y�8�n�Ȣ��R��0X��8��c�|�I/�8G<��>@�%Ad�v�b g\�z1�6�igS��֫���Cg���s�/�D�W�B���7�A-�d�X�0d�G4yI��F/~4�Ϙi��`�_g�!��(����¯{O�w�xlgpc�a�1;�R���b� .%�d��t;|��p檥��3���y`~�n�i����$I��No���~��P�W���=`�F�j�.R���D�'�S@'��x��7���Y��.J)�毜fe<�N�sR-���W:�A �i���K|n�	�2�lE��iq�ק��l�,�\�ĪFk�W�{̤c�ޮe8����0����;�]�<��GD7����ˆq�Q�h�ګ�lT�{ ��v�U.UdyOEhQRZ��,3}���~��[������4�&$Ŧ�w��xl7���mC��OT���_�V0���m�|Tڷ�x�I�d�(�Cq�y��j��6p(�3��m��&��L�Ъ��p����ڳ|8t.�?t,c��K�FO�z�7Sc�	�>B����}�����_���C��}P����~�R��x�=<���zWײ]=v1�=��! ^�φt=y0s �D��2�)
��f��ht�s���|��+D�@$�>8�����	>�dkx֟ϤL=���~�Q�ި�315�$|g�*Kr��D�w]�l��@�-X�A�0ǖ�	r��)\&3L�Q��D�# I�K�����J9���%�acx�%�-���l�h�׈4A{7eCr��gh�{@��Ķ��&��P�Gm^��9!:�@:��eb�$����;F8ӿ� ZyE"����2J�[�rDG�J!N����P��UO{��P��SCo�w.a�A��|�/1�8�pY싧�=J��x���.��� ��~�R`�ѡ�_e�N�C�i}3om}H�`1�Tz;��w,4	I�Ѿv�3�M�(����ۗ�5Jv
�[���X���V�כ�s}N���eG�p���ـ�&$m(�?#��{t��e,�:f��O��}]�x��p��3��'��}����O"���JH�Sh `;�d�b~g����Y� �� M����uf,Ւ{�?��=�8ɞħ-�t����J��]>!rڀk�^SQ�J:Y����Ԑ��gxє�g^ddHt�������eYj-�;r�a�^�P^���}�*���J���h{�SDn}n�/;[K�Y���`x���8K
��������թD3�X���5�9�t1S��[3{p(-�n���x���T���
q��P��?;q<u��,���U��5r(���͋�1�EsȀY�g��j������1�etB��I��e�u]��јz�T�)	�n8C$g���A{A��H![sS�_~:3rZ谶�c��}�2��7'���X��Nǳ��{�����
�9T*\��ګ$������\�Ee����J��-����8����K�M��ؓ����B��{V[i���',�hɗݣ�Cl�V����KJ�f��U� 7�K�����d�d>:�v2��'F&ԋ|���c�c��'����
SQ\��01 ��}�n��A�-yo��SG 6����K���H�Nu����!�AnQ�{O�l�����D ! v};&����۵��I ��8� ���%3�-�:s��?�*�c~�k�XBL��.D����>?���0?;w3�`|A��SWεrt���8���n��!村�B�;^^�w�	ˢ
�2r���#vi�G�`��Q9C敮#��BRk�1�;d�S#�<� $Jͨ��-�����ؤ]Q�D�L���#;,JJ
p��O��/?;xz��}W��=ySvVE�2+A+�_��?<�":�<�a��Ds�����'T�DVer�f�|�o�W��l�<s�K���,@��l��c�ɩ}Y�ۉ��~5��ﲉ����P�u�x�c@[6ih�%�tஇ�ִ.�F&�Z0O���ps;rsҬ�� 6b*2;�e����"<e�n��V�]��<rC�lJ����3G��Cє�_J*��<���%��"�P*�G�V�Y�Lt�"�w<'�� �
�J� fg}��������p	S�'��s�=�rh ���]��5H���Ѥ�X�/%6�m���/�I{���*(���軇细�c�ϰ#=��-�2�H��/�ޣ��A9���J�6;2֐ԒW8u�N��in�x�`��b��zFК�:��ڧ$�-��qSn�b���4 �9	h�rc�1��I�)�h� ��!��)��LB�	-�8+xa�>���y�����*[���tʖe.i����w�o_j8h�EgA�FX�]�[+O��bWdq���l3���*|Xl?���,�%�9S�E�E�b�50}��~3��B�����@ �z� WAc��G���[/Ud�>��b1ڃ���s/"-I@���1���χq9��;F���q�|C��(���o�%�~{Ո{����VY�	w e
��1{�O�B;r~��3�J�	*	@�L+����{x����is̉*�x��8�R;H%��b���0g��F��@�rf��o��1ҟIx�+�m���u��#��s!v���2^vU*�?Ǵ�{$ͱ���\1��ئ'd��ž��R!�����ދ]����1���WWc�%�.fOm��Wt)�
"��H<�#\�����-��<�z��^��d Y����ݻw�W"O�ċR�2�����@��.[���9~:�,wܚ{*d��G��K�,���#aS���V�?V�@��_�����I��Ƙx(-���x;c�/J�n������ڌ~�GF�T��A��`_��\�� ��K�}��3:���!��E9���l/��UL�S�X%[�K��_{o��*%�~�bL$��3��k*����=�����Ù��('8ސ. �_�c�;w�J��"�\�v3*ȇ�"�ca�vP&�o�42�$��{:QcZ=
�շ�v�&m�v����r�� wm8����TMڠ��c�(Jc���'��>�W��{U�`�7����t�b�%����̙���w�bX�q���s�U��mA���E����ŏ����M��� 6:F�)�;��ģL.k��+~Z��^*y�Ib��=�q�t:��y��ls�*�O&�h�L�������$n�ñ� ���N��>'m65��]���E��'�G��'l6M$r�
���'. �k>�Tq���S%�>v_���k��n�/Z��s�r����J����a�Ί$nn]H]�;>}��^-$�b�@�+���y-N&��` �`E5�ES��~���Ӡ������qؖ@��DYE����+=xo�sf�0LnQ�X�UG7'�n%�S{�Lm���3N�|��Iu0>�3�v�u�,)��Y[ג|��=CPH���&�p���QY��	�8j�7"����Y��I��v|{pЈ1�9����f��9P�v���H'X�.��S��'ڿ�D�ߐ9��Q������ ��%� �z�����ٽ��e�)��^�X)�����E��w��*�2��	T����=�¢����F뱏�������O-m�A���G�_g��?L��]e�Fx�	�����c�����IР��Wq�HŴn���)c�	�ϧ$�%��HcD 	�&�;Uf�qCPf��=��DNhg�Ro̚_���V��l;�v�sF:0w�����W�j��Hdt ��$�8�~�����'fpJrV�u�PÞ�����w_�"N�Ӱ��$b�wL�Ww��ud8�����$�]��*�(��<��`+���m���<���	� /����\��f�´|�pW(q�:1܃��64tq�C�:�F��:Ż�� �J��+��"��Y�!�чn�rq�#Ǹ�����y5z�������os\�}��ːqd����!r�V���]���M�X2טE��P	ḫ��W��Ҥ[/-S?!b�5��mk��4����r�k��W��6j�!no��:e��ҠꚭD& f�����O�u�$��YiCc!䧆�f({�r̪N��b�	�r�T��~ �J�']2B$����Ju�p���b�D��g��q�1�h˴����A�͍�r����RD,�'���y�l�� ��Jn����gg�_K7S�����Ytm�O"GPڵS��C"|� �V�ɷ�5���^���"u�v���r� ��ᶳD)5\}m�w�q!�=�}H\��g�Z�S��C����L'T�.���"��k�i��֟:ʻ�y�u����HTww�(og:����GO�|���~]��j�����1N���m�,1������q��\���zR�*T�*�x��I��2>���f��	��o&6��q,��r�}����]=.�O9\;k�5��a	F6H��1�s�(��׆��&/ ��9�j���N�$�F�a�?�=잽��L/����o�RCv������ً՚�ꅉ�
2���Θf��R�!�y�OvM#�A��R)�	�7Z��ձ�&��d�;��x�#�̘	E�W����L-y�E�b:�߹���@��N�e&!���N�E`��$�WI
YO�OL�#����D۝Noq���� 3���G~����X8T��3B''��R��$�㴣n�q����4oC����l�
kef^9H��)
N6�.�$�m`��M9=j�8�����Sc�q�C������O՛^[y
�|�L�˥��6@f"�'"Ҍ��s���)e\~'9���ԣ��n�Y|�z���e{j�)>&��<�;�M+�ˡ�j>��
�Χ�?̪�uz������~�>1��N>�0��8$e���K|�@'�Aj;���8��B�m�g���G_�?�����ֽ�7�����n���*9�g,�*�8��#L=s9����
pV��߹�"Ż��9cPLZ�����^+rF�e��/�A����!v��f����`{����!�5ܧ�&w�'��%�9��ah��c��>u?�%����ch_��4����W�1�_���P����}2ej�/{^TM���+	tX�8�߶��]�1�=�2W��c�r&�}�O!%#/0S�W<a��bPx 1;�W�ȯB�47|�r�!h���z#I+4o�l�8}�+RG�`HJ���a��Mw>�\6g�t���  ̶E����*Ft07FU`�B�� A�07_c�2-������M���O���-������\�{�"���LV��5,����um	��n�)��z*�3�ƕ"�t���{����D�+]�@�D��Q�ooˤ�S��J'�a0,�W�*�]���ŀ0�X`����|�UU�x��ܑfKbLf
Do�Aze�qH�0��ǡ�a�X��F�Y�����MϽs�\�i�ǉ$Y�����5���LN���<l�}mP�`�9�������F��a�����ER�<����|����E.z�Z�a����;'`w�j\�Ȗxaǒ�Z��3z�"�d����,Ő3ځ,��@�T^�/黧jƳT�7��G�_IDF�՝����(f̋���`�8T};E@Z����n�}+r1���z,�%�{�9�	$��0T�R�
3%��n��Me;ww!�����Et�B�x�����/L+�5� �(ή�.?�.�2m�k��~����[ZR-c�i$3#�6Q	 w�)�I�4p�κ,��#h�P��_�_�)�}q�D����x��@�-�3����O-f�/6���U1���ʍ�}�!����z��2�գո���:�U�8��
�}��j���Wh�ᇛ�6��ݢ���@�����a���"�X}[����q�&c�,(�D�t�0�>��ӪRl��ݩ�3���y��M�Z)�����������=�Y�]�l�Q�9�1��@�g+���ս���L�BOW�.K%j�1?3^�T>\��r�x��g�z����4�нjg}ڪ�j)�/��gD�����XOt��($��w ��a��_©����,�0]�&��)�"V3������-�N�{�j	�<z�ܙ(�iEͿH*��kf��$����ċ�����)�j�����<�U��f	�v���u��]6d�㤿�q7��P���� ��_eQ���ı��Y�j��NŁOx����(Q(��SI�F���B
H_ȆPEw�����A�am�<�o���v7[����:w���,�ۖ�p��1������(6�Iw�
�]�'f^�S�ɠ���:oQRJ��ӇQ3�.���7}��A����Nu���C�Y��e�O�z��W��Sw�,,N��'H'�ݴmn�:�r׃w7�j���Z���ؓ��r�pq����MaH3�qd���4�E��Wf?��C�K���ˉ���艽F����7��h�[��2f'4�D�,H������aYc�#�+�-'*߾}�,���D���f�3+�@�=i����*��dm�8���d��qE�����P2����X�~9KN�-�����$뇊d��ʀ�C�Ex#��xmz�9��ҥL�����Pb��:Օ?�a�G�uV�&(��`%�����lF�,�ύfO2�טx�#����(�G2�$ܷ!��d搥���X3E=��~vd�%=d�"'k������?C��Ҩ$�Gu��fÐ}�x��,6��+�[#�g�<�L�(���5����y_KE@	1	��ݘfJ�ā�&w+����	��# �>�!y��
3��e�B���U��%X}CNp���!�o��Q�u����?իN�� ^��c��;*��3!u�d���A�~�������aU|,f���;}��H�J�'q�F2����@	��=k��o+� �i����88<Ɛf_����	eC�뿮)�zvZ��	�v�'�$�fU�&HY�h[6�fE�ۛIdn�����|`46.�9�1�M�H��C2jP��j�_��v-��1��u�j����uŶ9�Z�03A�'��p �i8����Rp1�hv�V\z�ۙ�0����^S�u[�l���?(�p�=��C	������pEV�/Ѡ-v:�����
�m�$,�G���׻����_|b��t��t�_5/W�8ezh=���	��H#8��>�jTY�zn:}T�G��:!Z�d%^��i�"�j�8N�G��sxy3�i%6O�t�J'i�u.�4�\S��.u�V��3-5��NCw��L��<��3.e���v}�>���>�p0�}|�Mq�|L�Mw��sHޜ����i4�fԕ��؟M'�G�[&@x��N���X���3�Q���C*d�T+&v���ʱ&@�u����k`���	UQ�m�vG�ޖ���V������U�<h~_����)P�􆃴ۆ`��'D�KY����3�8�1x�=�U�0�$WBȵ�IG��E\~�;�����X�(X�^ဴUռ�����	a:w��mo|���w4�����"c!^(�-2�wL� ��w��ϛN� MqAY�`76ʽ"-x����
�Ľl�;����L���D��f](h��t\Z͐!h�	�>^U.���x
Gϡ;�a��U�[nt
0^l̔�׫��5�	�R���~����.���x\��f@�!�!�G�h��F�j�R�Z��!v%M���N�������m|�U�ʑ*��3Sx�[�KN����sXY��Xy�.vL�ת��&#�@:u��VF�W%/�&_�)<�ǎ�˞&#S}��,I���䠰�%-7P��!2��NbjS�6Z�ӣ� ٱhů����,s뙲zTg�v�}M�0�O~�}����Ӭ�X�� ��ڙ���J,��d�]�0oҮj��L_-_�pd&�SO���值�XY"\�t�(�Ơ{�|���4F��\�%����0��el�v1Q0�4�^���S,�ތ���+��nK�4��J¬X!�+T(���L��O���W�_�}
<��j|�_HP�,�\Y�{�5GJC�!�1�I�B��+h?�������?؁L���x���Rw�|��[���a�Z#:̍�7�eY�&�smbZm�\��v��B�[�a2�	K�3�O�|3��ϣ�$������N���� {/X��Q�� ��l��5p�U�΂D^�vv��ͿD��i v:%�?Q�F{�g�ՠ�`�;+2@���.��{�_����y�g��=���ݻ���w]��S����u�<����b�#ePJ�y�b�Z�CG�?"w$wtZ��<L
���p+�S��>,[�~mrď���xB��v��	��L�Xil3Z^�t�<�h�Q8yi���q�1_�����D��6q�
��+���;��y s�k��s36�[`����.9�.���,���L�1��F��e:�!
��B�N>�4F���K`Vec�v�*�6������}1��5H9�耓?�G�4�+��vj���w�S�c��MѠ�*f�SXg���_VT.G�d&���j������S��S�'�xyͲ�i�NJ�Uׅ�D<#�F.z�.7��F�q�\��M�B��+V�W_��/��|�~��U���7���a|�[�(Ϯr���y��&$�Ę���7�˧C�)_^�=}4[RP��v��WS����m��* d�j`¥�}�i%ഞ��r�cA1��օM�˴�'�Cs��<f@�d﷮�Y�6&�oUMu��TbfǺGΎH~ �H�~�V�ˍܟ�M�TO�5�@E�e�O��A 4D�C=Nyi��B�y�@g?<<���pb������b��%��4ի��I�~)-�|;��T�;��L�-����\�0�z[��Y��K�+U�x��g�M��.^���&'���)�?��������U������G����M�9+�pR,��JJLdyU���۲�H	�LZ���f����U����X��;�g=w��d�5F"R�%ɺl�D')��
��ugH�MCg���;�;Z6�#dt/�Ea��>��i� �v��x�HLqu6��0"Nb�Q�w��i#�S�s��+��d�g8+�(L� j�O�����!�Ҙ	��A3�}1hz�ŷ���`Y��\Ȟo�#xÛoس��MO	�n�Z7z�J�[�{�jA]��	��k�&B�Z��6l�|��;�Xź�" ew w:��7�o���v����\Z�ùY`���S���h��F�liP�@d�t��SG��.I�>���A!��(*5} ��b��<��ql���3���Ć�7�Rթ����M�w.��!�22S����~�Tm�F�q��w��,�u�I=�G��S��c��SArD�TE�my�ug�M����y�#}Q�$~�U�0�ۡ�5�E��Є��� ~�"�jL�iF]��m����v�OҴK ���N`b�7�ޮ�c��:��h}�����1�T���hժ�~�]2��]��h0�;)���l>6yx�8���+��U�JX����f��+JSɁ�`R9v*����	9~վ�o��?J4��8���sVI�\�����ᆋ�(�;� BxT�|z��?��T�)u��BoL\Ҫfl+�~I��s�٣�P?I�����6-j7O:��	��	�[#�ع6��9v�E��*l��!�����L�jgD�m'�1����kWEk]a��L{z���Ezbj�P�{��y�U���n�d�t��뀏���ur���Xg�> �Ȣ��t��� j`����s���s�~�s����e�g��?���{��ë��#(�'�&Qd� �Md�Lۊ�P:���d?��7^����ҏi�pQm�{4����O�i� ��l~]�}>��ք;�h�q.�qK�Z�=�X0����)�Ô��1�'I�ho�%��a�}�i�.g�?qN7�~�-�\w�mʎ���S�߈�&Y��i=�y2�ڷ<����H0}�Ny�?��d|�|WЊgSD!������Pnȵ֒��A�s]�s��ȉ�?�B�Y�zsF	�P*�w�U�ud=w���Չ�.Y�:�i9C������>7-�	|�x&@7���׮!��l`<)�(��ǞHک�'�b��C� �j1�z:V�RL��B��օU��;�6ME��n}��0������&��E6*o���Oמc���As�r!j%��>ƹ�޷"��q��i��2���:Q%Ym�!<{��]�k)��7hn.��/#6&�J���v��t��h��W�:]���,@�/������+���d���mJk�[G$>��cD<��mw^���m�QP���+��<�	y%���%Ы��>��B{8Vc��f)фdj��3L���ԏ�������?ʱ�l@�gj(�z� �@f��	��m��03ڶ�H��!��ߢ.hF�`X�k�We��!J�L`�c��ݳ�'��M���z�T��c�D�u�VcڇnX0��\��ٯ��f̝ӿ-#[�dT	�^�j��*)A���m�¾L��x��������mХ�������j
�,�e�4��5�~a�ƒ�u��jߗ��@y�2��L���;>��M��<�>4p�͐H���:��#�u���S��/Ѥ������oE�H��J2��w�䌹�3�������C�`��$�P�rb���}!��s�=�����!]��|�^9|O~����J��X��,�@˿��a�?�BM�Q���QT�����8#]#���Y�9�Z_�z���5�3�4�q�*�N�k���״6���0v�~�I���WZ�����ֿ����H����r�A	� ;W�W+Q���Υ@���WH�W�H�%�o���ԟb�_^�&�l9�\��nH�:�K��o�:@�d����"�T-^�����L@��I�Џ�yp�Wi;�`����D�zD1:=�뻨��0�P]��2;ۻ�a%�����3�x�y�AѴ˹��]��\���t���V���� b��N�:ΆtE�����(DA`υg���lИ�6�{y��H6�/`�JuS&}���#L�y���E�Fw-�CN}�Y5�Å@Ք���7�WM����4=�]i���w�j$}04g�u�`��*�Z�!�D4L�6�3m�������$?���=�Է�h5V����9�iY=g�T.�=�2r\&�j��y��'��^_i������;�1���tjIL���T6�.`>Oŝ��x������!<�4����Z�8�}�JT�t2�{��Z���l6O�Y�՘4�,��Ywk1�ކ�)��oN'T��}�l'Ҏ6	�T���l�R^��� ؍�Bv�"����������zI#_8R2_<���D���Z��)B�����`f����"8x�R���Q��O_fQ����*��Sś԰����}�h�>xS�+YR���Ѣ���~:�'�I��s�4�_U���������UE�X�ĥ3oP���q�oa��r����/Ŋ����E=]S�яߣ�w�{]5��o4������.>�?�6p�18�9�������C9��
���+pCYb��G|H,�g�Cɗ���>b�3���v�L�c�ƻ}�U.b��U#9��^/�޳�����"�Jq��� H�P����U�n�SܟMN6/�${�|;P��s����X�KR�J�7y�涂P>M���`%7rM��!e�S(aG�)����nBi������SaO�-U)M%��6�z��!�g]���Z]�$����c��M���gBVT��EŞ���j.S��������a�ꁳq�.H8��B�6�?�"�;)�;�{{���jsB4W��L��p��:Q�Kw´O�@xy?b�vK7h��Ƣ�a��I����B�^�;�o���Q��2J�L���JM�R�ˉ���h��"��΁,�"�n�N��9lM�8��J\΃"b���"J��Š~���O�(��)V:Md�$��e�*il_w�z-�=���t�IN"X�B|K�dUg�X6!! �W�E	� ';�+��g�qd�g�fv��A� /�]vA����;9RҌ��R�ND8��g��.���6�m��/�	��=�X�K@��]y�����ᘲ\e��)�����є�og=Y6�����Ǔf���(*��e��N�.�QO�9]�#��p���1˜��A�d]fgW��p�������h@�xh�[%�r(�cC����Q	��A�L5Z�~󲆿��%�'�$�,:C�Ě���`p-�m��L��f�	�6q�����7�չ���@�	���+�Vv�b"H��<l�TR�Y��T���2伆�}��l%gX7Ж�4�C�x�� ��a���[�4k�W�R�0�5zt�Doa�@���K�I�k����3���;O�dj�=M͠��i��j�r�R	.�f�:�@��Ȉs���������"�lD���RN�i� ���B֕mX%�f�Y�;k��Q��_��d�f��W��}4��i�
<%�IA�p�"��)$+��m�;ӲW��l>��.�Cィ�����S����͂'�RXN��ƿ�����R��"�`���[a������
Ωӧ	���A�gO9�L���ºQ-�&��[�U}.N��@Eȉ�@5����l/Z\���x_ͳ��p�"ƴ��֙Gr��!T��S-ЁʋفlÁ�E��iյ����V0ud5^��d�ǔ3@ހ��5����aJ��(���%b��g���iC���(�0z>�]7iV>�s���.����݊���M���j����"��A�k����L��~���2[�RL���˩��S�8��"�����¿'
w�
B�%d�n�DA����V��u�t�wN'G\PT'7�=�X�ZV�f�`��/+g���ԅ����s��ˠ��t�p���v8V��|��>���o�0�漚�
�sWEc��xa-=��aײ���~I�(�=���!N�+TS&{�*t��Qĥ��	�7C�~�g�.�w�{�8+�5��w�y�l�_�r!�����{��Y%/� |]�q����.I`�Ny@�f�ǽ.W�ra�܁�9eQ���+"�s?�ׅ6F����CA[�ſ�9�;�Ɛt	��r��:T�J����nP����P���t���2[���n,�$n@��\�A;�a��}��];�T�kb����Җ�;�l	Ԭ@m��ix�qI K�/��
��/�S/��g�A��D�
�s˟�;A�.�ꇴ�@Ն?������m�{Chh�;m�+�J����ʘoǅ��Ċ{�p�I٘�i��A�ۚ�F�ť�dO��5v��3m�]aTg��1�V5`�r�3�MR]�����M�d�~,N�S.�[z�|������f�T����G�EIg&���go^�l0�����I��[�p-r&����5:���s�x^��u��"<Ri�=�@m3#����IwQ�>#��;�w4p=Z���?)[r
a
� ��]�	��q�OF�h^{�������*]����\�����J௠��p�$6I曅W�k����K8ј�5\��_0?rE:��̌�R��i
�
���oz�^�Ŗ/
�_��zg���d�?�]�����:��?�����ñf�Q��jO�6�΂�E��-5����b���l7�N���l(c%���	�d��������ZxA�\�ϛ%��-���N�Y�����m�&o�6��Z���I�J��� :|ok�#E4'�u7�Gl�Q��;`����Nv�m1#��*�",�Y�#k����z^��^ȗ6��E��$U���.>jm�1Ŗ���]L���iY�F�&v(�
�ɥr����:��9r����K?x,ʍ�qdߤFG;{\���gT@A>
��A��Ϛ�e{��Rj��~}�9� u���
<�Pq$���l��ԝ�7cQ���@da Ź�!8Ai��Һ¹��M |���D��q+�g�Ɂ�,�U�Y��lX�sܲn-��e�E
�+,�`�8mb�l�Z��ֆ��X}:ix2���33�kn?��/���D��T��pv^�JŒ��$�{Ӭ����W�����V����hF1�u�ukD�`Js�E�=j�1Е|�)��k��oq
ݹ4��y�}9�ab�U�a���&&��k�x�I���E�LX9d*�w�I�B�|#ʅ��C	 �Kz�Ծ�`�T�yR�up��~�El�L;1^;���	y�[(F�l�����]uYES^Ƚ�eS��z3(���]�f��4�y���qH�>���$ɶQz�}����\�a$y7������C�_�9HV 됟\>m�%'�'|�S�H�J�P!L��ãc�E-ӫ�Ԩ�;�膘6�K��+�n��S7�LĆ����%ˤA���D�ozt	��9�j=��z�e3�)���a���i�d>�dS�F��s���fr��"7%X����E��d7V+����#ϕBdЭfA1\�	���@�>ŋB�K�.�oX$-��S�a�#��'�7Ɣ:�2��o��r�B��r�6�b�>~W�w-����lR�C�.m.�I~7A0=��i�Պ��>tLP��ND�3��X��#:�9,d{Rc��lxPۑ'O8�xY`��K���yִ��mY�w{L�=�?X-)
���E�����T&��I�!�e΁��|����:��T��%�KX١��~X����t�m�³��"�/IE��E�#�s�P�ΐ9J��"-nʋ�j��Z���s�����8����!ٰWN^$o	����0>D`����H�ؐ�fQ����(+���iu��6�VI)|y�*aݖ|�ȹ�ۈ QLX��1*?��Oɪ�:�ww��ҁ;��b�#��9! �D�%���b5K�ݹ0.�ґЍ2�5xK��5  x��kdV��֛�=O|3(�J����Q�|���j����,�2����k������?�;SIb�O��`�L�k�����e� yR�z���V9�G�P�K�(W'M	#n�1�lW���Uy8P/C4a�����Ex@*M�K�Fag%ig���\��4�B�l�Av���f���xq�1^΋J��h6O��ް�a�JX�F8Ⲣ�̺�m��;؁l�Vg��s���إ�⃀_��K���|�y?q^n���2[E�o_dC��q����~}�ԯd�Π��ˢ���DR��R-%&�?�a�>��6Q��{�Q���kK�E���O��gm*�T#�)�)�ـ�(�z���z����m�}���T���o��*/m���!�o1)��Ә���Ĩ��� P*"��$�0�E7آs�]�I�k�z[��Gk 3o�4�����>�K�� ���}�3�{�>-$�+7���	0�����u"�JTxqk�gYf���ruΒ�|&Уhq���<�Z�\^J/2�s��J���Bpf��j�@�8Z%j6v=�E��\w���'lu�\���^��@�"�ˈ%jmN�P��؋&���������M�=$ʫ ��pd;�kQ'!a��JZ���U��:�P�������~�~݌Q�NLS'�)Zc)�3��������}^/��#�v�4}�x�n�8K�}UP�&��e�N�{w�xA���bj���0n<�+	�l��
Rfo�k�NMNgs�4)Mr�+-��K����I��HS9>�@GT3�V»Td���Ns�0�=�b�
�'�����fc����k�7��0�����g�x�^�C�{�������4\�K��q�P��ھ�$��9�~a�b!��y��ё@T6BFt��1�t�lǠk������+-�8�����g��{���n���-���A����{'�Ei3�B{�������!I��2�t�s�M��d���ʍ���/�k�Xt�؝�F��O3�)�F]���$�P��L�� )�Tv��莆���M�vP7L:X=%��K-i�*�����h���W�l{SW�+��Ui��x6wyqd]8rˢt��z��g]+1�w�#=��܅DgL��?�9S��叡�0�B�\�f_y�IL����VR��t��@ ��C���(]��.���x�^�'��XH�`�� ����ɶ����=&F:�D���߂���-f���=�+���qܵr��G,Ѽ���}�%R�~��n�&{��R h������5A�����j q�~u} ��4�g���$h��e���K��+�e
H%��\K�/�Hޒ�ı�2I�ȏ�c"0-��hq�s�,{&B�3�Bf�M�l=��۬�T�Y��ӈ\^���.V����7�.��ʵW������Q�4�#��"\�X u+��o"mu1;��V�KNQB�+Jf��ay8{���,:r-uo�SA�ô��x}����[v�׭��������|iac^���w�7��FFM��ToZ�VQx�i��v�,	;�LQ��N����Y�1�N�����F]G�	AB�z�5�i5r��@�!��g �H��x�w��Ι �cQ�`Ȑ���wn�A��+��|��}�M�y�[d���Z3쫧4����*�yl�0l����)U*���?�3@���vЈy����S�ok�.)��u�����'�m7ؿY'�2�y���rmވ�dxH��K"d�ŤX�F�?�̴<��XoS=�v㵤W�Zt��`�����u!T����1�[���P�����wU~)m��}ǈV@�JwMJy����vo��\�i{���h�����>do"�'�����/�n�N¡��E��M|\@p ��^��C[��i��>���zCr�D��Y-U�A�0R:�+ς�/lϪ_��C�V�~��3/��)�Ѩńl:��+�2�B����uo��n��%+�YDw��%�a����6�i�":�g� &ӂ���=`��	#��:��<�1�!Y��+<�����h��յ'"Q�(�D��O�����u�q�F#t���(�#�3	�e�$h���V�thc���ꪬ�&aڵ��"��(�j�IO�����.��No��>�`I�DP�MF�kқ(�j2��^��, R��p3�8�|��� ��=���<���[`K�A��݉
����XPa&,��!�j\��ўR�Q'&�E#���V�jq��/L82��������6؋UN�?��),��	�aw��ɛ>���2&������S�9���
dkg2�[�_�,PE�N�rz�X����L,���v����Z'�>���f9�eb?��f�o�n�K���?.����B�m������MsJ��|�X���g��'�C����a��ۗ�V�%�hm�[��<��:[�� �$����������B�
~u���+6��|�>Q��>QDOK�b��=��$n{L$x�a����bp1��Q��jpf�}Q�Nƭd�J	�U�F4Y����jO�`��1/a[�*�V�1����h�x"���.6���I��Ĳ:,�{�#�{�Z�Ŵ�d,�~�]i�*��:�wƬ=>��? ��q��l>���K]���^������Ց|�L�J�q��}V��,��Qq>Å�;�x�D��]i{m�װ]���n�� �hS�a���d	�eU��`nS��u�fs�e:�bxp����ph��9�U³{�'#��a�*�	��P"�`V��p�	cʔ�IM堦}�D�Ǘ}��1�6Ǣ��͂�
\h+���7? �$��Ԇ�Q�ڍ�iC~��oۃ.�.�S]|�hh��'�f���H�T���=�4���H��';�0���Y��\����~�=�FZ�N4�y��m���{ftTB[O�GN�2��S ���������)gťί?\J��N�
�rg������T������c��|��)K�� �|~x 9\��"*<���7
��2�] �ð�2~]g��|�?h��9E�����[H��" ������!<���Q|�U��`�i��цO�\��t��&�% ��q��6�I�U����c=y��i����Kb��+����8{_��<���s����g�fg�������Iv�xJ�ȁM�E�X�-�=���,���[�t�_Y+ � ��TweF-�v�Q��bv�	 `��wd�m��0����b�!���Lw8�����%��	��]��[��4�~�7w5��j[R{�#Z���*"�Mz5
m�^�Q8Ss���� z���9׉$�M}R4��5�4T*0�,{��Q�g"����{Y�m,fO����s
�[������$k0M�n�	�@堷���;8�Ҵ��.8�|�/6w
&������j�����2>V0����|D5Էm���>{�s%JQ���i{)��h6d�s�h�-��"iG���ѿ�iI���4�}({�3�>Wu9����bإ\���FF�6I��+�GU/8`��z$C4�d�(U�V_�ERKs�������D��>��TߚԖ���{"��s
Xq�X�{����20��V����S�`O���Q`}��:q�K�䐺�!.�,3�s���sF��h�a	��\D�)$��� Uq��L1@,�AR�r8��L"Ȏ����(/�xr�0��w��G���������[#�T]ҽt������3=�0o]/��¨R���6����C�W���ج��{`���:���d�!�#fጁ�Ø#�a����/�1���
�AQ1���6�%��^�k���¨�?4Npb�z�f�r�$g�o����La���fax�F���@n��Ig�~�؁u��o��E4HM�b�����Ү}M%(���?����Ԑ��-��VPҦ�.yq�����4f:^�$󗀖�꿴�
�ö�"b���-��NP�/8G�FW�J��4B�ȫ�_!���ɒS
��L�ؙ G�X�6�Qbֳ�U<�iy��'����:�~EN,�������}"�l��k�I"���>>@�:�`�	�1��^�w�H.���{{2���z�?=\�!���anF�߲��`�^m9/��u�^2j!,4�lU�>��\�q78�>F�}n�%_�/͡� ���eO��\Lp��B��@ �q��1�`9��K���m����ʖd�eɀ���2��f!�w[Ϟ��㶬��_YȊ�ݐℓ~�չ� m�^3�e�V��-�4d�	��P�6'���8����7K3�o��*q3�i4��Y5'�aP��;phwY��i�Z��G��^2ҧ= ���沬�\������U��6~>MڪL��v�8I�	N�cv����J�JH�Y+��X�	;H�@��y�`^Z��1�o�5�0G�P5קM��l�&��.<#nBn�I����v"!@�2�L��������J-�Ӆ����9>43ܾ�loZ�/��kcǢ�3�yA�4'����Զ�/m'��ǺS�5ޟ���:Tͨ�P��YVm"���+��^U��"%']��h t]p��S&�089����L�����tnDu�I�h���nQw3[�Q���`}�B���Q�2�U`�l?�V	0cᳶϡ�Y�5'��[) ��M��އ`	���[�zK��c�S�zx���tЂ�	E�x�J�&�QɖUY����6����.�Kc�l$��U���!&=���%3@���8t3���	ev��Rk��)��[��jH��lo 1�A�v�^ł��N��(���͵��CTs����aCD����!�Zp��e�]Ž����ݹ�wx^�"��@�܍�v�aV��`��yJ'a�2�{d	Ł�:O�8�3�]�n�ׯÙP�DٿJ����B����c��g��r�*n�^�Q���؁�R&^j�	��J�G��B�9����B��������YҬ�Y�X��ŗ@�b���������!'���l�~�LY�SآV��B6)4X�t�sP�oZN���y�����<��C�� �nSD�tq;l尦�*���d�n#7p��#2�W�n��+N'��}mnZ���r��^��hΣS�2��:���V��mvD�E�����c}E�x(=���F�m���l��hbb�r�*ǔ􏕀m|?1� ��xN�2:��ě/����e�w��Ҧs���"�>�C�GE�q���Eo�ӗ�����C��3���\���1S^GT�Q���$ݐ�G����J�^�J����,%p|@'+ O�x���{�����ʳ(nCKN*lڍ���7�&o�֑ՙ��3�U��"�b�"ǲ��ǐ0��k����V^js,�Ͻm��6�hj5|����PF�h�KK
t]���ۛ�`K���JIt�}F����gtG�����b,�������\��g��y0I	�Y���Y��@B�:����}t37�N��ͪ�N,�[�x�>i����P&\�?��t{����VY@���ha�a�=���ڼ�i�Ʀ�ݮd�h��sPw>�����1���J�)�]�R�"�2�a�aΙf�Jab�c��IhR��};��N:��n����	$��G0�X�g�u=�� �I����fȔ�z�^���3��᳨Uq8�����p�b���w�;���/Z��ZUB�p�5l���u���Fv�V��/7�u�LA'���Ƈ�����W�
(����d;�-E��e�=Mv������Ib���?�����ml�+�]w�=��%d��F�hg�f�uexm!�L�
(|Qo����)�t�
;կ!���^��D_J�!�����z�s[����*8&t�Ԏ��5v?>�fS�[��f"���Dp��{�LG�-0�!�m���Qqq��>z7m�Dm/��6�߼^��P��<s�!�q��˕��z�$%g
H����a)�m܅	Br�W�z��O��~�����bC�h��TI9,��" ����'Qf<�[���W/:G>���g=sza��%�R$��'!����@qN�����~9��KE��Lo5� ƈ��G�qc��Ё��\���w� 0)ڞA^�E���R�6�T�s��'2��̂ ��15e��W��z������8��]�&�w��i"� �z*\V:�����֦�_��3��9\���%������nRb��ϓ���N_pc���jSR�0\_�	N�whꯙ�"���mզ�
�;i���~x#�b�Ȩ�v�E�b�(R�T���1�4L\Ed��+�,%V_�f�k��.����t�a�O�I�rه��񲇥��u�u�پ��C_�J�7�����E�q j�~����,�P�4Џ���8R������)�R���d��=M�6��{�`���$�T��<$4/s�@�_��\�I	��װ f2x�t����!�
/Ч ���@{��q���#ͤn������m-g�o�`1���<x�z������4�z�Y�h����IR��f/^�:�,�=�6��c:��6��s���Az���vl24���*X<�!&BBclT�)��6��6� �Z����X��]�K�O�$ci*-��`�w>��&��B���[��9��Dd9����� O)��޿�W!i���������:���Z�A龲C��M��#V��K�!�����ݟ�]�BѢ�]��/����//Jm�Q��`��izxt�Y�$�^DK�V��D Cܿ��P.Q�u`*�۬�d�n�j�!���	3OιT�X�~���
s���g�M2N5<�����n��[�XڀLZ���F�hCŋ8	w�ͅf1u�s�e�,N�/݌�FH��R�֭S@�GN�g8�R�����/	Q
H˚��p�*i��g�#��,J7eVC��f�o|���ԻÛ�SZ|�d�����?���#�w��h�8���"�ӳ�@������gj+�U ����!�"�*)R�}����p�t�t�O6�Ʃ�m�I��_d �� z��!1ciڜ
�酭V�(6�]�v4ςt�.�Y�p�sIV%�p�8�� ��6r�
��:~�K��ru4����o�R�m�E�b���g]灅<�gi�*O@1�̗�t�������Q/�3=k�Wo�@BC�ӠM9�|��}u�w�����_0n�}IH��-YN؎�X�u���~�'���sp�H�	�p�K���M,Y�2:��Q��64��l7�C���:�8lõ���)�~фS&�s9�Fs�٦0gC��FE����w�j���<�zC�V'�>��9Q7�:$T [��켶�+&s����ovQӐz��PU�|�?�G;�O<��.$8��
��&8�$�xat�"W��OW�Cπ�P��iˑJm��1JH�������a%,�hӘ��a$�H������^�D_�P:yy�Wॼ7�Y��ǽ�2�͕��Y��� I(��`��k[���=�������i���N�� ���)�]A+�xY��4���h*⤱���N�q�!�d��3�x�BĲ�<M6���rB;hx�X��1X�~�J;��n?�U�B�cւi�?���3�q���^)~+��Xb���"���uY,��KꜺ*��j�4��_�`��qa�D{��l�=�=iD��ju��>�,Ί�?����� vj[�Q!G�6B����9
��q���R�W�PA��0(�H<��I�1+�"ܮ�X�z��k&)fA8��χ���-��#[������Q�N���J(΁4�9l~1������J�'�Bf�HT��S&9�h��و�����M�a��+|L|ʂLN����w̯����Tnz�����3L�F^�%������P���'�Ղ ���T@���i�6�Y�����ٟ0i����gAyVU���'��B���eO�����x]&�&@ ���Lǔ�i�����}��r�
�|F�^kz�b��6J:��uH����w�nǼ�<z���.lH}F��vO��甔���p��u��.�?�X��RԸ��Y:���yU7���U�M�]��HB�*κ|)ӎ�weV��}�sqetG��Qo���Z?m+0�؊)�Vī�[¶�)�A�[����l�8����yD;�}8+s�Zݯ�s^���Խ�]j��Z��z�i]q�Fc�)A-��~�RWˋ���۟������us�&���9����Q{a��x�'V�j� ���i� )d����}&��C�f�B؃�&���
����R�1�Q	���=s����Ɲ:JvdYR�$����Q5�-�n��/���:�P��/=����r��E��t�������C���y�B�&���$Ԅ\��9_Z_�k��y�R$U�",�����
�D���_,'��
����� �0�7��<��@�y�j��(��c�O��[�����Jo�T-%f8�������dJ� H��B��_hX�I�!����b��o6z��?G�W�+J�@bK�=o5B�v9�=���D�^��FPq�ޗ�J�ʎ0J�:l2�4?J�7�s\�~�т�)B�������{T5j�jV&XP��� @,��y%�^���&ޛr|�Ă��خ������"�����S��5$щP����Ε~mu��T�,�����d&��z)�ɹ��'a�� d����\����AJʱ�vy��c��p�c�N4��c�lF�h�
F�k#<���{7�"�܀Om~�?f;f5��<+����A2�W@(""}=�M��غ��H�Py�tX@g�+[e5��*U�N5��.�L T軞X�n�0=҇��ƈk� [{l��"f �,~�~��BWeRN���u�L�s�� �d+�6L�HOfbdZK.h�ՙ'9�{�q�7ld�!�bƙ�Nї�$G�����T������FzLS#�dI�o�:6,�\A�0����n/ϓb���(�Yjt��v���}}p
e�t��j2B��sd�ހ�ZFQ��Mz���0��p�r;D1�#�³#>�2��NKE�>�g�DRJu؆B�{gakS�͆d��
�mm8F�FOr*(s�>V��: ���6���p�E4�d���w`5RmV��K�p���$)�ӫa4����O�����hi#W(�l0ץ?��T;6�v�6S��}o%�K�leZ����}
T�	�>���OKO`�P�IK��	��-���l_c��)��	��M˱�tĶ��&era_oKc�����؇A���ho-����X�P���Y�&���9o�L����基�/��M��<�a��-SS�@N*�~]�����V�q{��4�����@�1���BL�򩦎�X��q ���v�`�����c)���J{m�Ҩzٛ+�y��a,�U� �bˤ���_GO
o��^��� -�%��"4�4��KOV����&�����\�o�/��M<p�}�S���k���p[�vd��5�ar5��Ž�"�<\�B�E�&F�	�04�7��_V�`ii����y;'�E�
U>n��Q�W_��Hn�mceqA��zjG{lM�t�uXBt�s
E��ڙ���ɽ��;HS�@�ir���_ �F�]�2x�'I�� Ԫc0^�A���j��Mrmr�R��R3�-�;ӿ�u�i������P-�!*+ ��0V �H'P%c����f�^�w����D����\�\yڌ$?LY�"��4"XU�d!r.���)&-������z�������0�,�Ҁ�?�Wa��9�ϫ��s�j�A�`��2�)0#O�����]�s3��e��;k:�N�/Fbe��{��i����|4C�S���eŶ�D����QH��&	u��E�A�y$J�}�%:g��Nm�<p:��B�q��i��������S\C�FVx�tñ橁�p���$N�w�W�s �谏�SẤ�  ��� �04%/�ɄE/��G`|�%7�7m�*N���u�H` H,v��(�J)�T.^�Gr�gq��㒎��M��uC�'�swMZ&4�����p���=�f5���˽~�{�(�����6�^\��
���m�s�/Q��PG_ȌǳE�,l1a���1�z�KJq�5��hN3��6�V�Q�9+�lh�O�I�ኲ�
<x��y�٨�����%-��'��Q�@���ub���غ��v���
xA"�"ъZ/X��\o�Ԙ�����
���*@'hӏʕw����#rp/Ep�s�P-�����N�_��ϗ24����@Y����O4S��TG�-vyL�ܝ�L���������tR���@� Ъ��Z9�CS@M#�����*zs]ִ!�s�(T7�p�a,5ȵ�����*���.��$�^�3P��C�o6�ٜF�n���s�>A��4����Q '�~�m̅˕��.;��	�cͼ0�;�H3�-~!<����w�Y���0�d�)��:�dV	�{��'7��ţ���%��f��Q�5%؈C��fob��U�A�݉G��L�`�G$�"k�2��K. �ljz�M�]��`���}���e/Ƽ�8��1}S��v��%wh˵L��"j�^�4\
��w�8]r/�
XɃ+����z�<�������2T���Gl1�Ӟԃ�P"5��>��,RpXh�5wnO�ۼ��x�s����\���A#'s�f,A��ԛO�B���O�G�e���џb�F��]��������C6,�)�t����Os��}x83)������*��^Ӑt���y�~���i9LF��؆��4AR���)y����Y��Q���7O?=o]��2�2��1	a�>�{�}�
K�W�� �Gx
;X�f�˸5��� ��yX��j#Q� �1�l!cUY���^N/��_���
�F.��v17C+l�xߎ/����Ԙl�`n��Tʲ:V�R^1�ژQ�����S�ڂZ������sx,Ӧ���K�j�WF� ǃ�i��)IDb�e�:�$�?[`�b������AXvg$ne<֕�ԒJR�z?��`v��֞2`@.DU�����$��I7�K���[�����zZ?a*4����S�)ķ���Q��Z؉#߳����i��_�������-}�ٟ>Z=�R"�/�h]*�b�7'������w�9���H�	���c��]ȷ<!~�:�N�V��]Ѿh�~��P2:9//��d~��u�Yوz�QSMF���VS��r���sdОD��Sc�o�'4�BLz�(�ʈ��6��t�;��(���v��"�A==s�� �P�,��`�s��ec�)n�i<����H�I���5��8Ov�I蚗9��"���|��C�+�5&PZ��E$G�f���17��I� HR"�q�9Ay��9����R࣒RR�jsD�P�!�R��2�+��5�D�n���QpSn^�/��Qv��;�f�&����9Ղ��םR'B�q���}[0�{�q�^R�r8\��ӗLd�Y�w�!A�:Q6@�:v]`<���;�Ch.�t��������/�[N~e$`IgX{����uC^e
��������8�[ڷ�����F��\���Ӌ
q�91�������� ��*T�tG�.x��!򬽗:�m�:ћ�L�L4�.�ɍu��=����}�?T�
:u��pQQ�q�� ���Dv���=T �>��S���ܞ0��s1�R���
a�t#�� ���Z�����>chG�T���D�4�e
8g�cR� n>�J�{�]M�w�9����|���!r�s���p*l�7�},�d%B�O��;�o�R��]#ɘ���A;+&�aW�$���3��t��y_KD3�2�= >@�9(]]/-������nhCI{��eqrءeJc!��	�{{=	_�M����$�����d%��9�s�D�y�k���j�W�����M�L@�m��'�{�����y�_mO����[�`�0����s�XrN!��\�z"����l:��3�% ܇�^=��0a"�7��0�]=�qd��j��)�T�������`��z;O�Pe�Z�ǳ�}+x�w��$̗��9�$�wY����2����PT6�kf��rQ���쨩�Tr,�x��>�&G~^m��Ol��J ��hd��.��aNC'�<I���8��a60�/�tl�*F ������v�Hi�|	�2tQ9�Hcu�1�>Wq�y�T��I��S yuyn|�>�{�۽v݉VA�j4+ (<�Q>L(�7#w�,t+6Ш���J�a#�X֚*;)�̥'�+{	x�=�zj���ыN'�=T��kT�T��ڥ�8"ُ�TR���AP)3�J���1`�KE����G%Io��U�_���?T+��pB���Csm�9tt����ot�D=�S���c�k�f(t�8@l��k�r�W�T��CƁ-J�oX"͛������щ��Lި&���҂������Vzf�<;���כ����,e2��Tє��2��䡛��g��1B]���̘MRۓG���UTMH������bm�bV�:�I�* �#��$kNy� BwF[i����Oe}���@E��PUE�b�9Smv0ˉq/ċ'C�	���������*iEu4=�+3���UE�#SY�~ k��}� ��ߑ�3�t dt9��=p���$��0S��3���3� ���\�8]�0UW36õ�i�ek	͠ܔ��\]0)����Wgu��ޝy�b#`�/�g�"��_v�M��b,\p��̨ku컇!���8*�4�V� ���{���SH�c��U���P���$t��������iRf��9(��?Ikk(�8����ם��vޢb/n^%��n �|C���.���������])�H�2��[�vUE4�b7A��:�l�iA1R6�ԾeC��T=����y�~w��ݲ���כ;�~�c��V<�˖ �h�&˛�0���j�	v���`�%��5���K.V6֑�:�Y�z"����2~^�^�e�q,��=G_�$��Bdt{�ཬ��`��iC��2knluw�.-/�qb���������̜(�W��'-�=sEp��t&͑dO�a�h��(5_�4W	��G�{���T!#%~�D�մ.��n�����T�$*����6�-�kz�cO�Bjc�E��=���t  @v�NV�6�x�X�����y�i� ��fJA�U,����JR܏{KAr+���R������?ت��M-�Ҍ|o����&�NNS��5������Ru�M��O8�&9z��Zh�2�8
��\[X�c��8W������t����Vk�Z����'g����	�u��v�ݓ��Z�g+�6e߰c�衆<hɅu�?��y��b�}"_s�q�o5ٿ�@d��֟%�k�~Ѩ��/���s,< Aޮ<0��&�f�|�s�ꂺf��tV`���R�d�񢇢[���{��ǰ3w��;�=�#ʕ9*���.�)��b]�,�9%Y����
�O�dCLpX�(Xq1~�#��}���/�C"�(�d*V�rgN����h�
���l�l^Yr�i~��\����ogiV0�Ŗq͑ω�=p����x�G2.�C�'��j��4dKQAt�G���vy\(_څN?H.`Q�^���}n�d	�l��|��w��K2�\�p�E��m���ᦰM:�`����c���{����oRMOl�sgy^�vI��!wH�_��)yޞK�s���DjX�.�?����q��j�w"*�؈2FeJ�K!�Sҏ �a�]��HuV�g�4[�
@t֠�a��@O�T�	��f�q��-8R�N� �'�f5��ƣ7�l� �u��X|gG_�/��<O����K�|�G?�&��HS�ɿ%�������fKA����5WF6���X�����:5�b��B8s|oޔ��#�
�5�`GY̻=K�xc���R��ꏥQ�>����Y�rv��F��Z�Z����L�z&�# 0��,�ݹ�^ȂG-vq��Q7�g[H|�}�J9����?%H �ρ��� �w<Q�tғ"
^����z�n��7�-�f����^8-�h��i.]��X�Ƚ�ad�g��G
���8rZ?�i)�HZFX���!'؅i�zo�a>�%�v�  �|m���4zܺ�5��p˞��4%�t��cj;�[O������9�����ڞ׳�%�˝`�uҹF|L#�B� z+������.ayZL��Y���J��є�k. �˶i��p|,��yo���c�y��N�z$iF���b:I1�}"�>���Z��j��-��Y��P'���dB�QSZ�r�JҴ�����=\�/g��j�»=�^����fMdc�j+�[�7�h�:���0\ T�>'��7�zN��,z���=3G�����$d�·��&���g%37ҥ�U��D�CZF=���v�v>ԩ^{��z�y@9F[�o��H���z��?��o&�����i�DkF���Q���gQ��=����p��)h�`�O�¢�Qt���4M�Q��}]є'L�F������h�`n�~�m���}خW�܈�x�Ё���fu�C�eg����(~: ��I�s�33*ɶ��@U�JS��u�CRٮFvC�׆���ʵ��}Շ0�PU���a(����Q�U$6awjb�d�����ʐ����$��{-��S��թ?������1RXrS�[<����ߐ�)Gp���.Ξ�Wg�^c9��?	��&�(xcL7���� ����Ѫ�E9w�;D�f�����-Ʊ���`��>./���Cq��L�[2H��X������T�-X����F����n)q��N��A�v��e|GB�h�T�L��qn�Ν�aLa��-5���y�Q5>��,��j���Gz�G�ͽn�I`9�G���~^�׋�@%��fpf��Q�w9<�C�%�*�y�����f��yH�I�(W�可ߋm,6�����[[~��*F�[��7�-I�A�)�i�"�f�
��x�J�z��%�.7�+�}�������g�|)��q/N(xn����1`��Z|K��Sa�%��^��`��GJ�h��+��a����O���&�g������p�|5���j 
V��.d,I��6ut�7~�?�i��^��Nu��D��Ȕ$���哏�f�#����h�CN��f�}c��z N�]+Y�)H� &�g����g�f��	��&c�����������}D��Jq
��\�N�mq6����$�1>]���?IQEI�P�'�Kș�u%E���t�;�
����d�X�U��g?�=��4�TMɟ]��bR�x5B٫����R��*��<=۴���e�m�e�>Ĩnz"�<d�ĩ��W��)=`&E�%�b��*��&(���W���ְ8{�������_�ܲz������$O��1�#��z	��tZ>zT�ܡu(���Ht*q���S����6�n��Ʃ����xDx�#���V>(H�8�a��l_Y˞�Ki�7���h�~y�>�/ <���B��{nt�>�%�@[VW_��.�zߞʶ2�8�
�=b���Ud��$�O���w�B[���#�HS	*���Ӂ�s�z���Y5��ri�U�T��Tj��i���
�2����<�n.#��D=�0�f�@��k�j���jV^���M��΢�φZ���57HW�qyZ1H4;g��Q�) <�Ɂ��0|wRc���n'M�sR �:c�?�����8/��D����\@݂z'�������,��{{y�H������5$�|ct1GՁ�e��#Q�~mpo����8�3���c1�/��9S��ϋ�}2�v[8ރ_͢��ۢ�����l���B��������+\��=ml����c�R����+�D����PRR2W�����{�TAN�QqI���K|�'�P"�]�^�&Z�6���N�,�ER�o�7E��n��x�>+:bQTR��A�ws__�a��q��?�HV�A�\�l�dR-�A���
��:��oR�w�4,߆�m�:�O�\�`��A�ĝy�_9�jqb� ﱜM	))e�S�WrL�L���v��sG����Z�f�<�o*@=x<X@�sv+ǭk���*��9�)�r,\�;wLf�Ht>+��N���lKd�~wm��t}�T�Y�m�vT��z���92�!si?� C��M���G�ow�dGtY����bF���s/*`h��k�O6�?yjXn����JjZ����T������O���/q v�(!c�0sн6`�4�Shʧ�k+K�Ӑ��&7����_��>8�[�5�I%�s_QV� �N^<@�����3|z`X���F�-s����d=���Wϲ�ٲ���z�����?9�P��G�;q����n՟N�5`�A��VYE&��LJG�V����Uy���C���%�4 ����\����^��ɵ�onk��Fu�i�}�-���Ffx0����x���<�V���&]����ĺ����x;*V^h�i�P#�$M�^D��(Mo�3�Z@f��Â+
-��,���3N]	�����3��"F) �%=���<�\�6����C䃝�ө�h�C����A���R��a�TA�px*Ԍ[{����P�4:`�}o$G��>`����?Y�y~�6-��.&�a��Uwt�/�vJ�gN��65%�uC)_�#kL����0������~6=-FR2E\5$rº4|
�����TL>ywڢ�2�SS>��mo��4ޖ��:<7����=R���,�-52(��?Li��)]{��!�5D~��v?�����;q�`q�o�j%�{P���$f�Rd�g��sNi���y����`�²s��y+CeH/>�u���~?�X*�57|�}k=��k�2�xO��2:��'�A�-&����Z/���"��ʺ�,"���g+@8K��V���Q��)�ˁX�٤�bP��_�J���↬rV �R�٫��j�p���L���}9e]�0v��������SN�� �v8;B���lVO�Z������:��a޳x�P�D8g5Y�4�3�r@v�Q�L��|e�'otm��V��2˶��������0m	�M�Ce�2�v����V��M�)_v	:$::���:Id:��b�L�Q�����5� �c��_�X�09�~ �� C��7�vv`�|8p���XG�KF �zm;��c���#.T��	���QW X0�{r;g�]�XtB������\��5M��
4!�y|{�O���"b�-�p�Y	P�4�8#������q>6���z}��ʖYz����z�j ]���d���s!�^�ţ�#�;=�{�C�����x;{n��=	�O��*M��E�i�y���k!D"�*s?����)�w8O�V�"�N7	}����1|Y�2�����1����G-&�˞L;���MhMɳ'�2�t�k��s���Ծ���XeǴ��N����!;�jm���UM�9��d�.Su	�y���H]�2ZI�Ъ�\�sq�EN���o�ַAR:ewD�2`\G��3�O��&��Ɉ�ϖ��w�ev��U�+��7�JT#l�TԴ�X�G�i�UUҲ��p1�-I��2�g��LTeV���A��`#t���v�5 5�"�p�v������טp4�����������}���\�a���n�)���c�=����)�>k����J��$�5â�@cY���w��.�I����LOȯ"ڥ����c�%Q���J�6vр�;�{\b�t�0��+B�R����_���D!z�ݦV�� Y�nG�
�{���������v�W�=���n%��s�~|h�ir��"!|�|���g��VDYk<�2�p������8�v't����fW��]qd!*����ېN�P�x1V-֩��ɃI�#ڴ�0m��̾���,ćv�qlm~>�L<٦X��]�\�6;<��W����!�o�ya�������F��Ga{��.�L�I� Ag��~�&����Ҧb���M˾���JE���@km���I����r�S��ǋ�c����avfo�\�: �DB�a|��^�=��_��Υ�e�w����42kOA���4ա4����e6����v�8��--�M4ߞ�TvBR\�����Ó�r�h-������䑥��7?�8�����D*�`�r�����k$� y`�8d4�A)\F��%�#���<x?=��1�n&b~j/� ��?j����x_ă�y6���:��X�wQ��$���Z���ۏūB��9vlc�.�s��}-*�L��h#��(r��]P���X�6����A6jӮ* �Rʆ3I���ʞ��Ko0]�o��j���n�|�g�P���>�߻}7���ck-�n�EʧᎰ�W�C�wk�i�i ��n���I��2�Y
�_�qY�hI��"�EO���>�cf��LPo���EN����5��L?���%#s֚�ț-�;,&(��%;���;��ms�������3fy��GK��8�E�y�.B݆��o|R��r�A8)��P�tP�ɔ/Y~�Hg*_�4�����iF!���A/᢭�{�@b�zHr ��p]v �_ꅎ
TWq_)b{(+��+ooXɗ��U.�����]C#�OeM�W��.�� 0.�`� ��Ѧ�N�_����
8��L����ri9am�� qQNx���� �[c�O����g�+���+h����ъF��9�I��j�����?2����~)�m!����pg�ܒw����I��	lC
�X+�Hf6����W�% @t��z<˩I�޲�.����=��eA�u�/���������5p8�!	a�,R��p��I�(J[έ;���6!,*��>��Lem+=?�$
q%���·�b��t8��0|P�ܡ�`kd�������gXͿ3Xɝ�B)8�����H�2}3�s�wO�t�A��U�m�wF��wp��U��̤��pDՖK�E��9`�zi�������ll;w�6�r��4�S��^�-z�DV�m%8q�W�$L�(�+�zЈ����ך�����d�l7��Ёh2�W�j@�IP���/
E�H�g��`��f,�ʃ��W�_~��pfJ:XRQ@���	<��c�&� ,E��/���bUY����Ψ�+�u9�TGO2U�]��!d�jCs�F�	��ti��Cg���̻.�S/�v����i
���)x�.oW�*���D��c����"�*�Pb��.��{�%(��l��51�G��e��e�eU!8P��ܔ%s�|�s�2H���ھ-�BA�Q0~����Y�T�'�XЂ��WRK�*Hʥ���i��j�m�M4S�;z^��2*W��7@^�����(O��-7�׫�X� 
�ej�>�_�;휲�����ݷ?8�*�2г?6�N���yv�T
qc��j(7ⲃ������KP�c��_v��>�}��&�JP��e�;�~℉�>xǺ�K�dy���c4�(�Դ5��o���CpdA\��I��ܼ{��ۡ�4�2�:����8E}���  鯃����2�ڷ�~'�]o�%�tGt��MZp��r���Ʌ-^[ШH3�=}�Ӽ� �?��,d?t;����K�(x���d14��Zn��Q�
J�]�0pc
����ٖZ��V��Кl�d���J�5<2�4�^�U	.�iIře �}�p�o~L�����ܲ�2��mԉqs/?������u��Ҭ�i�9.�F�NM��ܧ<ӌ�9/!�ld�UA�J�>�U�^a�Y]Y��x�XV%.��_\
>�玟i�K����1�m�a��<,��žF���Kw�Ueqi�t����P��[�\�
,�Q�-��p��n��Y%Ϳ]%�c�\> ����9��t.a���w�=�gz��pB�+yh����YX�[��Y�ޤQ�.�!N����x�L�=RR��V�P�D4���d��xq��ipɒ��Ӎ����r���H����	���i-��ex�gD6�
�6vS��X9���2�x2@�=\j����'RKm�0n�j����yӘ[F8O,�f�B��v�th���M̰���#9���I����ot�&;�/��%AaJ�2��O���H��6�xY6%��K}n�a�W�{W��b�crEl��ݚc��h>�O{���|}  �;��ʁB�ί�g(ګ��FC}{��-��6q,��?i�ȀB�����Y�/0�Nko&�f�4jGyUh��������󢛺N�R�lE��&���:j����3����K�hxz�	ZI��D�
��R^�X�D�L�$Y����u����x��-�/DJL���[ ��/��s���t@�ѝ�x�T]V���1F���W��9�����F��Se��c����:5�+bRC>����3$ ����vō��]�{�Z�)d�l��w3qO��7��͢^Y6)�йlO���d�I`UN�)�u�ξ2�b̩�E3��R�q�� V��4,�y�o�jɪ�5�Dԕ���d>%�Cp��-I��(F�/&F��Ylc��q<�����@����) �{
��?f��؄Cb�rӄ.�5:Q�8��_H�{|��ꉜwh��o��X�����m7֯����r�(�L��Y��g���%� ;�Q�v�و2:����8�S���U	��̎��*R�4nײD$p�3&h4�6�.��?����}ZǙ��u���˘���]_����L��E��qCy<�\����]�[xN��ҿ�ٜ��Y�P���o�Cpk�V�SUp��Ѵ�,b��v[8�A�/�It��V�q)����)����#7���E#�%�ĥK�k�-Q:�\��id�`7����&|�Z6�.W��o��X��%�ڬ~@I���K�B<��q�y��������{��B���"G�YD�3�_b�����w��I�|��$����-0�#���&�3���Xn T��n_�9u>���&D���+UO�K�iq9Z��<(����XE�Vz�i����l����Y�)��>ۏ����0�ų�Еue�.�"�2�Kl�ɳ����S�"֞+�������ﾋ�/̡'VL��	V�uNމ��BN�)�N��-"��+=!Kߴ�ܡ>��M,�p����{P�S.i(���.d��|2�isy?g<I%�2����00��(�;n�VvƉ[��7*C�d���\�����T�DL��jlLI�$n���`!�hXCZ�À���Ńy~2�P6!�(�D['���yb-~������X�j"���$;�W�˲d�[�A��gD�A�X����s#Ƌ�]�*s[L�T��s��44�cy1�gH��)P)�?�ĵ7p�"R����Ɉ�1#������X�O�����A��K������0R�|JNرoK!�y��tr��
�=��)�N���j��^����d��F7�������Z4?������I�S�צ�L�ߒOG3.��:�fT�3��1����KK�$$TήR����1Hw7(v�F�˼��۶�Fj�c��M��y���L
�l�R�l�u9C�m��S iN�UB�X����g��!�hz�A�|"աh��"�����\�Ϭ�|��@U,�=R�'"ǥd�,/�le�ΪA�H�ۊ�/�lg���,6>�sX��U�H������	����37�;�������%Jƶ�eq$�����u|�J��G�Y��./D���&ު3;��� ���Trsbl\��Z��uS��_�yw��!&�۠EGAz��0A[���W8��Uy�Q�g���#<��sH���w����Z�`w7�0�i.�����S�K�a^v�>�j]�9�@ ��nx�W���\�_FiP�퉺��فjLq��z�#ߐb���P-F�]�8���9�߲�E$B�	;�a))@|'����1�:����?��~lE	�+��v��[�	РDy�K�n�,jՈ9���P���$�I�ƙT���}��m��m}Yal��Rr��L��� [K��K^BN	Y�<i���2��{V��`��2	�Äg/���:;��C#A�\�VH����	o�O�d~�(S���P|����fX/V�qˏ�,�JeA����+�7.��A�|�{9���
7���ڇ[3�Ph��J�B|'*l6�A%"��7!T�	�9'x��Ɲ� ��������9����´�w�4ʨ�H���_�n�)*�� ��A�/� v�����\ ��#M;�v�w��G�׸-AI�;I��Z���`�����B���n
l����Jk픦�<�����C�j2S/>`׆�jqf��ro�BLgן�M.���͘�9չ-�|;�����a��oe���#�l�ץ����YU��R�\ö�g�4�R�ј�Xg`���6	/ט0:1_D̧Ż���L��8���iL�\� �����ak)~��)�q��ż�i�,����=9��"u����0�X��-�O���^���vPS��u�n-��Ǫ����+/��Z�����$vw�b���e�j"��|-�5_F����׎�X������Xr��A	$q��WdH�$��`, �r��ϝ<Ū0o̩0�wK��
��(��*zW�_���L�5��h��!�C�o�OG2��1�d�5:��dv���c:�WA���T�m�k���(��#�v{ne|�9�'�q,Sl"���yT� iC�s�:��mN&Mj"tk1|Dw���W���1�ѩ!o�~�v�&s_T?�����1ҝi�G~���ph�
�Mp��Ӗ�zY)T m$��#�?�6�h?���g��Oee=�IR)=�6��^1���o,��ת�%�Q����f��f���f�[p��679{��c�7oŅ�mU��<�2N=�q��ݙ�3����+J@vю�z��	����~�lY�������\(���ݏFA�2c�'���m���`�#`�!/}�$w��R��V���o�d�b��͢�l@�<<f&�3[H\�U��iej=�ٝ�6�L�l3;��or��E)ǽ��0D�4|f��+C%�^.!��ϥ���Τ0�@9k�U��n��nls<�&�yz�
1V �(/)_���z8�*u;�9J�+1Y��P	a�������&i�ږ�I��5�a�&���JH"�U��38g�|�~
2uK����Wx����j�������#���B)����;r�h�DTt��r
I��e�U�yu�a
����/����.&܅Nq�}�Ed��=`mʍcRokr�-�9�E3��G� ��>�/A/�`#�R���3���2.qi��f`{��^_�iD,�2��
	=�Ĕz��d�=,�������r�uY���\�$3���%1�?����<�	��������KZ��
O��ړ�4���p������<�gn�:F�_���7��Q.)Q�est�T9�9��yH�&�ߏ�jg��8��	<y�Hɺ�G��8�5j�@h����o�up���!�)�>�F♭©��f�a�Bw)Mp�9�.�h��↸q����n�H��甊׉����# � �?����OP����@v.ъ�=�Ilf�	�p��P@6k��F�긥�f���親E�q�s����IX���R8N���K@�eL?~�!��o��䃶g7K�	�lk+1�*��ôࡘ�����3W�/hǉ(��	5A�c�MB��ug�������j������B6�U��:x�m���ӭzމ���u��/L��˴�S#Z��ϼjh�GpC
�c�<�s�i3~eU�Vb����$�{
L��YJ���ث�r(��V�8�ֈ��R�2�zp�\0��E��gK��8�����~��ݼ3U���5�`�bmQR�����\I�έ6���6�����Ӭ�WF1�M�
�o�did�C��Hfy��wY�R�?8|3���UA�g�5*�F����']�p�,�k��f���q�s:��9A�?si8Z��0�AS�.yj��79�!#z	8L��y�T1���J#�D�l��џ�^����0�nH��d�䈒���.ǺrI,�98^�ڐ�1�8\�P>���[Ӑft��y�/�&�s��N�E=TP���f1p{�K�I�5DVM�`(7�(�7��*���Y"���� lx�Ķ @<�s�e���f.��"Ut��Dɿ~��j��O��.�Ps�S���q&�/\�JҾ>�_f�2U'�d���(=��o�k��ĩ�iC�so{�9Q��&k<('��ux/!�G4�(�H+}��Q���V����4�K�Ec���!�9)�ţ�GJN���Q�M���(��״��1!8@rk���:�AÖ�%�,�뷟DJrŴ�b�U�{K�Pj>LDJ�����2�K�Z� �(��|: 0g���H�&(�V���./w��E�$܂���v���w|O
~����H��,�����[��2b8&5�8��x�kr�l�B�̷f�s��%�#�z$Q��
����	�'=�X���}4P�,��TA��vW)F.�S��v|�'��З��`��Η7�~���m�W�d��q *�H��~��,�p������v�?�zz5� l�{���3�h��.��e�d¶]iW��L���BEJ�&�\D��2�(�w6�G��^�/%�Ū��U���&KDM�g�XZgu�@�L2����f�e�9g�\��d�n"�ު�����¸Cࡃ���jL���z���;4ac�^�����-��<�36+�_;����)��'̍�(w���lg�F��5L��bΌ�~�����9N�on};M�����}&Q���9u35��fX�q��@GC.=7��D�s 4$�E�7"�I����(� �v�T���H�`Ȉ'��������5�� ҕu�{!���F68����]�]q��p�g���[��b\��F:�����,�Fh��{C+�b�	��X��!���уT��ɠ��ϊ/UےΠqD[���(gZ���V��e���R���m=����¾4fֻ����P�2ip�i/f�M=���lqC�ö3Z�3LT�~ ؕ���i��;pΗH�f�q�dpq/��H�I߁J�f2L8���^����{m�U��������n�ID[�p���,δ��&_i�#��x̕�r]�.�8��3��E&����l��C>�<�+��/_?�?��*W��|�q��\{S�+�dO��y���Z}�����o�!e5�\��hb;�4?%ۉ$�l]3t1!�
m���i�Ŋ�D�upp����+j���(�5]ﱥ፻ f���0�� #��mE3�sT�'ȻX'�x��3���^���,J?�
��%���4R/��(�<����D*�V�"�ݟ�s���b�q�������h��d��5G��(�A�Z�p)˷��2�>�%�[��?wX`o��x��k
�E��j���jȨ�������@Oμѿ��j�`Y�N�������h��Rқ����h$j��<,b�h�k�Ցx�"%�]A�}8����	ڡr�c[&2�ZB���b����&�t����|�O���f�R"8}͢0ʉg����<�����@`�op�� ����a�4������� �٨�l�3c�)��6���� �������폟!BܥF��[�r�|�$Ē�B��x���v1�g�@�d�9>Y����W`NC�t��y�
�x�o����x%�Q1@)�m�d��1�0�j΅g���؃�1.Ν����с� ڍd��v5�C��\9�����R4�n^S͍��z��V[�Q���PD�;~	����b�v�����y#�*=�]QI3����2��SKښ7����U~�7"�wi�K��@-�|�mn,�Q9�OW��~�5�������O���?r�n��U��U�x��¹#�\��V���#���byJLNJ��mЦ���ۚ�~���7�w9�.p+�7]���"�?�G�3Wg#�.IE7�3�W��U�o����z6�bAdл�D��v-�ϔ��ٍ�ٲ䝻m*O]�Me�"g[B����,@ MƏ�X�v��>����&{c��#i��6�a�ѩ���ݗ�v�_�.���d����K����q��zF��٢Z%:���Xg��Z�+ G�
�gWP9��͏�G= �?L�Թ�UR@�gMR�AeX����	[��������M֌T�g���|M���B˓���i�ԇ��֜����%j-�S����n���@��я����3�޿x8=��i޿l�쭷X�*=l"3&�8u6��M?�kj�u��Ҁ����1a�U��p#�@�<.�H��j?��١m��ơ+4�	v� C���T	�D��`B{�MF_�Y���ic���`��c�t(-�n��x��&�Ǖv�Z҇�,��&� ��P�E_��/2���v��S�o��>���@�M�� ��s]�Lh�]�o(ߡ��1�c�ִ"A��T��Yı�/����>X�r��NU�ʵ�p��9 �v���=j��7&��{��͓���@�5�"'�&D�\��P�7�-aV�ۣf���&�$�l������@�R�{_��C����lyy�mn�(=ըפhn
�X��������o�T�2�	14�/�*���|)�$�U�?䨚C���g�RH�)z�1�=���6j�Xzt�r��.W{BE��UH�[�g%�Eݒ6�,���l��,���
.�H~�ի��s�m��5t�"�֛��qT�D�#�-D��$�,�@�0�_��I2J�	�*��PҵC���l�D�'�hW�����7}W�f�1邗���WV�sf"f��C�3y��0N�P����~[& ��{h�E/YnC�:�rZyi��T@gC�'�[;RK�D?r�Y���b˸5{pCT���ѕ��#���YJ�~���H��	�����H��c�&d�5
-�Q�����q�ڹS���J����y5�	��(Ͻ4�O �`,���lݫ�Ҵu��2���[}X8�	�RF�n�2��ak>��al��Ѣ}���w㏪ �7��)��Cn���y��J-]r��EN�=8I0�.eht��Ί�"�j��(R� �U��z3��'6CQ[ZG����c]B�M�4P�=��ȥ)aa5�s���f��ō���E}� '!��@�$@��e���__�󘏤�TdX((���e�<8ʃ����:�G�Հa�r���w��.��u6]��q��ZԢ�����j3n�*�J]k��Ώ���Y�`�;,�f��T��x���fc��Vr���3w9���H�A�WB�˝��x�K`y�_1�h�2JJ,x{�Q��_���\�Z��L���	��!��6���b����
�W�I�i߆�:2
���ç�h��E�U��ś��ؒ}Y����TU?�D��uN-5:���c��2�q_3��F����GB�4�u�>��n(!��r]gy y��_��u蚷�I����I4�0�y�`�k F|�QѬ�����("EW%���_� ����P^�w1R��/w�|�E�m7��h2�]N	�$ρn��کn�����h˶������R��ZFS�E�y�L5M�g��E��%�|�.�) �q4��r恴��$�D����+�}Ι��=���,������czgjSFq�K��T�Z0J^���T`~�*��:X���(�[E`ҴcD6���8��T��<�fv�]�{��;�B��L�̓^:_7�6Ua��$!�%;���Ai����N�A~�Pa
��$~�e91��`��^$9�pp�ʅ���@c ��[Ŧ�1wOJ n�~ߊ�ѶП�%��8�L�1��.�'ɔL�ᒬ�J����+R3���� b7�������*mJ���}V+́?�A�B�bo��1��$*Y��,����2��'CD����b(!?��n/����-S#�F�}�>Հ%�W ��"��)7���_"q:2i��dx�§�(��$*�Ԁ�oμ\L�Cj����Ja����X:�	u�̐:)�ܾ��'o����}���ƅ���\뵷GD�?M�)��y@���Bne� �R4i�[ܯG`¿�D1� [w�O 晸7׊z�[�
|�1�ݦ�-q��|�&eh�Y�%��̻-C�'�����|XGw�.F
ֈ�1�x����f/���r����=��)h�1�)"㍺e]lT���#>��������Oz/��+C���֣��/���7΀�����՛���S���#�şxo��`d�<յ���_��:MvQ�)-\����a8�Eߺ>�V���[���j�ym������%O7���.%O��W��쳭U�dQI��L�����c��Q�P�r�x�Sd��������l㒗�7�Q�~hA����F}��#�v�l��~Rz�/WP�M��3z��XFs�qN�=��!,U�㺟87y 0��?\tx�P��?��G��eVn;���i�/�����4bE$�A^�Z;�!]΂h0�z����y�Y�5Ԉb�5�����A�|_��\sJ<��f4OoD����kt����2$7o ɗ����{�@��k��x�iߒ5���[�^z�h�]�xZI���u�+�m�\�ٵ��}�V<܈.s�6�v���m'�B�����Is���ӫ�<��R�!�uΎ����`�P�\����~h����3�ɶզ��h���]�c�N� ���E����>�q��W #=��bHI‚b�g�y7�g	6�G��4'�~g�"�^�Rq�Rf���<��:�&E�?8a/�����j��޷��d���)UA^G_El	���2��w�\c{a^�&1��Ra6��W�%bKK���Z��bJ��|��Ɋ�������V͘|1+;Q=�H��e<C���JKpk�J��0������5P	��0��3��' @B8�$����`�#�	�S��-w0��i���(*���i��� L���Z.Uvߵ!��M�:��3�~`�+�[P�Z��L(�)�԰��ɷX1>;~_M�v�P�㼠��}�"z��^c��k^�RV�����@�hC�Y�!�
Y��A��m�gk��MW�S�XZS�B�[�a6JY�K�48�PШ��K�\�9�[�]�]����и��^#���OA�%o~�c���b~��S�|��	����I~�*�!]�T��r�.�]���\������@�fI����
7x2q���6�(A�E�8M�Kk����v�R/��o=�A���	��W1Ĥ{o�۾("2����%�&���&�Rjs�ZY�r�'�o��$[���p��A�<dЮ�t����I�����&$�!�Q�&ev�����co��h@P
��f�I!篢9>(��{b�Km"	��M{�����'�=��oVJ�X��YX*�ě���~�/E/��M�+~g��.��捃_���O��q�U�+���s�8��sP[@�\���+ΛD��e�(p=�LL�t���p����ge���
r�/��z^�u=��r\Lvg�葽�L��YC�.Q�D ��B/����kN����VX�b����'��Lܢz<Gp�d��D?��|*�V��Z�]��W�g�0�~8���$��ߋ�>0Zp��VӦ����D��ؙs0�����#���X�*�
�W	|��21�a�D���E`n��E��������P^�Q,�Aꨂ�/��L�HH����#.��Y:/�����+�=�%2��0C��zX��"�����cS�ȇ���=��ث����v��ɣ���s��Ɋ_ r�I�\���ET`&��B�Bi����	���y��̖6�YFZ�s�Kq�����nt_:H�~L���:�X�,ė�z����� 9MY.�k�/G?!}�e5��͖�Àl�w�'4���$ᅭ�958a;��&7繕��u�L�l$��<�6
j  ��K*7��K�K���5/d�"��|fT����O�!�,�n�㨩���6J[��+�gk��ޅ'�A/hҧ��N�DIireTJ�X�#1��弋=4�B�-��QX�d�O��	:U(CSۆ�`�Z@�� ­,��50Dp��8�UP�и�.Q��ӄ���k!���(��!曽�����Dr���Ӹdl,��� o5)	+�@Xr6ܔБz�4��oqA�$�ĳ�XY��[lq�{0���H9��냬�ch���5F��+����b����aa�՞����e-�p|���=����u-٭v�bTX�k\�li���l-G�A���~����~:�J��t�_�h�6��i���9��Ʉ����;���59��`.F��$?ᶯj�7�2i�(ۯ4.��� �@�v���LX���ϸK��+�N��gY���F6�6�)`Z��ׂ�W��
Mm���a����m�P��2�[�WL5g&�	c�r���l��wV�il/��թ���t-Oǿ)��g`ݲ�qs�x2�s�#8=�W��k���lm7˧���F�j��GDS[s�y�"o:��.��X����� �ll)ª���WtW@J�~���JE����>�}9F�$J��)'�(�G��&���.�����8���{~(�VF�ᅼ)gX������bA��^�g���v޷��P2n�� D�*/Y4,N���C��Bi�i��E���p-�%N��#v�@��0������ˎ����
�{�%N�Ϸ}����e��F�\����>7�L��+�<��w�ٴ�=��$��;}�AѪ,%�:�I4�8*D��D4V�f�%y�6�\�v�:�"�g�%��7��>�z�A�o�7�Qvd6=A6r�|�`�6���텓�2g�69�o��D��i�P��`)�X� D�#��^�W���R�)g�c�xsE�S��������[F�MpZ�9��S�������4�aNҠ�uX��?'��������09�1�#rw4��j�'������\�v��� ��c
����T��i�\��R~�U�L ("���<3�_���a`�M�v�9�9�������{��Q	M�5�`��Z����C@�y8b��z+�H|�ү���`TBg1�O(�ȏ_d.��ӐL��=�y�vlʻV����簈�`ޫL����>�L���F��a�4��1�+ez"K�A�R۷J/�a�U���/�1W�
�/����-�g�����j�-&
}0��s2���&�REl��5���NZ�;a98�$��^�t��k	��<��h���Ϣ�nD9y Cy㵤��i�Z_n���C�k����J_!lJ{�� S�ؖ�������9�?��{��8�]:�ت�m��\���!�Z�{0Rq���`�� 7�u�_É��f��d�v-MkD�4��Lv�&���RB'SW&[Lq3qڕW�킒�1��/���7o�8�b�|T��`�sG����*;���U��U���k��V[^����b�d�OZ�����ՀU�0ɞt�_�Q���O�P�w�H |�� �3�3$��P<�|���~��h�emG����]hD#�8x�!�	�NS��1k���<?�$7��*�7!X�@�˚���C�v�\��8��YNUʃo$�ƈ!����s��9`b�z�Z#��~�*��^#w���� �!�2����	�?���]������_�r�`��O�	��R���!��8��WtL��lFY��F����/��оd�E���%eyJ�0�!�v�����E{.ԔuA75�����ok������>�xOT"heZȵ�)c�e��F����F׌���A�$u�X����6��X�Uρ9�:v�o�%!9���D8�������f�/	"ap5��$���i�9èٹ2j�73"#�v��3Ԍ2�$c�yK�ϊ&�̅�o�֊?��Mַ{�&���qC�7�A<��o��.������u+�8*x�=�+�����?�B�#S�2���y�~�=��:�φ��\��6ކ�"��u��I�Jf�j��P���>�du!J�}��h	1=�K9��h}:)�ܲ��dU���sNk�ҟe����L�T�����[��A�k�0=�# gkMd�J/qЙ[��_W�Ү���X����R�7ОԼb=�ǈ w�z�_֫?��4U�C��йu���#NRT�Bu	��A�F��b�2|X��޸�ě2��F��iu/0�7v˜�`2�#g��x���x\	��}Ւ�zY�������e��ǈ��~���U��p����6g��Hn3w�g�NAh�ՠ��C�Ƕ��O��ھ�Kf�/���+�������4 xlң}9�=W6��aB"�g��Y���W�(����:8v
k�jw$���+�̕�vh�Q3i�w>v]k�yZ����`w?~��
N��c����2�s��)^ �	?κu�s��q�!���^��,�؃��n��Cp3�8�j��jX��@R��RY�L�]�5���?�gv@K+\b�y�X �d1	�bC�G6���q2S�ǂ�� mm#�n��k���G��B�L��	��(�Ɨ���+x��4X,�d�9-(�9ԣ�:cW7�p�zջ*�J��o�l-�Ͷ�C1| ���;n���8�����6|��@X��d:�q��WH�JD���*f������BL���
�	��' b��!�Z�W �(@д��^V#�����*�Q��{T)��g�p���'��r��_RyQ_���|���f=4X�?!�[����.�dַ��N|>�J��aG�B��N��=�I ={g\���+9;
������_�(��=s=�u5T�=/x�V=󶢟9�=ԕ�rGe�c�u0�yʲ�] �}��ɑ��K�q�jq�P-YV�fL������w�hm�f�O2704:H�8PZ�<�HY/�`�b�&G�.f>��-[?:���X@}���bw(9$>�*�5h?$��8��<vi�o�K�]� %��4�uؘ.�2���F�����2 �m�z����� h�T%w�!�Y�4�x�᫓f�Q)<צb�>�pc����oRZ*����{O�"LĲ����c6��L���z����'�D����QAJBJ��3����h$�auK)�p�$J��֞i{��j��@۫����ʷғGͺ��F���8��͐l��Tru'V��@�cT�ug�*ۢ���7��$Iib´ʘ����(SM�QO�A�	 bv*�vߦD���z��uu;DbQpg��q�"�^��э�'��1O��=UT'��o��&%H�G�}B���98+��v|��»�u���hˤ��4�V�c-�p;���x\�U������A�G�*���-i�'{m�eR��k���!p�7|ழ7�ʾ,Ki�^Ge4��'���܋?� �'{�Xk�#D���W��[#��'>�k��I8�Eni�����M4��o;���7Sʹ=����܆]sgȋ&CI'�
R�r~�U2�=V~~.D�#*ކ����o*��r*A>7��7]x�<Ģ?N*�S��C �����}2ȩ���nz���ڭf^���Sݩ�:�V#��b�kRCv�
��U��F�����-�����f*����q�2�j����лS�4�A3z��Hq�̀��n�.~"��Cf=(
�EZ��V�r%J�OF�����۱T�K���d����\��ƺQ4)�1���Ʀx`|Cu�P��£�
.Ny2�i���=/�g��X����6���9 ]�u�@g������)��_<�0T�3.��fy��iǼuR�&w7�~$+�r�R����x�S�O�V�
d��x���]��c����;�������$�v2�@�"�-���;�bx�%1���u�����<�0����B9]3�2tr�3{�ά��UK_���Z�,�����h�Ú A������@��o�{�X�i�$��@���u+B1ې ���\m����*��A�i(�r.B��LZ�~���z����!��T�6���-���+7dwɜ�ӧI!���zM�Kw{4_#֮_��h�?������Ѵ1m� '��Z��}�� �%��i2��g���\�&�q��t\�Z�]Ǣ$�G���  �����G�5�*����ىz?Ij�/�e=ǧ89����j��ʣJ��P��נ@R����в���t��-H��ε�6��gP�,���KO��FM��[<q�1+uT�"����4<�w��d�j�uĦh����XY�fh-iOO������-���1�e���a���T�(7Qc��b%{&��&�ñ�8�ӏ>��[�r�a@<��T߯z�x��8����	g.���r�}�|D����w�����g�WzBע��Ku�'%�q��@A���UׇD�	�LY�i�Q�H"��e�\yy�:џ
N3�#m����(� *��f i�����G�nB��2������RA�	e$~c��s�F��Θ<��Xr}��]
H�r��ca-E͗J�P�ղE�{`���\��
���8T��$y9@&���A�ҷxo��Uc�?C~��1��U� �t�����~N\��r`>{�]�F�J������5��֍�7	�:�� "���V�W�ml����b�=�*��(�X-�QP$)��v�oz�V����C�\(W���6�s;�_E#�
F��{tD�PH����tW$'�S��_dU [���y�E1}Xc���K؈�F�D}�O����
���LݷL��e�c�{++m/(��na�n��w^�꾗{� ��Δ�Hj\�,X��n�C���R�}*�n7F�|�l��z���"Q�x�v���`_F����6��Pl�v �fς��(")?�����(Ȅ��}#:~�M��݁�Ū!_��)�6�5���C�1��N�ekD�\*���k�ԚZ(_���U�2'W�{���R����m�����z��ֳ4�ԁ���<�Rp��a]�A�Q�u�^��M���٢�� rڔ�,k� Æ,��A왴�M,�T��u�|��!<.��
MM=�T��2�aC�||=�b��	
��D��4���]�sZ�|�uh��7�!�Q���ڑ�7n��?f;>�r�v��wj�$��}�J��a�-i�cQ��ht������,���b�Y�{#�U��A��rteV��Q� ?�C�ݡh&M�����=i{�m��w��K={G�A@(.�a���0	�����:E+~�`�Ѷ;�{�
=,��O)��q�u��{&٪B�Nj�}��K��v�`6 ���Lr�<�!�p�w�tt��Csf<	��+{G��?EN��!p|P����Ysָ_���s�V�e��Q�IF�>pk ZycZ�M3u���#WEλ.��.�j��v�q�m7�=�1�� �,�ՔO#�rm���FG��v�=��l:�$e<}�!{o�\Q�[�!�y�I�LݛL�?|����u�����ж��U%_%�5炘�u�Oi�!o�8ۯ(bO3T��uMƤ0V�����@E���Dw�߾}�hgg%ؙ��/�Wشǜi�D�s1���F�k�!j�l�.�<LS_�U�s��t	-�}����N�����-H�lt�Ǣ��������
���f��]�T��8M�1������Sjq���!9 ��L#tg��r���e	�Z�_*	c�;�ĳ�}�������z���w�"�c=��q\1�֝*�4��F�g�N���yeAUPª�"g��O����{=��=���3�;8�B;BA�)�=�xL�B:RA³�3���/��V��v7���;ߋ�L�"s5!Goy�\�Z�++�y�>�"��,I	k�a0���WK�^:��c8z!Ǵuo7s�B�l<�u��5s��g�M�КS=�O�oq)��r���.2?���A�f:x��V'K��p���F��E���s����f.�z�\�+�I���ر�Ke#�r{'��UN(�m#\�Ӛ85ĝ�C�:>��
W�7����$�u'���&�� ��1��(LB����
��rO��t,��5�6�������
���Ȼ��u>w��0�b>=�R�8i���b�cA��/��/�򭺂��w���_�V�KM.-'w��+H;��.�t�r |3���S(t<a�]夑-)���a���//[�#���.�K����Ү��P��쐎��k�'dXZ�$y����QN|8��4�#5�o�(�o��_�Bt�T�k�P�0��]*:�0����$?E6�9{;<��rQ&֚ր@�&�I���<�Z8�ԡhI�Ȏ	�x��r�E5�O���sQ�'����S^1���H��"C����ͮW,u�9�EWj�<���5��c��b���̌_~�&�i��M��g#�"TSM����$x�<���R8t��".��G_$�A�&�H���n:�O�7O z�k���)��N���P^���[�C h�����}y�u�-+�Yk=)�"�����?���`?mw^�E�+ʫ6��7���5:�/��5G���a������<�U�"Y���6	��qgT�|&�w���~�]�"�;��Ek�9��'X��>~	����+-�ߧ�����>;bȼ=v c�Q#[U�OD���e��ô�k,�J5����-v(^�р�F!iR�T:������S5R���t�X7�1�%=�uUL,c�Z��Gf�3���a�c<�=������1#1��,oK�z��!EO>�ߵŒ)Jzo�O����)��L�r��ҡz�n�'�I�(y��~�HA]b����C��(<�y���;	�g��u��M�Z�Ń�O�&�� ��Q��HS�!�H�KT&3:u~�?��y�m���»5m8qS�8�1��d ��Ox�@�RS���U��f��I�ջ���D�h
F��~�17��n}�9�GO��/a3�*�i�@P��:���2�7�AC&[%>\���A!��:N��Q�h�z�� QDWs8�Iî{I�ן���Q�8�x������IZ/u'�����$ɓ����J�����00��R�C�T>���)v��zٶq�Ed'��� ��((��&���j�+I �?*���ӒA�^������'��!4Z�w�������*��lE�?b3��Y��������P1 ���2������\��1��h�(��ٕ��f�����v�v���B:�:� +ё��.��|��������X^}��V�i�1���;3\�:N�L3�N�cd�)0�1�������7�0�8�a��B=�&�%VLA1�}�REA���@o���n����� Z���HF�#bXe>�p����z5ȉ�[�
�	����B�&��@��'��|��7�n�Z\�K��� o�`뤳�%t�'�%�<�oƦ{���\Y�l��=z8S�z�C��Ģ�j0Zl���l7s}�mz7̈���R�%Fk(ˏ�V�Z�[�O�#�l�ܲ�u:{�i=� (" {z�ޗR��zg}F[&��:M'��دp�m�N�4_"
	�3Y��	���0��u���wn9E~ٳW5ZN���U�k�',��e~8^��Jg��h����YMd�m/�tu��";d���`�Z8Y�t�q�,`�	U%s:���S��+��n8{���ß2/s6�0�,������E�N+wU�9诟�-!�D��1P��Ɵ����C{�[����x7Z�W$
�&�>(Q�e�6c������^�\��T����J�#5�U@��
ē��8*���L�Ӱ#�"b��X��jM
:HxC���M�s�'4Ǡ&|���z�&3w�˳|�[W2�^���vi���\�8oS�g� 3�U=��h�"Db��1}]� �8_}��`?��/[l�.�	9�!���׿�[`��U�/xKeա/=M2Ad̵(;�ռ�'1�t�ſjJ�7��3�����Q�����} a��s���_h�oZR%�|�Ȫ6ܟmH����r�����9g����y�P�e�Yk";��X�뤵�U8�?�z�H.��|�<�� 2�4t�q^��J\��a�Ye�o䧚I��M1? �c˩i��/|M�h(2��֊��rX_(.��1Wi "S̳g���8z?���oo�c�.��O�X����HM^�e�j���S%��!�hȚ3����ێ*EP"�p�Y�׊�~VA�<&��A�k�:f��I9uTN칚cV�[��-�}c	�N��Ώ:�^�f�3�"t�����y �]���R��9t���h��"�]``g�bt�ߘ:k���KޯR�(�$�!�0衠�z?hk�����נ��IQ4�n�������#��������&?�E_(�ǡ�7�7wL�i�����/�o�M��ۃ%�pr��.��� �IY]�'�1A|E<⧞XT��lL�5�*T5p%M���+�QO�j|b���c�'���lt���N�+�5R0H?��ن����Ζy*�ǂ]p��P%{��P�:��u}�3�e��FY�S�����MO�����AI�b�ᶀ�� ����Uӟ�8�/'�+-�<X�a�Ɯ�Z�cd�
�WnAU���Oi���;2)�I`.هm�,�����S���$��K[m"%��=�M�PN��9Dk�Hr�
JȺ���s�]���Y嵌%�l�K�"�������W�S�nE�9O9�]��P���ei2m�Y4æ��z�`}1	�<E�LAz�8÷�v=M�\�����i���@�4�:ˇ����,U�lN�#��X�2:�]������-*H��	�>�$c���v�9B��*�a������x����
<Fԭؖ�HA�@E8����bV.@�6��=�t�O'���|���]aS�m�l:t��	N��� �U_l'���ΕJ���}���)���������IFG�|�-Z�3X�B�����
gT/v�u��p���'�Z���.�u��}��q�N�D��	Ѡ��tw#v�vk�$�J�R���۷.��:���D[U��岦�Vz|ϗ����_6�NaJ� E��Y��vz,ߩ*u�8�P�����EZ` S!j���\`��/NH��r�y�k�b�|>+����/��f�}�;n�=<)��!(żc^/"�9z�kd'�j�>�Ip���)�PĞB�4�.��/1�����ٿ'p�G05V�F5��՜�NY'4�f���q#��A�^�}C*�,�>��6�����U$�/�e�y"=&M]�<�ᅥ}����RN��ȯCJ�H��Ѩ`\���g�%�4J8���4��=��V#�3���_a����M!x!]����
<�ܽ�anQi���a�x�֡b	*&�P�嫞 <�P0dP?0"}����Y�ڊ\vѱ����R�E���>��1���e�(j��I����ʜ*��8@;���i�zj *+�i�X�C��%~��o�Ƶ�ᛉ������ϫ��&_������/b1������m�S���kUᴴ�\�Y�_���~��Pѹ�Q"��l��� {9���k�W���d�`�B��:��!^J��V�/3M��6����72�{\%������I9�+����i&2���#z<�%�;b|���W\<�?��o<��x���ɜa����4��_�KZ��e�I+���X�o� t�#�
�5pK��h�Vm=l��xi1)�J2&r��� ��_j���	ݶ��\X2�O�q$�,��O&d^;��'��`�Cv��ܡ֦�iSa�{vf�[ds�}�0
��I�Y�'T��{�oaч��
��ѩ2��z��i=�X����2!^��]7;5��~���v�C��0DՕ4��8�,$ԦM�c,��+ BA�8�!�ԩ��8a��tI��J��zU��R&�@�F��s�����0r7f��F#AU;S��u��p�d�d�_Ҽֺ�͇��b;��&� I�vYX>s����9���Aa���N	m~$V6�h���)�/h �@���ղ@S1��i�/l#�'�9h�g�z*��/��|wۆap� �˥V�*N�?����n��no�O��fm�]�M(�H<�W4�w����xY_Pٰ��U����,!�9B������_�nI�ܳP�}a�TFє����DV��!�kY1����]!*�b^�C��k�͘L-w�}�1��"tLQ�x9>᜖p�>�8I��HJ_�$*��V	���
���{�6<@�,e����M�Q��S����IZ��ҝ���
~�u~d�_JB�=�8fQ2΁qF����C*q���� l���H.��ĔS�ʙP���`���}?�F�]�R0�?g�K���p�iBG ��&�ͨ�c�Z��>5�\�X�h θ�K�{b[�l�Fv�j���p�FF���m�nl�8n���qpD�놚Yln���L U����|����z�$�n�m� q����==N+�[��2O�5s�=�KI�z��)���L���G|��Ї|<��0e��kQ�����^���2���B��Yq;�q�Vd{����NT|ݩ����#���y#f�ٖ�ŹL�����kY����N�����Z�z����g�z���~�Ⱥ�o3.7~�8�w�|���e_�ux0�BOĞԂ�������cY�`W���	�t�Λ̝��&45@�*~T�,˄��R��TS=�e��>�Ǘ��_�P����~>���>9��?���jh~%u�8����r ʰo�������TTk�W�2[�dh����,��F��8�nO{U&��ջ�B�	�y��mM��6͆�߻ru����1#L��4��:��0���6Ax7��l�q?�U��)�.I߅�S��w���>���Ü�7{*6�.v&B��&H�`�w��R"m�W����9���w�!I���ۚ@��ğڎq7T�Tnc�;�G������a"�:�#�pt�����@݂����#>�G��@9h+�hi�ϻ�EO���x�/���	�.6L*F��Kmy�a󹭈�G�}���6V���km{՛�Q^��C�r���E_�pb��N 2��%�
4m���TD�7�S���r8�R|�˿Go`�����
�E:����][���ڸ�DKi;r��\�A�_Ԟ���3���v��p�M��9�U����XK)���f�澉f��f��7Ou6�(yX���[>��0kG&�0���=��2$�w�kP�g�Rx�:X��	�K#hn3A�X�c�����	��Wb]�lq�T��`X����K�n;Āy룼t�����R&aGX�KkO�iA���Y��U[D��Q�b�Zs-�>b/r��սnd�X�g�g-ͬdAv��P��Z�N�b�S(�лW	QxXOpDq.����p�	�¼�"�B0�>n�yiGw\�"2mq" }hЖ�e��3e�}D�вi���a�l�:$����c�$�W*�0&UJ����e&�m;!~�nX���|���������z�G-�0�޷ �\�A,��C��{Ę����t=ǽQG<8��<���`J5~8mDpw��}�w��5º�O�n�2��R�~�okF�����8⢮�ע߭Lj�!v�8�`�����~�Z6��c�hڭ~= ����9J*��1ޙ��s��*'�͎\a���Q5�8�>�3N��ˬ�a4�6yª��q�(���7VTq_��Z���Ќ��r�؛R� �?-X~��T���
⽎,��]ܶ�iiZވݢ�K�8����i�5S�7I�;,�d��f�3�n�Q���w��N1t[B�*g�z 8W�B��:ߴIϑ�kXt�|�5ֻ�-�	���}/�*(Z��>=�&@��}���a.<�{3�(P� G�laEDk�"'HB�[�i���L� ��9pcp�}����{V��sL�G��΍��uf���X���lg,�x'�	-�,����Pf�ڤxM�P'\��{\z���`#+G�)o��*�w�,����Wby�3u�sp )
��q����5j�xm�o�/9�.a��R�W����L�"R;4��50�-� ���-���)q�D��j�݌"��
�����PP�=�O�h��c���ʽU��"f����?9GD����?�|�Iz�������� ���]D:�)ü�	�V�X�Y	�-HK	pϯ��j�J2� w�0ت�)w��
mD��Y-Y��d�l׫�@����#��Yj�@m���14S<%�?S�wA��U�\�41#=�l�ЀL���2����*���Ri���f"�B��G`s��L���%_j�FRE�&�Y�� �Peq'&`Ĩ,~z^��M���(�J�z�Дvl���;!4$������IX�穕䯱��뵜��,�o��g�"���h�d�����AĔ�/��3c,y�n�i�fUH1p�{2�,��C�p̾�Á�Dq7c���J��,q�k��.G�+p1ȷ�#��N�#(���2+��譿p�_3LB1[s�W��
�g!�T����q~`�ڟCp(&�����:��̱p+јe��,?��@�?��s�hIb��z���� �5�(�(:iJޔ���)h�ћ7�v�,�ȆP(���*��{Q���pY�߮Ȇ�lq��JNBY���pR���C�5��X!q�W�� � ��q��^:��ͽ!���q_�'���O�-ͼ�>\{�Mv��UR7�'����<VF�E��f�qS�f��F��h�
[�a�Nm)�͆*�@�=x�4��/e�2���{�)ڙ�&�*8Mqq=��.�X�����\b&�uA�~�3:��H�rU*{ߠ���p�ƅ��м�%ɍ��+�[���ҵ28�u���G�����rթ� j���
ܺ��Y���1i˹HL1o_˾ �7t�b������nC\��i�:�_�ë��iH!�ap �@6i�u�xs>�z�Bg�(�$��x��8�P�c>�i��������^2c�#��dV�F� ��]�L(��Ue�NA6՛��9�,��V�n>l�p��:���7�ȉ_Y�V5�,Qټ�ȡ�"{6_+�ER�_FH������M�]kJ��~��_�E)őJ�1X�>r���CD�`�J4��M����/e���& ���9^y�Gz�GJY��i���v�7��)��Eu������04���r�@������DKO����}��~_�qW�'\��w�8R/��O֦�x�Ύ�n�`�Qsˈ��*��clK��|E:y�QAT���j��-Եȝ�~ԥVr�'������%��c6Cƹ�}�M�X�Ȩ ڏ;����i��!�E?D�H
�O�PtP1R�(n�P��Dw�x�����4з'�#k�=��|V��R;�ι�!�4���Dq;"�-�q��*)��gwi���rX���m��c�t�Fs��߯,�B��՘�c�^�&¶�����#g>�D��ʝ����;�P�8f$��P5Ap{;�7:�u��=��L��}ck�,���!`�,��k��i��l�a�W��w�D6����)�Ì�3����}�wuKc0��j�y=�p2��F�l6&VȨ��6��!�F?�R'y�շ����.s��XeX	�k*@�b?m-g`b���7� �,��UHD�⚂����j���m���c@��\(��K〾�j7/���v'�����kUD��-Om���o��r�9��Y��@�b�O;l.�ޏ��,��oe4J�u���2�� �9>�m:D��n�~���T^����x؆��7L�]�!м���ȐVs�~�,Rc��yA!�T�f�Q��Y��<����	�|&�'��C`=�RϛOtB�����-vVf7���(�?`Hj�1�+}�$EX�l]�V>��b��zQ�B��(o5��-�_�1^�h";�_����=<492���R�5��J�b*�~��JO*	�4|g��ĉ�hKu	��l=EJ%_̒�Uj��݌�����yl�u�9d�������E�\\a�ܬ�bE��V_>��h�Eƾ�).��U���U�Q��T�⨱�-��g?�#<����ҷ�|7l��@�-����D�������Y��=���Sj�;#M��f�x��
R/w�\���E���%%�D�Z�n^
��R�k���I��4���� �"6�Ǜ�����_���JF�l�1�[[6�׈��8�dߍ��C(�����+��dX�F Ce���j�FJ���tk?���2�u��u�����M�P����
�0�����&b<�?pD;�Q��΅N�{�X��m�F�_ҟæ��d� �C�+�75�F�Go�94
 v�<&x�§��EB��s*��폃g����6�=`h"s�A����S`P�x�m���1P<A1��o9�����%4��ibN�
�B%1=*��T���o����@i'c��x�3,6B��ԤQdX� m��P�q�l�B뒯�}�Ę�_���@*aO�#<B�e#�AY�n���E���b���݆N����Ԛ����\�d��R{�7��Qq˔HN4�����/k�����P�-ά��uai;�k3��h�����:���nX����7|�r�+toꎷ�O���pS���荛���¹C�.���Ֆ���Z|��+O+��gȏX M��ec#f�&si���wV�8.�n���ېH�Z�u����Z�H�9U��2����L�����+3�xly��"f&N!f�v�/�o�.(��U*����Z����GeG�pt6m����8J�3�ݰ��D��Sgm��8�frS�� ������<�7��+���*�y��x����,���k#Gfŉ\�4�Z��{�^�)�֭�Ý�����{��`ܞr+0{����fPR��z*^�K�@�{�s���3;�v�ga�%�RHrh� ���LS=Lz����͐��Խ�h�r��,DE��B7�ʼ[�EB<q�C�I "B#�7���n	��%�Q��	YŘ��z|��T`D+zI@��5���9��\Ί����F5:�8Ï���p<����э�^�|Y��+�dJţXЪ7����%����>���0YՁ��W���fS�!2+�\��Ʉ��Z���܅`�.G+@��,�����^.*I�hL��r�)` qlK���<����~ �.��|R*���D�`W�+2�_� ���ʢ����xF�3n��Ȳ����)��*��L����W��F���a��2(^a�}^�*�a��+��P{0Ю�k�ߏ���5���{�Y5X���������Z�iazY���� �]%:#�kU��Ei"�'�t�U�'\e>Z�I��&qZZ�^���%��Y��&C�T�܉�?	���»m��X���#>G7&�y	�_�uz���K�����s������B��mx�Q�j��#�]Ig�wOWϜ�ͤ��K�R�ю��om7���E�b��$��̢�HY�V~����""v��m�6��z�CZ������w�"k�<~��$~�(��+���/<��dJs �q懗�̆Wx�%,p���[e܈ћ�#��/<�[�� �Tr
]�������
G:|�wS]�-`���z	WэG��)�דc����f��=��de`�,O��P9,�?�r�E,�qH6�l۔�tG���~�!Q�����(��v=�Q���'�!Kθ1;K���$L$�1�;��[\�:�:y�)�\!Z����Iq�F�ܚ�h�8�c:o��j�x�/2�2��)%�_TC�Y7���.����ۣ�y��k����Jۛ�����d�RK�!��TX�4rxy��K�' ��ѱ�Ϣ�h�#1������Jr�ݒ6��L55��x5Gr���@Zbؘ/�O�φ��W%���g��˭6��-�w���lk���� `�����a�WX�o������k��ګ��5��R����+�7*{�_�C�fBZV�9ԕD� �ҴY
������~cT�n������$�M��u�0�B��{����?��΅Y����E�e���>�:�+�g�Q��Ӏ��9(1@mk�>�ei9Ԥ����tuCS|
�k�]�OK����/�5�gF�!�ᣟ���$��e(���i�'����BH��ϭZ��z�4h$>Y�m^��1ƥ(��I�>#�ĩ��L�W�Oخ窮eY�Uc���i3���{i\N�/#AL���O���X�q���Ch��;pP������Pi������?�����V�ɟ&��"�K��7�G!5���B�Tf�	�a��_6ѣ��3���RӪx��[PX���T���dt�˓le��!z��1	#�~eB�jO�%��L[;u{w��dh1��E�^K2���N��Z8�\T�V�F���B�c�ؗ��6F�����QM.o�mAu=����6=^���
V�)��Ǹ��~(Vޖ�4l�G�R:m���޾�7�	��zѶT�ZU�x0����sٕ�����M���|X�mr\�ѥ �w�>����2B� W��$����m�{գ�ց���B�k�E��{qD\P�̲8�ܲt�	,�rH�BiW��������Ee���������"��u�[�ͷ���&�l�s�.�G�RF������=/=f����D��Z�u^�)��_(��a[Yڕm$�V����8�9�lՊ�h	\�v�2���vX����u��7(�ٵ}l���o+����������|�(�e���i�H� ��c���ѓ���	�lE/i��K7��(�q���l8�p6�6��Jo��G� ��t:��;wpIc�ȃb��$�y<>�?��Q~g�x��Qy����1Z��'��,%�Xtv)'�f�&�?���Ȉ޻�����K�������	쨶��͋�1t���A����q.j5ŕUV��.�o%͙	>��ө/z `4[�Ɓ�s>ԝ�?�,�4O<5�y~�S&�O��=b�O�}��p��!N�p�}F�-��sw�2���L�l�F8��E =m�G�Q�{��2��{?�ф��;�k�SL�w[ot8�OEѰVЧ0��D}~Ai��<�`�t�QF���ͤn;M�Ub�9��F���~
6]��!�S� �G�v-
_5la%�x=0�93�ͥï]��7+OBK��ߠyc~n����L��(c<}�q��ɥ���2I�9L��Ɓ�ϟ?9���lY>����A��aH"a]k��"Bq�W��׍#m4ΓJF�\7�xFW��zw4���������� f�wN� @X���Ff�� w�����å�MY7oC�O�o��Df��s�I�Lk{רטu$��o�I��P/ձ-���t&�<dFg�]�kj]���9!/�}$�3����s� �����{�x#(Pȗ`e�;�V���{��H�͒��D�#��!piy��l6O&��kL�0��w�W��$������"��i\�B�<�!h+�h�_�y!G�y��a7�5�v�Nrv2> �pga?�!l�(�P_��<��Rr�Qot���h����;j�G�k)NS��r 1��q�S�Y^����v&4^v}�����[�ԕp�5�� �4���$u�	�H�'�/�*~O�f��(�
b�ϾL�>s�h�E~��p�q0 �|?bϮV��=E라k��������'/�x+����
ͦ�f�s��`d���L�R�O��N�&����� `1]5,m"��{��,Cc�۱�'=j������Q|�l��A
��g���ķcK
2�A�4�>ps"�N$�|9^��$76a.)�?E��-<`��� R�so3Ё�F�=ȇc��·&��/���|� �3a�+��<u;�.F7�� 
[	j�<w˓lY�X��񀪁����߫�[d�TѪ)Nĩ~��U�g0��+��*�FS�%���������3(Ŕ�kѫ��()2U#%|�6[��g�x�E.Vz���l�C�<>�$�ڇ��� ��|�E �;ɺ�o5�/?����#K�����&7m7`��a��/-��KI|�Y�hTvz+_�Q�?��d���ڊ�f�
�U�a����k�~�czl1=����q�
>M��@�����P(���L?��j4�G��(�/(��
Ò��Z�|���J'��B^E��E=�g��gzMJ��X��\#�,Q��9H�� \E���1q�c�BZl�_`w5K���Q�a�FK�d!Hw��p����i�1Ѓ�P����m�௟�v�[oY;����a?�I���ჹ��8yۘ-=��6��5,`��Ä��w8E�Q�	?h��QL�ǫ1(�ֳ7�z 
vu�J��K��Y]/��xů�jJ�ze�D�xI7�v��v�%� 	4ة��n DzƑ�(l�%���z���r��o����{�v{���9�&�4%Pm�~����6!ęu���A\�1Z�ݵ����Z:��HH1V!�^
u���X� �ܪӱណT6�q��@࿰_��r�� ���pv��L���ߊ{oi�VH1e�hr��N�~>��,����SM>�w�ƿ>.�;�I�y�D`tU���H�H��r���͎Hu��,����v��g��Pg�������<IC�04բ���\
���i�����&��x��O�_X�Ƀ������E�5��ģ׊�-Y���C���7��*c���9��w�l�Y�9�D�t λJ�����~6���������'D��i$�h��O@yt4���9]��ƀ<�y/��0�y��+���y��Ks[o��2�،����`��b��H�G�`�/��H<�@��Eݛ�M�Ny�7� �B�B�E#�7BZв}E�sVR?�C~
}���1��s-��Y��h�Il�y����bK��	ۘ?Nd�����8W����K�扸���̐�w�T�3���\"Pj~����b�����^�ZF��x����mL��P`|��O���%�_#��}�O��}�h8�@�5>���)���Q�0�7W%����po+�yz^S� �#|�{�E�%�N�G���I�T�⣧2���x��{e&�r���SqӱXr6ũ��U���W�<�pE��\?4��_5��@�e��S�:)�;FĨ�s�.P�x!��;��~�G����>��_z�����+�!�7�8��ß�� i���W�m75���Z��|OF�y��(��� ����gE�uv�p蝙Ş���Ni\_���9��� OĎ.�5��k�:��_7DX��>ӌ/�)�3>�ڷp6s�~�m����Q�k&�v�+$���~�BN�vMცJ����^h%�sG?�.� zy���-�k��b$<'=3_z�W"߃������n�;ј���Df4��>�@��7w�9^F�B�Ν�p�|�!t�B�Ff�7:+@�2A�����ro�����l�b�S��KM�]��İZ��~~�b�w�|�>H�C��]�����	�!a�;�8�H�T�R�Y���[���1ߍ�U��k� ��/v�'��{��k� k�&`�ʹ��kcU��W<�S���a�m����/[�m��)~$vf^r��������S=�-![Ʀ5��EiW��Z��P¯fd$O�4�u���δ
�`h�J�i��l��������!)O�`dO�H�HWY�R竱���hb��}��!�f�qVP2��b<�Am�$�J���ұ�����,Y��b&�.%�u����rc1�H���E�N=5R\�{)��+��ՍkU^�������l�5����)ܢ���>��V69���&P﹓?B�T+��87��eJ�n���u�RCi%j�{�$��C�@ Zo���9|�ř4F���u�{���mv�� �o2N����y����G-�.���
W���>o8ߙ���!"���puJm��,+0_��m���#��Á>�e�O�r��u2�M�nޓޫ�$����c&kR/� ��Vb7�hb����d؄X9���Y�U?�q\=�|�|U�:���4M�6ҭ����gc)W=J�+�F4�>r��	�e�|�����T�6��Dn[F1_f������`���g���u���.�0#� �a�|L�Ü�դ* �(Z��B�Z�d�T$ۺ�5�l�q˟�N����;�=��@��5��k������ ]�ngw�,oܯ�K�b�>/7n#��lF�2�۠1�F3���OҀ�urq)�d6���_�Ɔm��'ﰩ}/g>ChG[�N�ۏ�"�۾��\�wڻY���4����(�xٌ`�$DH�F��,�VD=���3XG�t�)���D�{��--!,^J�<��W1��� ��	j5�������
�K\�w���A֥ߊ�	�%So8�ǣܩ'�:0i5+~t�{��y��#�ݳ祏%-E��_.��]�q��7�k�E0-(�Z���8�ͼ�5ٞCE����QR�.^/v��?5{�\�N^��󘓨̩��nN���X�
IĲ�K����?�<����"sha�)F.�`qLGX$P�Ր��ߚY)��y���1w�/�����<�w��mk�3n���x�-��v�[ꮛq�2
붔�n��p<�bw#�(���M��[и����_a��d�������o��゗��s��l��8�V�'�<���5Q�}�9��L��z{.`���4�Ä|�{�V ��ۚ�R�N���ݷ��ZMh��<���`4MGO�{�ʰ�ʯhk�9�<5.�{�V��o1�I!�F=�%!V����A5g�X�b�	��� �R-��񬠡]��[�9�\q3��,��A��v=r���)��3�S�Y���=H��׸�[�L��A\ٜ�)��>0Vp?�Kҿ���>���}�F�:7V��<��}:�Y�u]u�]kj��"��q>p���-�OD����*v�E�m���n��l���E0�Z��pCxv��Wur�ې��d-��*v ���)��F����3=�鱞kd�4�	�ϭ[̰J8 ���z�F���_����;���n#r]���B�
V�n����\n���#��nـ�1�	�����O����+�j�#���ֆ}� �u��l��-��udsy�Rr@���ܻYc�|��/&�����G��6g�p�n!УU�qg���L����	*�!��m�D�d�u�|3v1���'�C������J���mo�B`������`p�#����]NK�B���t����]7O�VH��=0�Z�����B��W��!R�QIV?�!�g�)#�W~0B�OڝծY6%Q�ߑ����l�Is��>�O���=<�tI�6Ϲ��{8/Az��J�+�<Vc�J��n�`-@�\��k� c�����P�����QE�֖�E�����f�j�߮��S�qo� ���g��AV%����o3q'���ʘ���ŵFp����񍃑�&kN��\��dǣ<B�lG��3B�EK��F��`�V���V%9S�i�B8�/��):���M�s�6�'��ۃ�L��̶ރ,Y��<`9��IYOw�:�a�!����SƑ]t��5/�]��%!�<�PDCTyX��e�	�P:�y��$�Sy���fb�4;�'�*^ؚ7�]�J�U��f��0��@#n�1xf`�t͜s�q���a�ʸr�=�m����O� ͫ��_�t���ۡ��@�0,�筬S<+�L�H&�� �k*�g�]�����V��$�+<�?����]�+�v6SB�'��{a����uZ�8��
#�ǲ��H�u�qz,0KW��覇�-z�H�`���[�Mak�9LmDA�����Lu	�G����⤛I>cہ�p/ħvT6��m�@␜�CXpsʂx���0x!Ňv�˷�XȬ�cY��ؘ�P��� ��8�lȴş�=y~*2������j��!�ׅ@
%L�9��V��̷�K6d��+��&1z"�x��O(�\���!��N��jS9Tș�ȯ��:]���g���{�	==��g�O��j�wհMD�� t6H��}�*W��<�D�2 w�_��}��[�3�u9����j��Cr��1���R��G�ߣ5V�3!���-���6@�՚A�<�ݥ�����D��̰U:B����M�H��}v��O�1�� ��]�8���䕲�x^���9~��_m�}��%��a���������V�#7��F����Qǅ.��������o�ʟi:�I� f� � 
��6���3Q_O���y��E��zFlZ��XT�����J�xN;�x�)eY��1C5k��{��a��`DWlq`��ф����1+x���
K�㭂�>�4�?�5�T%�VUҜ"p!�Wv��2��(�P�/h�â"�~9�������Nw���d�G��^��b���@h�a0�u�dK�&hR���k��X�����ɫh��B�+��"�?�>@��KN�&�Y�0a\&������u�F %v��F��tϺ����haP��N%��Xf(�&-S����$Ɗ�&��m}c����5������p9Km�O)��Ff���*́��o�����#�sj�^`c{k�}�Y����_�������c6�~�"���md�!I�~s	�[G��#L���i#��O��3�>ؔSj\bB����� ���]�,��c����z)�.Z��L��8�=��$@SU��ja��ު��XyF�>J��a_�s.�~���r����6�C(R�ukV}Aj�%
�))�򚆷٠F��F�;53�O���M�t�ockbN�B~B����T�C�d���+�
��?�$Xd-\�w�)����a�1�R�	�ޝ>��|��T�ӽ��=�6F�p�!�_���xK�,}?��`פ]
����䟖�c\���й�%��f��v�p����Їa�A��)wV%���]�q�R�����ԛ�l�L��s:(�
r�h�bR Y���1L�������R$��[%1#.K�����t�A��a0��~[�u�V�F&7�3�z�,]'�4K�x��Ŀ1��]$	���A�?�ζr�(u��<��s��,��t��>����n�0�ǥn�SUɩL*��;�_g:��Ð+���ҤcCh�tjB���3��e�;贛Ά��GϽ�	�)����K1�$Ds{��u�
b��,^��D�R��T�f�L�΂��?t�q��l=�%�k��'�ʢ�"G���~I����/�JH�m���u$��͎	��kL3p��������xT� ó��l�ȱđ1�i($;Q��Ԥ��`�U��o�'��&�n�-U�IP�~�������{M�1�Y��,`E�I�V�	�"��z<N�8z �$����I��C~�+t�:锱�F������p
�^ņl�����e�|B���_����)+�8|q=�淸�/�/�1��fK{��ygbF����
��Vj7�Z#�⿴5달(���Vt[	F��
����4���l�� ]e�1L��b�6���<M7�a��!2�MC�7HO:ao������ᒹ�MW*2�?X��'Y�U��G�p�N�(�cY���s��Oo5�gOD�
1���]sG8�!�e$���t�E���y�ּ����zT���`�텳��rz��]f�BP���T��V=W��j٬d�N�Jd���}�;d �'�^�|u���8@a���u��X�
Ec7��M���(ξ�l��LS?1���T� H��-��%�S�M�㖍���PD/�a�M��)���@����յȓ�j�!�ۓ����.{f���9�L�2��'�p.�V�R���um)]�%��*�h��PY�;��S<|,G��mS$����Ϩz��xH������9Y*��
�aS�`���%����/&ZY���Ȼ.-�^� ?\�&%�%i�BF�z�5;<�gx��k�HV�����aǑW!��Hy����w�ב+�Go{~ߪԡ������^k�"8�����\�U�;�Ǔ�N~?���G�V>�b���o���C��I�d!���sW��&P�ɒ�8|8�w�����K���1=��u)�� O�Q{,�Ϸ�׋���v?�r����^)�a�W�Iq�O��`�M�w��� xw*�ZQ�^����j��(֤��!R���{������i$�[��.j�9�dp}~�6�8�`��� kk3��Pr"l'����@���#?�cSBi��{ڀ�L�hfq�B�ͣ5���h(I����IY��o�+ڔ�D�t��x���e�O���UJb�H&H!�����c��	
=������P�-P����+ES��꾗���;��厢�7";�(��ܲ���s1�`=ر�Qm�l=�G]��(��lң��w�c�+n=;9U|sDA�/���#3�prZ�-I�{����;����
���e}�M�i�f���(�X�E7�m��aG��K��7��+C�L�>�[*����_��[*ɡ��ɨ3�_��>�U���IQ��!(6+ޠ3���Vh~�0��yl�/dvqt�����W[oF�"�х]�]�M?o�|NP5����GS�]�r�ӑ9��dn
�p � K�:��� ��^�^���1o�,~ߴ��z5�l;oc�鮪!^z��ZD�'^�n�R����>�]:������S
)x��X�y�_�r��p7+!K�g,��#h�e�yf�x�_������s�i���+��D������#��{���
MHA�P�PiJ���̛V9��OhC�/V��{�HR��a�:��߅i��M*2��ū~x+�H�@�� oUk;��f"��p�7S7g&xY�>Y�$��Ҭ5�O�	$�7f霰 �d ��Ux�}/�������1<���iJm흣�v��ϕ�w�(��Fg�̙�uU4�1�X�Y�~t%*�_6�Og�df�ffg��Jl����/j��	�1҄�d��Q����hݘЀP���)[�R����m(�hHqǱ���apl���N���hJ��9=5���r���Կ��[��,a��r�#ϯ�	�&��4���su�hB�Q�{]����D�־zv�=���L�!2��)��m�u���?�Kc������UV���-��ۖw�:�ь�0��5��J%����\�l���،�d0ԫ�l˾v��Z���x��+���U�R`��i-��4�}��cj�WпB����n�(=���J�U?�f&4[��Y�G�c�G6�~5Q!:jN,�k&���b��}�[=�'M:+���*x@/��߬ЂkS~�y��Z���C�+�$W�V����5-S��=Xd���h�3�O�8�r���Nau��]����:�J��j7�[�#2�.��g�vưβٝ�O�I�=�.�M��	���"vU��#�T6El�>��<hu�Ҳ�=
�2LM�^T�H�h�Pl�$�$���bSom/��p���w�k q����ؐ�����d��M{.]S�Ne?Q��A=���T}�Z��Y���5LGY8r���+	�.Yc(� ���x���_$1�Z��?�N��3��4���U~��Q��C� ��v�Ė^FxDq4$�� 2��yW��.� �f�����he_��ϋR��}�;��)?
FD�{eY�Q�΂�M̷�߆���p6�\��(0��HY�'~�]qY�ޑ?��Ϊ�n�6fs�@�i��Y=
��yb� ��	�����Q+�]�!�x�,._>��_�K/�{@�Oܞ�s�0�x#�A��0�e0`te^�􁅔E����nQ���8��iwzV"x�d9�S�=��`T�7}C�P��V��0�W�l�Ϻk9�~�
��a�����ޛ.`Y�҉Ð�^ȡ����9�'U�.��>� m?��c|}i�QRW�$hH1�DZ�З!X��A��J��%�[^�8�KsQ����F7����V_~���^맰G�l<Z{�2vmf�Z����� ���c�H�����ǭ,U�T�
@f��)-�C���b{R)�i�q�0�VѾ��)zK��֗#��^	"�s��*��|Ԅ��F�*݁���L�ʙ}ҫ����{�'���m,h(b�I�^{Cm">�@P��'�k�\Y_���L*@+�A`�����]�u��>hE9T��Nq�`_�����1�c۽����7Xz����p�Ju�����3�Yej$�
�ϻ�}%׵V���sS�@<�3��=��O}u,��I���P	!����a��{DK4D���_E	��!f�~q�P^��[�+_��D1�)�K�v�SCF���E0�ٰ�!��E^i�r��z8��j݆jn6��'
������O�|}6�px�x3?'lp��(Jo6��H!�GAl�YeR���xx�Q>~gO��4r�mh��U�ę��̫�j�u��Dy�R�����@7��������#m�VS����b��'"T��03��J�h��T�� N��/V<uc��rL�yr�
�X��5C����M��~ݜz��jc�+7km���=���r.�#Gۘr*a�D־Wsن��Jm�5p�AY;�!�u�������d![��� ��*|2��a�P�x�SЄ����F3K5"qP,8��`���eK�^o6�>twX���w�8P����R$��!��R(�:ӳFC/�����@�?7~Ӡ�8�A���2�[��W?�1��uC�%����q(G��M��1����,�(��'j�/U�\m���ZW�C�,|m�cv�\��EV'<�ԑz����"2�>q�A��s�=�e��ܙ%�zh���i�Ϗ�$��yk��RO@��Nu����p�����^�Cּ!"�P��pz�hһ��ڭ��pRt�"�	�l�:L������M�����CQ��˹8B�^ҕ?�c�k���k�;�0�c6UY!h7si�C_���5��P�<�9	���n���^�EVP�؋.��\1�J�(6�n�o��s�<#�%qd~�S?��|W��q��:
La=�Jr;KHty��*���6�����ܪ�}��?�p�����M�.\�9�zLQf �K">���h�ٌ�j�"����U�������G���3y#ڸ.��'��G)Z� �`«Y��u}!� ��oK�N���;�ā)�@`�Ԅu���%^����lR�׎�I�|��0�3",��X���\
�Ѳ�,*�渒���)�䟚5��~=��	gc�#�Í�w��|�wU��V�c�1k�kV�~m��k)�S�;)�^������^0x�.���AW�,���@O��v�]���^L��c�0�Ѭ�YpD���	����p�,�|�s�W(k��v%�]���0f���"��p���̡uyJ VR��\��阮=�p�9�Y$��Wja�^���- �w�8]��:Y(a$�{'��q�;�/{�%�E3X���.�LG$�#�+�7�YF!�?���{<<[R��/Ђ�}��Jص5'�����0:�LQ����Q��2����e����5@�T��Od��.�1����^v��s�q���M�H|��#`��y�*G�v���J�7Z���*g�Ǳ\���6�?ฐ�8m,R�']3��\�����S�0�/z��g!.(7�;r>��#^b�����6@����P�ӛgw<i�*0�.���by�C7�idme��nhPx�����?>� e�Q�0oG��%�Vڴ0��'W,(��~�q�FT>%��2��Θ�����ᨁ��0E��{����ϬR������*�;'�@���`4N�~'r�H����%�\:��y\=�|*�V"M%B�D�͹;���f����鍾\0�"����tiڜ'��_ ���<�^�}����=��ϼ��6���l�R�U������� |����g�d`^���I2s��o�!�GI��a�dRл䑃Φ������m7C�9����,�da���f`�S.�:.� �� ����^t�e��3X�
״k��#��m!�'�%�Sݥ���^:Ẇ<�*�9�wK0�6�5����-�p7abW�k��1�F�ݠ8�FX��.6$rJ�{�e�jyS�3E�P�w�_`/˩^1��Af`I��+�d�J������E�����l��Pї]�xi�U2�GE])Р���7)l;cU��Q��h���\�qQZ�ٻԂ~��~o�1���[WwO�z�ܢ5��hǏ��g-%۲�z}p|�+=���;$��ǧ��/����r��\&>�_��:��������'�`f��|9�a��h[�ͽ��/�T��+�K�"�>Dw&R���9_=��V�����7���H�@f���7��O�
�5��ދӥ�� ���ֻA{��7��G�d�4[�'f��K���n�8@,���~~Ϝ�¦�#�6��wIi�t��ض����6H���2�Eؠ뜏[��(v�2Y�Q��Wkr��G՗2!���$��rp�ϓc��>ѓ��9�,Q��<���i�R@�V��.)��|�!��M�W-�n�TRY��sB3�6�fg�w�\�>���o-.�Hr�;	ҷ�(e7������C���Kv�	O����]qI~u�c��;S��ݢN�1�띘��2�6�`��r^SXx�%TGI��������m-��s��Rmx��\���&]��p?������WW�3k��
 �b��A�[,��#%�Zyo��&�8�=Z����4{>,?���=�g�k?�;#N�ѾZ����0m|�@�ʺ�&HJ�b����t���x�Dg�$��NLy��[ K��P��Ij����v��lQ����3,���J���{D���%4G�`�GR)g���?��S���Ht0�l���i�	����4E��A�-W-�;1r��hR�t���o2S�����S�iqt�
��I�\����$��l��OhFF���U~��|f����MKj�K5K����A�L��N���0 Fa���6�燚#pN�������C Z$�q:�7�(F&��ה��ݼ�O�~kQ���LXa#����s01'IPJ�ñt	�[Z~���95�vf��A�c�i����}Ӭ�I|�^]�CAR�p�j�!Y���d�;��]��m^%����Q�(x������Ѽu)�I:�*����:�˖�ծ����H)����:�Ӵn��&Id�{3��V������X��]�����A�Z.���Sm'�.'[�~�)f,���џj���ݬI� x6��{���sReP{/=��!�������C*���'>yeq8?�0X2��<�#DK�D��Uʱ�&�ͼ>(�N{�*��JDAU���*T��a�(�z�~Z�b�-��Ks�ԏ�++:���>�W���钛o��+A8�j?��0.������r�8B%桄s����4_m̬^�gm���D�tQ|PT8�z�p�I�L��q�k�P��Y� 	uGL��Q.�-[�$��O�K�%ߐ���p�����/�H�:��ń��;Em�Mʤ��n�fօ���M:!�h�ߧx[�]`��(T�k�ז������W���)�( ��J,K��sG	q
��7�=ߔ����S�1Ff��tD=$0���Ι*�,z�0�I��y#T�;&;=��mr=�����w�Q�#�(�U�� �j�xm2�����5���2�l'`a_>��~@k������:�2�j�p��}�]���@��>TPV�[��%��_溋� ��������#��rN����;��n��$TD^�"
'�,�K�Kl���^3��:+����� ��qgv�吤I�nI'�Ĺ���o4���m������������ g�E��-�� d3r�D!�xX@�+��wS]]�mm�t ����(� ��C�z���V?�ݽ߃tC>j+/�ܜ�깂B�-����Cg-�^���2A�a��ZFs���c����dy�[q
j�g�e�����F�4�Ψ��\
2ee�M�ֵC���y3�ɼe��s�����ڸ���}*+C�7#5Oz��Ф���&`�U����֘��p&�r����Ǘ���D҇�+}��D 68�>���HR����/%�N��	�zN��B�!��C)z�$�I�r�^m��
|���E��R��X�z�u�H�	���\A���r�1���Q����XB�] �ZBV��U!Â"h�
�Ύoc����ߊhz{���z�����CZL�QI���'�p�w;|?'9�ۣR�E������n�0e]QMm���z%�U�BM�dN��)6sd��hht�W[ښ�$Xe��2��&�C86�b�&<�)��+f�sT=�\�Ȕ���H��{��5��H��]db�	�9�C2�}�.��D�]����Z�d��S��J�~�I_�PލIU�c�4��_Д%����.gz7�/V�	.�t���yT�(�AT]	�&<Z���T���!��U#�ծ��ug .	�N��^�\C�0Rɥs��n��¦,�xr�R�X��W�)������֔��T�����c�OMj�H�� ��\C��G�><`�R�g �f]	tU���#��c�D�ڙ(�o�g������J��;���|���5:�F�:�)�Y�5�3�������f!�Z��2�����Gqo:ӒngщɡR񥼊��˗��	#@��ղF>�7�.�p��~�p�MQ���v�B?���b�,��*j�AT�g��JO�Qd# �˛�Èo���<vi�mh��.�Cf`|WK��d���p�`�Ĩ�3+��!�ybQ�]a��	���Y�f��8�fe�UW�9���}�Ҙ��2B�:u �����/��+΁�#зQŴy�a�T!v=�l
��_ ��'h�mv�E�q����VMy�V&m�ȏ�#a Z�8[��֯�^��L���Daf/\�io@��^�VÅ�|�|Hn�"�gɕJH��Ֆ?���p%kE�SiЩ��;D��ٷ"V���p�"Vye7$R��Ha�0�ī�~��a��W޳/�ď�ե��Չ�-�.r?\�V-�������ty� m��@�=�F�d_3B�c����.���y�B�K�2���i�F��_p�nG���8��Yy�=M b�V|PL�C���p��u풎��/a�6h �����X�]3�8���gd$���|U�Ի�R�\붡q;�U��*l><\��F�q;��;XHzS<�Z��R�O� S�z���6���wo�Y�s�{p)�i�\([�+���w5�>��fo6zj[��*9�;W��<���T/����3X�Mq��)���Ti-�h*���de�@^�uGV���g�E0)X�t|��fHD��pؘ�:#ŵ%�2N��o"a�osw+��q�h��@?��0��fvf��y9������uܫ���ܿ�*E
�<9�:�Q!�8����� �����kg�ݮ\��FL�F��]Htz!:;��:�j�tl�U��{����K4d`��e[�`����z�m��Ǡ���H�+B�%�z�w�o��/���ϦU#9�Q��F����6�kSd�my+��z�	c-�]ڬ!��F��bK�@#%�v�U�&�[Պ��΅������B�E��`��	
��PW�/��.����Gy�6��7fA�f�/>�P��	"9�)F�^��B�Ý�$�a�k{�Ò�s�w��Q�@q�z��no���g��&�ߊ_2���G�3�8(�R��?!~C�Ө��r�ѕ£�xdP�R�^ 3�~���S5����i��������X�߇��%R�~Ă�n���ͬB�ͽ����*��5��@2+M٤�'�f���Yo�-X�;�� ��Vw����Dv���˗�nLo�M~����CA��ph���-0c�_�s#=���.�r-v.9�u��LL�Z(3�F�]��ө4у>f������[����z��S6���R��=�??,8����	�SY��7Û�Ƴ>%�x�!��oU8L�ޔ����w��(#�D�Q(� ���I!ᄾJz�����<��7����,�]8;AB޿�r4�/iĄa�Y4)������ɉ�1�]�%0��K��Rh��A�S�!z��i�0��3�}�81Eb}2�@n�+a�q��m/��P�1
�1�?ٗ�	�TQ�_�A�]?/��H���J��b^C�K��ńV<��3������f���ϔ�����}��n�G*��w�Q]��{Gi���?/*��:hh�A��T�_A�m@=$@.�S����Q�Q��l/d���s�i'�ɳm��ʟ}�:ޖ9\�x�YA���~�GE$i�RA� t���+)$��=�?Y<y  o��w[>����^��t ea�1����W�0~��0=���0L�ߴ�"2��u�ZAŰ2�������4�DW�0��㦒������<���XM*�A�>��c�FG�%�������R�������&��fn4~b��	ED�q�;"|C����hNμ�	k�;I���0,yx^6�]�z�>��X�KGu��Y�ҷ_|vb��S������qx<����vd�����n{e6�f�G#���ݤ�����ӓg�$t�e�(���>��BuN�o"������o���c}����j��blX˻=��c�J��c�أ�񏊘aơ&��A|Y�W�ݲ�g�.�=�o�3c�w��w;Hɐ��cPi� ��R�6�)�Z/F�����>�H�ju��L�rӵj�~rW}.em[�>���X-�1�eox�9�!�"0�c)	�:q�	��ٞu#O�A�`�=�qI�#�>�*t[
����-i.7�*P܃P��߸Қu���d١ �`/$o�G�x�vC�T@J�Ǭ��i!.9����	qMc+>Ή5�G�V����9����z�~�b爅X��j�#��o��9���;`Ry�w}��G�T�h^��|�^�ߨ&���,��<����ig��f8��C(h�/�
�mѻ���I�O��h͌ҙ�ܱ�}X2�YYN��	`!���Է`8�C;mn��r0[ygsM)����9�+۹�Xg,3��,��j*;-,_�s&����,ý`AQt"߹�v����&���@�O (>{&�j�E.�.
�֝���=K��{d+���3O�������P�ST��?�Jp��h>��J�����$��{�y1]{Z<�[�e?p�L�t�E��T����ܪ��t2�����J�O�{8��μ��-�i (�E��a�z
~й��Z8�����ER�_�{��Ҵf&�L�/"+��n��/���G�]k(���G*�w�u���?�{�o�@#A�\5ϯ�?:9���#ڃk�,j���2x�`�I_����FS�}��(@5w��֒���L$����}6҉܊��g����(���̵IxQ��m�9 �v�kZ���m������o�{�
MX>,��$#6-}����g�-;&�
��翆!Odbb �Y2Ғ'�W:u�v�e��r|�i�o�^�0��q��I�Bi��[F��-Eh�Q`���4}Zv�pg�!��$� $��c(1��-�S�9n�N�.�ܴ@'}ɬ'�d&���d�GUݮ�O�t��ʔx���cV8�,��"�uy�,����`X���1�������<�xj�H��:<5iM�%e�RY/C����Y/�1�1���B��̌�,'|0!��W�����P$��_!��B������F�Tfq���zȅ[��p�g{J��4]L�ߦ2�rr?@<�� ����p�ʳl�W�K(RK��Ů�/˞c�
��)ΉS�e��-
��݃�լ3Iq_�Ǣ���Ğ3|� j�ϊ̶�K3�P��0��6��� CB�F���B���d//��9�Y�l8�d�>t�.tBg���!�TD���.k"ܰ�@��D�q|]N��w��K�ȓt1��~J��n[�i3��h^�-�e����R��>ク)4��&à�O�
��܏����Ǥ�9���H#���f�Oz$ͼg���"� l�)�(�\�Wg���2VW�v�_6Lof�����R��(�(��М�e{#8 G�a߼��{&>��K��v��S����6�b/0��6@{Xo�[�C)>�.d��x�<z�r�Kw�G�jo�d"/�>�Y!�q�����eM�$ϼ�:�9�X��.e�g�k��X��|�˟w����#iE:���	�tWQ����MJ�@>���s.�a��eY6f�<xK��K�9��������xB樻)X�ۥ��>I��~��ܥ0�̻��8����k���/I��}7�� �`��x;9˴�i��Mɮ1� v�O<λ�
�v%�坘-1ڻ�o��w���� ��#O�@�����M���R	���FC�Ԅ��0"˚��eB�q˥����.h�(}�m��D^�8���\�庾�摩Ll�uE��b��q���
��C=�����v�O�����@� �@�'������,7)m��2�>I�O�L10��("%�M?���ͨو(2��E�ؤ�i�^��1���^��������bY ̓l\�=�2|�����.���{�+���]�@�^���)!҇�0���>Q��G"o�Ȩ_�5p�≧�9�o,�*"\׍�c�@���\�������u���n���|���d>)�huA�:w�� �r�b��"W0:Em��Gh��߆�A<s����F�R�~��ɀ��W���r�8ׄ��uz�E٢G��{x���t��'��b�}�f�=�H��������w�F�qM�l�1WF�@�߅��ėD�D��|_������7k��j�=u�6��t�a@o��eOҗ1ˢO��R����)�ڬ��ӄ1�j�n��t��Z�!�	�u%66Pͦ�~~��>�`�ƺhlc<O��]8��+��d�k4G�i�e�����I����x�A�>_��\-��K�a��\��?��Q� /h���b�������{�Z3�Ȍ����,�������#8���r�j��	Y,�=l��E���ª�w�m�md�'+��~��i,m F��pH�=����'v�����U9f!��v8Wf#^���j
M|)���U~�;���xe�#�յ�x�2����l�9��_�+Rѵ�x_, #�`!-&��f�P��tR$_���1�c��m�>�s��⮮ʉ��-�ĚA��ňz:l�d���3)6�7���SW8��R�KQ�0�N5�K��C7�BV�պ}S��4�zI���	�l���\ۆ`9�f�Q���90���a~H���91��53:�'��o#�0KI�tb �_{V� �[����j�l�Kj�}���԰��������F�����?�9	N2��z�3��^T���"\t)�GTS���I��Z�\������G �wGuI�����o�ƨ����1o����r�S�*��W�����L�o�v�r�{�zՋ���`m@ܰ�Dݘ���V�k
��B��j5��IoF�N��_�H�$��C�W
*MY���v���1[�*V��M�P����=�{q�P�T()��4�e}��ƈ�ڤl�ͪ*���LV�T���q䁴?�cO���c��!+7�c���E%�KXx���9[�t �m���9s{F
�$"KE?�)އ\�W~�ӧd
�5)�J�P���y�th�9��n���2�G �`�����_i�|#-�!ED
�ɤ��d��V ky�(�	$t�{n��<���p�� m@R� ���0�ʸ�J͒�k�˼{	���f�B3;$� 'e�.E���m�b2�v��h�O������{����u�&�
a���x��z�l�:p�VG��4|UR�'��{�*��"-PbCϋ�ggN)����j��'���X1G�Θ��/ײE�xiH �]��pݔ�_l߂=Ϋ."~W*F���i�E2ê��*X��5�*�L��\9�����З�k��}�\7�r��	���[l�`	a7��fk���~&��N�K�'�+.5'B�cJw�[Ҧ�)�iׁ�|u� �ub���be��弝	7�G�:��Qj� py�)m��I�X�r��6����8#���m-�3���o��Z�r���{��C,� {NRʻjv��h*�����c=������<)J�y�k���k9��Ct��H¼\�l��F���ݗ�85k0�7����u#z��!���b�?5���T�YY����%H�BInPU�r��������%�U{q;��7K��p��N\q�^儕��� �]r��?�s�1.L6M���0���ZbЎ�O��\���:4����Gx4��J���^$�RF/T(.R�`�?�\aa��Hx���6�Y���ی��CP�D�U����>x���[���/�_�t�*�Z�Q�o?9�_�1p0�,:N_2��I�^I��TIyn�綻k���E�v��Q,UU	��,��#5��5�:"Jxa{rj�uu����ޔY��F�~�w!�a��P
���O�vۗq�!��׬����O�v)̠�58�n�� ��ǈq�/q%�^rv�@��A}j>_v�v~�f�FM'I��@��ڧ�VZ9>����?�w䪜sѐ]�|*IT4��x�L�CS�fJ'��E�?�O��/6�/��so���f�75υ��X؀��!>D�k��]��f�u-�\�r�@X�:�z�`���O ��=�N�Qn��4 ����̣�!�<�9F�H����X��iM��;��Ʈ̛���v�%k N��!�Վ� !�l<z0�u]9td�FN;9��b72ȻP�L��E������U.��.�p�1��`!%8��G��O`�ļ�-]=+���v_kW�L�k��(v�ϕ*0�Hn]�U�N��������=)�Q�l�[^���q�]T�n���{h����|���[@�.b�ϧ9�{�"����J���3�;W`H�f؋���<�9�������;�D��A������X�|����O��Q����
��\��H]+�G�W	�^5�Pc3b\��ņ8C?�F�>7�"�������tp4|��|�w�ִ��B�i�M�i��:I�Ρ��Nǖ�$e9�6�&�2�b����{9p�Kx6��0���/�-�œ�9n�\�ĝ$�yb���6#����l/1�L�Dd��d1b@�䜇��Q-V�&�Дg�Pߨ��:�(���1B�\�'ɖWޡ�E��YB���0�;K����^�MBn���B��sρ��y�,��7���0��G���Ikˣdu;%'�i�Qz�l]����뷋�Jp���Zɠj^�z��bz!q���+.�����ڢܼ~�@������;(��[�+��*F!�R���[ �u��_�o�����T�>4/�8
���v3�� �Ȁ���P��TїX`\k敯\e���z�2����Dm_%	�b)������ �,�n�~b��<��Z3�RBQτ�k�OA�7��33�wۉir�W��pne6F��M��Kՠ��{^����%�[53�{�������JI�☟D�����Xd%�OP�!�Z�}����q�#?�8�GsT�eoL`E	�`�P*�M�� ^s ��kYk�5���װ l�ŝ�|�3�[�i�%�d!� qi\͝t�v}~�dog��^������.6�=5��-?�D+m���j�hv�5ѻ��K�����I�䐻����57�iGpL��4>�Y��k ��5�@�muf$w3�h�;uI�0��2X�r������B�\��We�Aj����8/rHl��:[ &�D�k������j�Ec���<[�#��K�rDR�����q+
�Do�-�n�"�ۡ?I�,RFT �9-�Jk��r���4��yFJT�B&~z�2�d=*���D�cj�n#͕b��T=#y'�4k�s�oZ��с��u��'g	�nj��8��P�:�w�HIR%�#΅��|���%܄C��BD�N�#�)� J����^!���XB�~�[A��.�A���鬖�l�V9����e�I�Ĭ���M���s���ܛES$��V�O��m�=��J� �.8:]^��J�u(�j�;$)��=���r��hk��B"+e���+��j_{AO��Zh9�tO��*C� � <�$�#�\Хu
�ILB{R{���GYF@��K�_�F����:��ksM{?��n����C����~f��E�N��$����v�G30|���i�>CD�U<�b�}D3,\"l���b�6�y��d/�b�\&S7$c	>cd	�&�+�1�>���5f�r��sH\�yNtp�j�+���~��-[���CȀ֥����φu��xX�X����O�"e�,�9�I����f��#;)i�si:v�`���ϧ�Q����k�}�
3B��J�l�c�=SJK7��j����ǋ�q��11IM�)]�C��V��@D���B����_s�1�غ�xf)jsB!.��u��4�D��+��O�t$��-o(�d�<H!�ӹ�cy��؟*^FtW4�Q�?��Keީqk��WX�Q�"�Cq+�# q��=��^{7D�]�0�GY�����y��ϤK8}�p����Tq�U������bW5��c#�-#��2N�gz��`��9o���t!M��דt˻.*��|�{^��=I���	BO@Ni���Ԉ��'7^��)&�j�#�l*>~��;R��i�3'N��)o�2(uT����̡K��m�O�Q��K��ycb�K'�ѓ�״d��`�8],�
*z��L4�Y��%�U�N�1p44Fs�:��y{�B�~���mrr�1C��S�8�~���ݺ�
ce���%U�,�7�A��b���ܜ7�	�A�N���2R8�}~Now�6ـ\���w�{��A��NO���|A���qko�@j���yh�LM2N(aCn����߀}�5��拫&ߟK��結�=���rKRa����طϼ�A<V����!V%�PiրG ط0�yy�3�����(��+Tk�n!�B]0�s�ՈɈ^ţ��!��ܮ�xXu`7�s�^�46)����d�a��U�l�^�B����&լ@QG�8��eW�'�ٞ�lSU��|��u�:B���>M#��ӫ!��rr��`�]��F���d����Rk��6�s�u�v�WA	@Ї��:�^p�Z��ϳN��kZ��t��(����K~�^����Ӳ	������Ū��q� r�gA�������u�@�*�7��G�2���7�a�2k�í)L�K�s>��f]� �.̋�*)N#�H�,Kϼ j%Dau��2���\�@����k�aF�>�(�����Z�ҦƲ7����8t�b�}�S�I�82�����B��iZ6�W&>G�q7V!�� �"�� �9_�|RcA�~��3j]I�;��r�S���N���O!8�|�'��re	��m.�ekȒ߫�ͪ�%�Bw##�g�����/n�;Q��x�k/�)��m��+q�=\�,�|9x�"4rlYXƗ���RN�����S�B:$S=ſu��jw�'k-��2�) �qu�]����g�N�������ƚ�u�U]������;��'v��x]=��	Y}<���q�w��C,��9*���P�;��&��}x� k�� �k�"W��	����I#F~1u�ӧ�̉��q�'}�{��!0����mB'g���эaN�M��7�i����H���h������9��h�(��H�m`��ZИhB�	q��[�I��`�tVxqo��y�� ){hQmQ��8XL�b��&Bf
%��țf�-�1�.��c��'�*��駽X�H#i%�B���ۆ�{��~e&	��^s���c����Ւ
��<~��ȩ���)ܲ9������nG@�ZN��:��c2�{���S��C<�� �!�_b����W0�[#{rރ����Q�Lx�7�r�6�?��'�t��L�.EU�� )��y��/��=�XJ"5%I]{�.J>����CB��zǢ��|�&�oĬ�J�D�o�ð��
��!�T�3k�fXߤ��pՍM?���-�kz�&92��w�뾂ʄ�1@T�X��w%zեK=�L���,���Io�9��6��zDm|�uz�36��@(���� �0����۪Oo���j����9=�B��[��St�<��H+�􉜮b}�!:�g��-��T�H�v�ov�~g�x�OZ�%��á�����C������}�R��4��Pz>ޥ�G�?�Tl��D,�T�e�R���׊db�/Wx��;�b���4|h���:nO������͵ ��%a(@�� �2�~�A�b��3���ò��z+�A����)�.ئv��j�jcE�u䯬EҀ�Fv��t��g���D���p4ԟmOls`Us�y��xüVQ
i�G�`�V�]N^�E��dK

�����l�C}~h��5��N�W�mB�%g]�� 6����곓^cס ��8�	j�<�UO��)ߚc皏�ɿ��G@i]����)ɲfS��ږ�����/}M��Kz|$8�j��"ȑM
ED<t����+H�lv
��KcE[f�m��C�h�2�I�S�4��|T��I�F4w� )�%e�HV+���z��)��7��lKf/Id��p+�.�}Z��x�kA!�?��<�
+�Qy�tW�M��a�d���u�%1^����(1����K��<{���#�{z���'�=j'CWq�kN�z��;w�?b���]����@NN=:L�/,�mun�j�I}1�;@���{{,���zv�`R����4dm�V�l�<ҍ��辨}4
}��<*T��cj��O��Y��=�2���Y��M��EŹ������l��+������C�Ч�C�[�,b�(�W�D��p��S���X'�n��s�iF��9$���y�F��I	�=W2-I�Z21��r�$Q>�#�큖lY[�lג(7i��e��:]kdf����s�أ���a�Z�7o��S`�ڲy�Q�۞&��C��tH@P#�,٘�ȝ��Cs���6R���8�v&-�ڕ[�:�w��� � G3��>`(fS�@ :�N�V�"�y�%Y�K��(����S�}��Q��V�t�m�z v�5��-Z{N<5s�5OJ7�= E��(���.�>�!�]���v�s ���B��ϸK�l��P���P�O�Beү� !h��r�6�B��ms�@���C�b��{��c��Q������?k�ʅC*#ynt~����&n�{�ѣX�U�}gr�l[Ow�_�
���\'�6tf0<[:v��"1ϟ���p�Ō|(�	�4�W&˺�u$[K_p[����Yr�>�F���������іVz@�W�^�W���UL����`/d�HA
��RM�ӇOw����H�N�r�۲�ѧ�hR<����R���Ru[P��j~����w`a8lQbs��ɢ=�)�8�vmK*BC��#���������U�:��2�q�M�}�ѱ����Q��>�'�`$�-�[��;R%�����R-�Q�r���Q ���E���� hp�T2;��2q�����Ԧi�f��|��j�g� �����F�+^X��f9;]*�V�1��ی'�]�jm%r;�q3Nnv�r0Kе��h��&���GO��H��/��4ҙ�Ÿ�WY���+�D���� ���"{�M�]9�̲l�F��4�3g�(v�����
j.1P�1�h��V��:i�Y��J�x��5��tr��u̘E?���!���`�C��L(��M}��ؤF�W}Kdw��Ǉ���]��y�Ҵ�mj���:��������k�<�F�gF�'	�5�G�&�6���a��a�"m0#�[�ǐ��ЋA�B�����!C);4[V�JsT�<|U}Eg��#K���n�E�?�.�5f��,���-99n���+�i��g��{]��A1Y��1�6�<��䖮�|;�J���yXH0y�j;��>�K�M��qTh���G��07�	5	F+�V��H�.��Fﬓ���#9$:_�$')_� 	4�nv�n�z̸�`��u�������4��gM�zVb��lr�?)��m��v�U��|:���R��"�Soxl)GE���	�~�D#9�h���+�s�^������=��-Iضg������T�nM1�;VN�"���`��P�wTMgJ��B�c��3S����GQ����T�k�*���l�G����� 8*!4E�Z�Gfo��L>ۍ���-����A��}�B.V��߹�F�=X�`|��}��8��`�7���{Xw`'Ba������M~>�d5c(��8��p���������a��1sU��6��V��>Թ8�쨻�Vɫү��!��][o���5zBb.
*}��U�GbK ʮ�*�T��w*�w�_)X���Ӻtc�� 6)��3p�:������cb��_��S`��S��Ë��%�'&!�}���
p"�y[*�\�%��k2����Pڏ/y���e��D+�:�)�'�%m�$`�u4u�����%Ka�N8тRʢ�>��%w���@�epee�C  %����qVt��OȞ4���+��1��ǒt}I�6)+R��R<����\�2N�Re.��A��E���=���5���n��xz�X/-.L2�%�(%V������k�����WHx�NOU���A�.Y�)e��3�wNe����AwD��7?qJn��++��!�X!j��w�ss��@{�v߷�`����t
�"n����5�l���@�I򚍞8������Lpxk�"0\8�i<��H�铜�ۏGr��3���
|��b�%����(X��Ū��^c���[7��T�(gb������4�"حs���gB�]���kqeȄW����N�7�N���{Ӽ��V��y�+vwi!��Y��94>Nn�/���p�.�(Myt+5�U��V�[n��U`ka<�=s���������S��j��bI�od��+��b呱�Q��"yZKR��B��z�2�D�r�Z�9E�J�pW9goܠt����>�QaN��D�oc�Cz�h��0����mqVe!���j��tfv(E6p+ċ�M�����N
L ���Y}X�Zє8���{���y�ݲ�%h�<�aA�,5���u{Ep+gI�w,��#��<�YK���E)	QI'���V��������'� U�?;*�C%�p�0��➡�BeBnAqb�	x)�߷�����A:�����5�SZr�xt4�$NlN�o1���kp;j�$����?V�i������]u��O��?>�G���q���qlf<��$�?U�7�T�_�S{˨^�q0��Q��K�SB&�W���c�僷�|W�%�D$y� �y���iwν;�X��{/��hz]߂9Qg��|�z�^MA��0ʕ�զ����Mʕ��t8)���4����2f��tE�K�4�]�&����FKST���ů��Y�(b8Ӛ9]=#��x����Wo�� 9g"yu�5���2ou���Q_u�kּҫ�M���\��Ko�O�]��ϩEǒ���Ñ�F3�/���b/~+l?��EqgE6�<������v�ɖ��\�/nB'�c���� S���ʡ�Y^!CY��D˪��\�`���W�vH(�B��_`�7� �D�-���PS����[U��U�<�H�:e�Ѿ,T�Z���aX�R�.�2�����oJPK&x���^�CN�J\g��|�8�.��E��h�.�j=G�[�OT�|��3DS�x�gz���5����U��P���e�ckM���'�,������a��f���~�Úk,WAɌp��qR�#|B�L��(�Aִ~����n�<:�u�?v� �y��*��ߪ���}����W�O���	k��bh�.S�[��#d���j�'w��j`�{��<��׭*J:�����H�n�o�j����m���ܬ�ŷ ���{1�ڝ���0
e����ID�@�F9@/U����
��l�l�b@T��d�f��гk.՗�C�}�S�pw"ߟ%N�F~�q7@��j)���D���$��F�;`6�3.Ҫ�q�<h[B��) �"	���9>@k�1ئB����)C�?�7ovD�ѕmb~�y�j�߆�@5\3�nNh� &��7 ړ����d�5����{�yʚx�-N�%Jt�;T�w"�']� T�!��GF�I
Ȏ��C����g�&�0����cM�E-��W
ܙ.��6��M�	�u�
��� |�S��WH����+�
����U�f�A���Pц&��s#��-q��O�Y��,
�^p���!!�t�-+�������D�&
'3���������S��`��gҜl�.�&�$�Q+	��0o%���;ς��{�9	�ף P>P���C���N���p!�{6�q��=��l�����B鼧M��.�,�*1�e��ryA�ף/P�e��M��F�;��-�9���qr?�F08)����n[	I+�Y��m&S����ב:΋�_�g�bMW�G��!R@!��Q��ھ��ra�I�}����x�eM"��=�5��I�=Kx:���Pb��Ӎ8;����>��o�L�݋�6o�r�Q�v����Us�����ykΦ˄�;�%Fl�wƭꨯ�m�V��G�ש�PS�҇�^���#�` '��V'��F{N�DE��	y�9�yAz�B6�X�βH��<Ǿc�9�.ٔ�]Ў���`w�E�������?y������	��4@�ƣ��h���vQ-�!�ۊJ��D�{�G���.��#L��<�k%/��O7AI��\&S8�G`0�w��i���w�q��s
�s�d4�A��]�	$�Tζ�݌@n�.�x���7jPg8u��B�a�s�T��O� ��D�G��&NJ�a\}v����wh?ٷ���Z�����e�O�j�7L�>-�@��t�}OK{;P�Q�>���i��i�,۝x�Tb4	�9<Z�S�(�[�[`�[/[��/�l 1�	.��UCvqg5���^'Y�a��z,nǹ̟��霻#V��	��:h#�H�T�E���	/�������pk⤭-q�0�HN��q�5�f�43tQ�1f�k_�p����젯Yh:6��SIp����5����t1k�{�aIH
6U4���^��K)fYFO��_�M�F�:�o����w���RKC�N���H��H;�h��뤆6���|(�'��͉�u.�}����cȸ��\][��
En�u"뵔=����e	�_ ��*1W,�ք�+�d`����2W��n��];�R��Vy抺�� \vj�w���ɝ�~�:/v�5����q�!gH�_ʙ�yl�_�:�V�s;c���'!f��1�g���~&�@��(;���M%��>�O=ʽwM@~M��)$�r�n9�B�z���L#j9�z�ap̊uį�{�(M���^=�#L���7+�t��"��!�T�_3#��]�O2�܀Z�IT�m%�n�p��zy4�/��Tѻ�
����-y䭉
�0x���g�#�$��ʮDv(���3�"Is����y<�t<��� �!�c���շVQ�1�v�.�LG:�Vbݰ���K���
8 �,�^�e�l�h��x���8��T���sM�.T��h�����c4�[����͇�I�ڵ����btUX�TR����a�eCWxB�Ll��-LB��
e_�飙k�c�&eA u^��s/������g��kw���W���H�����;ӎ`Q�kjfú�M�Z����*j�$~�����TC����H�)��7a����tM5:{X�w��bH8��b��<�۠ŌP������Yl]�ʼr|w3�}�i��[Gz#��]����˜�� �:"�H��*tGH�{�b;�}���!m.���g�W��ti&$�[���odҺ_����V�zǼKM����^�-��&�
C^4��P�����8#Q���LS5����J�A�W���m����6a��η���)�,�08����LoM�:q���D�g�as�V�tIG�Z�>�]]��j؀�`����zr��)��>�ya^���Vd,��L��D5P��ᕃ7+�R��]+
c�[�J���u@�\�PO����v�J��G�8���wm�3]S$2بE�n*����WIC�+���>���ǀ�~	+���&�)��gy1��vfT��"H�(k���0��UY6�R�S���@���9��Z��>��G�aIa�"Q<�?�ʻUs�ɑ�i�9�������j�����}D�at���Kl�u5i��M�{F�u��͇l�5���
P���v�w2�ꄤ��'��ټ������)b�⿋p�[�ڱ
�%��;x-�B������<A�����@�	F�,c,9G�2�č��$���� Q��q��$+�e�Rm,=����22uA�y�Dƥ�C.��(��Ml��!}Y�ۏy*�G�<8D�w	J�V��c� �'�?�)lՑ��j��R�Zu�/γv�~�@e��֙�rK�&�:�#U��l{s�8�0�ĈD+	O*�GJc���-2���|��X�6�!�Bh��Ȧ��!g����Iu�����(�y����4N��>I����\!�D*�}`��������mX���A�]�=�BKj6A)�����[af�~DΧvo�� �Y�Y'w��+6�l�9���eqn�-�Nͬm�㽒�.�JjB��~nId5[9|���~��MM���``�^�5>����y=ʻ/0ޏ�\�U�[	��ݻЖ\�?�e�;�'��.�O g�I�WI팑���=���������}��� �v���d#�3yCI�r�\�%��ȄvWb��>cH���?��4IK��*S��{'#.�L*֡/80ޮ�����qI��Ǩ~��]�r�������BM��զ��D+l2����%<;��"�Mf4�P��/[F��)��%�{`R�{�J�(=}XK��;5l���1vu��np^Gto���XQ�g8���A{��.���\�?Ѐ�2YM͘�ϵ�Eb�����Yy��y6c��:v#�bԴ@Ӆ��#��"p&<��P�S�5�|���h�^�J�R.���16Z�T���
v{���|��鶫䝈B��L"Q���"{��A�������ۦ��	ޟ��Q���B�2��~7`�g�uEi	x�>���\̈�4�qJLBSoR���W����@<~������w?��:�?�m2Bk���2��-������?�}��E��~�eU0�N��T�h)��+���5�G��>�6,+���3=a���,F.k������A^Z5!�4�&�]%_� �3�G-t$�|���U�'\Ӡ���Oz�>�)OO�k��#��=��������u;Cle���/70�o���������Qc�f�{!J�cK�0���V�f�ot�R
q�=�]��/*Q��3f/.��a{�X�P��9��/����wUH�QM~�4S���tֿj_�0�)1�ܤ�-�]�ɞ��(cc�^����P������J�}�V���0�2���p��DV�[�uWVZz��uWO�Q��d�`-掩#�E���I�0FS�c�m�a}0nT��V�*�`�'l;�E������N;w�~�p�rZ�;��d�[;����΀H=e�� W�-g��9ǟ��+�s:6�p�5����rN�0+v���(4V8j�8��<�A?�zT���D�:�p�Q�g`a1���q��[?��씸����E��j��~f��:�KM�QC1��p2���{Z��.��͍s��Hg��sr�_���z����A��4L�z5w��`Aٸp�`c'i���6� �� %�������Hq_�2ۿ���h>�n���/B���تD+V��0����.��~70�=@����ʖ�d�{KN�����3������|w���)�TMVl�6��熖�Λ�j˪|˵L���v?��W��@�+(=hL5�(�]|�>��E�|��}��VO���ӥl��Xۨ;�W{��]�}��)�H�=䔆ۥ�C�?͵����^�6���{^tc���/��ѥ���e�q�$����q��Q���e��?��� �j9R�`����)j�Z�J�$��?�[l��0o����+k`�� ҷJZD�=��� ~9efd�k�I����.`�LЮr�m�]���&�q�4	�9o&D�Iܧ�сۭ�74j�{����88/�,�@�|N��#��w�O�;���(h��E˘[��1z�s�5NkW+".�,�Қ,c%�2�ھ��*����i�K�������
_�1`��!�GC�݀��u%��3$�=�J�8g�x7�ҏ��B�Z���#~E؎(sj�35�&[9�o@����gC�+`�F�u�'��M��^�S�_t���c��h�~�'k��C?�BW=J4n�ah�y�8���,�^#{��j,2��[��ٗ�+���>=JY����&��R�k���%!�/�:�'�
��n�B��c�74T&T�*�5D������]��wQ����_G�J�qe�+������Al,��[G�K����㋁�"�"pp� a�Lj��Bd�{]v^^ �i*�H�cn���`�ǚ����m�=F���8�gEQ��;%.7�T�Ș[q�f���6�9��.�%/��(�ǒ���-�y�a�ꍰÊ%ծ��ZL��×֝Wfm�>MJz�8��h@㐕�3d��O+�JO�
w|�NЦ,�T�g?$��2R��.ck�����Y(�u0ꆓ"Y�F���U�%�8wf���A���i��6�/	�����rC����_X��T�IRH�+�{�K?~]G��qMǨm��~5_M_�[X
��k��3ܘ�6%�,��S���9���7*[�M&�����:��Q��BP�ξ;~�K���Ye���S���^☽���J<��]�L���0A��0��[� n3���%��ݔϦ�29��B����R��_: ��f���,�_�Y.-�����ֵ��h<4^e��X����A/}+!��щ�B�Q�;E�����O�/�yZ�os_�FΙ�7Ѣ&��_<^�:���0�y0 .mF���TI)�����R��{CwI�Pdҿ����'��\h���}�Ȉ-?{�u}�X��I?��Y�g�)jػ�YW�E��u��-��CĻ���|݆�8Rc�<���۹��^f�Ѹ3�1�+�c���Z�N��HBg�:�u�0|5dw�
$�6m<n,)ta~'�薨��5�q�G>z�k�����'��V$U��Ŗ$'ä�R0���l~X?*�ʵACk?'.�t�)r?�_y9���5е2_}n�{gA~�S��cvOp�0��ȇ���U"��R��| /)�Y��76s,�R�Ł�+Ug�_u6���!���5zȿn�1Kb5�r7A-�{Na;�tlj�d#�"��r�ꋢBOa�0T2B,ᒆP�}ʏ���:�}O��'���>�`�NȫT������u|EP��pQW�Ү���<�z�P���w|���~4P%-|i��i�!m&������t(0�6q)~��7�mD�2傶�t�d;r7�p��>�Ҟ�ֳ���+c;�襐�p�����߭�[��˕�M�\.R���}L\�A5 ,�v�[50]�k��k�2��>w"�f�M�o#i�.��Xp|�FaB)ĝr*��}�C��&\�AMW]�m3\�8�5�]�v��m�v���F"E����?P2֨��mcRe}�R$I��>�I������t�㍦�N�_C� �`�
Q8�C�S _�K=�h|i+��C�@��z�0Qu��_�0��WU�R��bVv�0��Z`Q�[�?�����T���W22�v*����R�V�La?�X�P���=u?X��'s�l�	�D�s`B��N(p�.��Y>�O�qoQ��2��"��Q�
����1(v��"?׎����K�~��Z˔E�I������/=�@�"T[�3'#�rФl���ϟ\�� ��Q^�Ii��%G�>I�J�XU�&D���')�7�%R�Qy�k��5�σI@����8�}n$�Y��N���*-'0{~c<��~I�{��NTџ�u��NSk� L{�!�eL�5����������()]T奿d"x+�������8�#�K�0*�4d۽��"�  �D
~S���l1�Ɲ���.��+� 2�Z[]o\�[�����"�$���d-7%3���S�7�*=g����j�Z�D���D��u	�7 S����M�P�w�!���1��N&jpǼԆ}@�F�ƫ�<e,_�ӪLoR�x�C3QڿU��rs�?�Zੌ���Y[ǩLڀ�h"��/�&�]"M��FA��y��	BӲe�z���0\�g�Z�/[�y���RUI���X�3�a��@Z/0yG�ˢ�=*��8ۉ�U"��o��T�+Kj0�����G����#�lH ǝuB�	'}l�h��}�ng�aN`)��"�$�����85E�|�J�9Z�M�����ѫ�%��)�����������QS=�JzDh~��H��(�-^t�4+�A�b�y&Y�wTjrL�X����^�?��,"�&�$����#k\�Tc�ht/k��"I��, כ��j[r�=��pbױ7� Y�KF�Y�lJ*k6����"9�	�R7�m�]�+4�f�t�6r��,�lBؚ�P׭c����R�X?�+[�F�TKng�"�\V�Tq�����넟Y��x�&<n;:/QN�벪̓2WB����hT/�é%�E-��ĳ��=�ĺ�j~z�b{�UD�~�iL�rU��#�ǖ��J�ݔ~�R�8GONd���J�����IW�f���iP��ėOdI`����>e�V�+�\_��Pm��b5�Vŕ���:�6{�>�V�hp�i���`O���l��UNoRP-_Pt�f�����sյ�"|S����B����-S�b��g� �o^|i]k�(��T� �6�������d�ۖ����&WDh�P�[#���Θ�TeQh{�	�]6�on��K�T(��G��  .g��}G�������#8x�h���vn&l�&6n�]ݩ~������!3�u|K���fȟ��Ss1;����m�����)h�˞X�#Cw�$_������@�=8,�st��U�ӴΤ��y���z'g�Y�`n1E���e�4������y`���L}`���q:��Q��s��N��i G����y9�T2T���!���H5B?���,��x��R��������@��p@M��ē�c����4��46��-��~���}:[�A�Pt/�_���Ut��pB(��[o��"�!n�߶�#�R[�M�u5�Z�P�g���#������Q8[s%�;l�����) ���д�cA�oD+VP�6<�߅�(�DҕbF}�s#�����|<���9ל�ڶ?�>�	-���T�#�di����F��c���&#�"Ņ����4౔���i��3����j� �4�&��4I���ez6_�a��M��m6�녧����FD�yp�i�py��o|Ek�i"�w����K�L�W�|�`�ŇB��HO:Ϥ�Ӛ`��e���KF�T��.�G�R��ApI��N�V�����G.���;��@�`�HL��}�N ���3�/��2uҕ�[�_PE>��ΡbԻ�?\xi7�A���"�gq_e��1��N!4��Iw��c��Oi8��xW��(��	Xkv��b�AыtG�8���bcI)vь��^� �KF�4�t)8���[�"7�^!�����x� 4�6q�h�
2���޸��;�X>�\#���w+!��&)1�n��~�>��+�g�
�/R�X�}�,��n� �Lō�����#��{�O��}�%i6apt6a���dKВ�����
Elɑ��F�_a)���za_�u�5cg!�x:^��_sĶ�@b��#�g�y��g�H����}&�WH��H���9ӳ�����j��+���\g�ђt1�6�5��;�(=׀�Yݨ��`MT��a�I�L�*������a,��q3I�	�6�~4���-v˔A��t^������-�sN87إL ���������b�F�A�m��b��������q��.}���M8��i�|�L�º���ւG'��9ƹ��l�&~x��[�ɷl/QK���v�ȩ@�[���&x��
�ݚ����t,�i�o$�ԃ�@�ɔ���.rW��&v3
��':���i�)KE.�D"���������Xl� ̋k���- s�/ �e��a�KtЄB0HS�1 �w�t! IBL5oS��kr��~H���F̜hf�Z?��b�6�EQ\r��}Ѕr� �K#�o����ҾZ���b#��x��s*�x%�[_�oM=7���ȯ�uU&�����GO��KYLf �ԢYA
��g���R�5&و�~��*���f�ÛF�\9 ���֕f��G��������ɗF��'HR�l7�V{��)Q�q'���� �#�UC�M�r_�MT�����C�A�1���B�Oc��hr��MP���� K�1@�~���vMQ7���`�9�L�2��m0F������ҳ���w�[���f��,
���M%���͞���cri4S�t��Ny�!bܿ	G��C~67��e�:h�]{�Y��T��^��|�b�Ӌy}κD��Ze�9�>�r~��E�r�-D��Pe�E�|�<��60~�9\�;�U<%�eL?������K3`zy���3��ĸ�CB���7�`����o�������g}������XLt�C�N����SyW�6��\aH��g`b�+�ѕ�M��r���5������2�$�P�O�������l!�i��x@��uK�\-;�O�l��y��Z��샕��!�7�m_k����I�.�d���ȧ&:�����%�Q�D����}f�i����i�5��ᙥ^��d��*hB����h�y�[ ��ͬ�~��~����~�U
�/��[�	}u� ԍ�;#������\)z�x������?x�o�4��<�d��Ʈ 0������5�L�dj��[�q�\Y����L�0J���ܲ7P�i�Q����o!f;�����5�@�[]Q�9Y�ے�M�=�X��݉
�B[��yx��Ua�Ko�k��_��*Λ+	�h�V3J��x.�gvo?o-�`d{ɛ?��ͷcD_n��
9�{��
y1{��-R�^��+|-�n@0e������iv���e��� �!�(Ӿ5/>P��l�f�OV�H�B)Q��
�?��֜��5A�k��4���ɝ�%Ex%N1A���	h2jO��0n3X7��X)�ۑ���;��0�(9�7�M:>1P��%5f�P�T�2��t��/�Ԝ��j�yaO���0_�0��S������l�� �Wo��G�͜����HI��H'��{���@���h����(�;�s�3��n3�K_sd$����%y�Kh1�Zn�]s���*Q���r�<��`c��}n�b����q�ML)k�D:/�kp��u�覠�U������4H� <�%����~"n:�ꑫ��ͻ�������j��Y�Ua�]�y
 �w_.x�D���!����m�F��[����lnvǐ�@i���!N��OR��:0VQ���1��Ŗ��7�=朗|�O�����w�����<`���q>�搶���uf����bx�L��j�e���A���Q;�Y�����J�JH���$��@	g]����^��d��.����]�����o�T�iL*�8S&t+���!����;db�t�pC�lyvi��r�_�s4��E�@>_�`���T��|����{N2�ޙ�4�)cR�?�T��μdL�89n�f��+��}�v�b�0��v�	qx]f������b+��L��o�����K��#��
<؄H�7U}��j�B�2�ml���)K:u�h�p�SȪ�~��ڦ y�2�;�H[��NL�����@�5�Z�(��M��;��K���<��U����	 �Z�5!]?�6�"۠���s�K<�����E���������7j&�m�
���O��_�W�W����g�!t����VMpR��A����ܶ��� ��X��kXHb:+���H��	C�_����X�&kڃF�Z6࢓�ʑ:��&QW�瀣v�zh�,��7�rT�<�f��PJ�~N/��^k>� �س$�W4u��������f��@W��6[
y��+)ob�ajc+GHU�p��c�e�[��Yd�}��X<��`H/Y�z	<�e��ڄ���Emd���;;���e�@��ճ��N��'���ⶲ�tD�������8�";���Ka*���0���n$�a2�ZR�nc�6c)��7����$��@F�Any�<Q��W|>� ��_��Ҹz2�h��)���Z}��uZ�"w�׍�=U�������p����p�HDo�*�����p7��������W�&����w'��9�p�qOt����4`%`lt���_=�����aD������>���ٹ�O�a�� f` ���~Yp��z(X0�]c�4?�GA@�;߬�M3��P"R�y.�_�����6}t����p�
��lx`���՘"��D_N��/�X�<�����j��c� $�%���+:E�#�����qS��dہ��{�O�~��l ��G��Ѧ�V4�餴`�q1�97��&��H;��՝G2$�u�]�-���Mp �D������^���%^�e��l����Ik���}X'�L%�e��-%#;����v����T�<*��~��fvǓ�w�׼�~S_a��'��_ݵ�|l�S�;~�X�' �,٩���V�Q��׌_@K ��P/�{d+}q���#��m?߉�BrNK����qJ���Y���r�����)�Fy>䙽4��V���4/	��4\��v�D��v�;�c��9D�<�`��\z���z<�jRΐ�����
r���;�{�x��)�na'��R�RD)�{Inh�
H����*�?� �7��Ք&Ap���"��خ��ژ�Q�ߗ�u��|��Y��腯��P��R?�s���xb��h*1�|��OT9m�Pv��lLL��z��ìݖwF���ӟ@����9oZ�b9E$EVs��(8!>$�:ڒ��D�{�9��$G�²O�NlY�jL��������3���dnV�HD)u�ѫ���f����O5����D��-��LpEs��J��Z�u�Dʣ��;���;x�����G�X����vF4Ƙ�~����K�[�iF��skmt�s	���������� �0�X�7,Pa^^3Zƕ"^�e�G��r\�
%B����2cm8�-r�fͿB��$�OQ\3�sPd�C6��K�"$>��+?�x�=.�T���DJyg�h
�f&�	8P2,�u���!� L�plS���ƚG;3�Y0��`9M����̺+���A�
#���>}0H��S>:�P�x�6k4_CJ�*U�:�9XI)��nF��q�hX[q*�s~Zu{S("��OՑ7����6��b��� /f�yT�>�%�	V�ҥ���n��2("���\H����o�([&��R�º!h�̙�
Gx�=�����ȍ�9�:��c�:��Xa�wkñ02�"0~����I�U
�dW�q��tA���E�	���S#��X�/Be١ ��|�󁴗��IV��{��"�����s�L�=�V%?����:�Ǝ@��D�S0T�A:S��	���1Mׁ�DF�ē�^q�X�����3�J�(� �~���8΃�[��7)B3� l5�v��"�ԽG�G�vG%pX �[�y��{"���T�;k[�&���0, �N����I^i��\�?�A��w�R��pb�"F�k�<>5�{1�G:��ƓHs]+zpv-N�><w���V�2 	�B�dWz��/��� U�XW�M`e�ʕ���G`��'R�=~%9o���S?���?T���맋J>:�Cդ��#��]�ps�@N�	r*=�q�Z�
 %���2���~�0� �����[��#����2R��L���]�8*PRT��F����^DzT�^� W�1Ͻ쓍O�Ӗ���R��zI��d]�2��/��r�D�i!���5�1T����.0T)���rR�Jd��Q�_g�RnxDl�:��_�M"��P]@m�3<ͼ��P���t��a�m�f�����ػ�fo{G�������x!�_��E�xi�)���������ñ@�������ｙ����Ė�a�C�]Yt�d>�����yYU^�H�:��қ�#�'���6��ŉ��m�\D#���$���R�� v�x�K ��;TU��Þ��� �Wn>��4�w�)}P���z�C�[-�W��zP�.;����8 ���A��4���ɞ-���'}E9���(k�	 L�/�y������X�M�ν�9Y[���3�?<zO������vt�sϠn����&��U��w;Vp���]�	��)a&;���8#P������x~,���L:.?E�͛�3���DFR�8q=P`?�z,ߗ��*����sŮ�|6�Pٹ��;��Қ��?+��gn2���d��S֓%,�^�Rk�}_^�$��8<�����7�%�r}��fx�,_�.$H3(�X����Pzq5��	����Wxm��<�.����h�U�J�N�-��(QY-��K��9Y�h0�)�#�۩�9��|I��O�M?v�� (���t���zX��lY��X��3�{p-,4���`�����<�i�WZ��Y'��밸���>��f�?-��Ȓ	���gS~��H�#Ǉ�j��*�
��I�d%ﺊ��v�^Z��t�Bqg�F���*�m3|i5!�~��?�JY�H�,�b����c*�����ÔW��f6h��\q�SP��Z�0S�.�#tQ����u2?Fg��]T������E�3��&1���;�B��Y�p��Jrrίx���B�e�-s >@�ݝI�&�)>D���1n�.��'�)���0M)���?�2f��d�01V�J��'��WĖ��ő�4����BQƿ�=W��ew+n�Mv�ZkF	��ҧ�#�q>߇�̑�i�x���-��6�M��	Z�C6�uq̆CR�x
r��˸�@Is���[��ZI_��������|X��3*$�f3ݴYzP����?��iPB���t�ܦ��0t��	$C�an,4�m���A_�n<��t��0�X�6|:1��O�W�t7:�		�����*5�jj��C�B�ZW�'w�3܀©.ZE�&��kYUf�����劢��%�O��{��L����鴝h�ugU�_�f$s�;-��U��)V��C�5_�Ϋ�Zzi�3��1p�G�d�9a�[,��R�OF��7HH�?��M�"ݑ��T��aqLV� ��!��KwuY'9"(Ӑv��1�hH�j��5v0��s�/�Ѩ��X���4
d~ܡ��,0`�m��PFT� �H>bwJ4B10?�"�9�= 5K
5�g˲B���jJ5T�ƫ�La���G`6����w�|����T�ps7�n$��p��똧��Ҕ�'�� ��ܬ��f�����gTc{�I��qa�Mi��ٸ�DM|�Wt�/�t�L��ʧ7���C�k,
���a��2����c��v�r{O�~<)���"��DXYW��nn������ ��S,������+)A�0lK�O��{H:Q�֠v��hJi����4^s0��A��S&Q����c� a��䔲X�x�}����4ZK��D�/�J�G��b���Tq��li����"},��i�R�X��������3C���ol�c��4�������#%����`&�p��-潧�AZoGXgyw�R(��p��!�����	����״�z�Z-�B�8I��t�1�D�_QSVs&v!z_ڌt�lM׳�{M:�S��T:�=�9=(�l�|=�0_n~U��JQ�����?d17�2���Pkeg.k-�,��fGYδtIqb4d'�y�$�@����AXq<m�%3XB۟;���"�3��
��c��d�zd*�ӴH6���'c�35oc����	(:[5̿E��7ܭ)�j��Xn��Z\0�Y�x��&�������A�e���a����)K+�i��5��gްT��d�mSc��\�+ik�dȱ}p~ئ�z�齃� ��/����bxZ��H߭�[?,3�  w� X�`�s�u�$��?�99ʩ�G�~n"�t�[�,�b�#�F\��l��Fi���(�k���mF��P
���^S,6���⸗�t��%�Zϲ��a?�傠B5QL�[�h��T��,"�G£��凾�b�A~w��0O� Ŗ��zs�K�P$-��2(릹	�yk��E�𻉷]Bz��y��S@dŒ\��Ŗ�@��.��Ub�@����ҨYu��&���KILrѴ��,�L]��Q)8h�QK<�ś�4ɝЙ��s�^�:8�:�a�+�]2�RY�g@�'��h�lg��?A�G����m�_	��{I��^x���?Z�+���$Ֆ~�W%#�u�J!c��d�*h��]��]l�lXƏ��S�����7���T��u��VVN/�x��D�]�ɠ�M��K7����qX���@�0���{>�&��ɞu���rXʀ�Ue���؛��"���t���J|�޹�#W�&M�y�*�T wQЁ�`��=V�rxZ����%p�d�9;C�
|�dR1�Rs��f�4�S�� �4�_Y�'"��G�3����ؼ���>0��\�$(۴+v�l�,�0�2�� W`8���)�F_����5�	$���;��i<��S��Ϥ15?��B�o#�U���;-@�<o�m���}��;iVJ0꠵݌�|��Q��y@U�������64_K�P�a�ܩ��ET�M���|�H�iIr��՜�* �+��3F2�M�c	�RQ�Č��cv%k��%���h(VD(ه�ϲ�yft�K�����u��OE�kC��׎y,��#��3! 򉐫�qC���d*�?��*)��e�goսw���(ɾ���֍	g�i��01O��m+�7��x�L��ҐS��x�O2J���7���wq���#�G|�e�-6:�DaT�[nx�	���`8�͍���`J����=M��7�yDLY?���{C�
�o�"r#�z�a�Q�fYcx��~�U��)ꢵ��z��S�/�<@ҹ��u�y����<)uuBvx:�|?"��Z�y�b�ϊ��H��h֫/���اC�3��3��������ؖ0(�����%�!ݣ?����f����Ov~#�L���L��S����Uт�)@	��QXh��'㋕'�C�@>rhE�g���ƸA���^&"UI#©(oಟ*C��.usfH��=����(���}�6����o���kʬ�C��>�,?@��#$�'c��E�7��7,�c@{td*�{2�h#�tL9I���$���/]܆`��ٱ���_��0�}�D��Ԏ�*!��ȁ���w|�x� �������'�7Bp�Hk@�p02^㗫�?�R5)����h�Xd�3*��V�k<O����<���Q��#�USΊ6�`y��%%�4����_l|K���_�5 �s���ei"�R;�`>'}�:�tUiv��F^��V��&ĺ��=��̖�7%� V
�S�D��Dr���Iѿ�Hes���[�Ё�����A{����/�$|eǓ'Y�%��zS�;�����A1S%��mĨ�0- ��-,�f��'�,�X>\ϋ�����[PK!��5H��X@/��8$�����5�U���PU��/gp�pQ�=@��X�%�Ej�.,rKJs0��j\\oM&AfN8��6�"l��5Vٱ�5Eµ��c�uQ#��{�� �M���l(��2��e�q��H��4<�T���J��<�	��1���|��&�ɼo�{@"�a����ͤ��������S{��6YoD#EIO��ň[�U�A�w�w9:l����9��E��@��G}V�폙�n���3���If"TT!L���P�	����}��g���=�G�n��7�`�J ۉ~M"�d�a����0�|Y֭��Χ*$��H�j�k�.tL�#�x7R���V(�X���3��]*��݄e�Oc�5�5@����#� !?~+q0�a�;�x�3C�!&V3�J�e��]�i�BMߚ��6�dqE�{�f1?��z��,����f*���I=X�0�BI]��(C���է-�ꠣ������ԟ�z��t�ڹ��ѷ;څ������W�$�rWH'��"6'�[�'rU������j�uD������Cƈ=G����U5)�K��X2�S�eކE�&��r`��VCx��t@�E�%{��0`�/�9�c��"�؃����Vo���i�0����Q���<�-�=�YKz7؞P��&M��:�PjG���j(�����y�����lr�_�J�<���T,��b��(!<�Ǎ,א��rC,��q d���Φ��" �b��Z�+GSd!�wx1HW�j7�D���d�����t�A�����b�n;M.Cq��:={J�_�qA�p����=�]Tz7 "듕|���Rm|BDC��Ut+ ��#�se�?���v��#��G���e�p��8５XN�wd�)Q|��C�}��#�Q��p���ڗ�3����ǁ��W$�ëM��, ؼ�t,.4��w��yq��U�����jr�AC�7(���{�N�;q�MF������;�P��M�#�{I��$������^��h���� b�����|��画)z��#��=�.{�S���J�����w%6�{d�rq�oz���q���?�e��Jr.��`���d����;�/+QX�
RV_��5��'�jR&���~��k!0W�1����-�ztM�N��(I��/#�܃����Ά9��@�H�HK�l���TSu�i� �f��G��Q�c�*�Z6�_-�o��QJ��k��f|Pr��{|��S:��t��UF��
�+�����c�*�����ۻ`�l׃��R�E5�������}�2�!a!~).s�U�����C4U�b,m��D��l$�]���׀S���tk��)�\�jPe��=��֘e����L�I2��0�j�%ӷR��x�Ry\Pe3FXh,Y��T�G)	N�#m����-���Ds}����'���"�(>��P-W�#>q�0����FC�[�w�e#�3c���*w���y���o�/烦Z
EM����3�4������l���N�:f�px�q�OK�qv�<$���H�qR�ۙGqTػ3��ku��<�^��G��{S��悍�Ya����]Ȥ�\��~۝��3�t-�+���F�'�1���+"�LM�lG�f����)vT��Z;X�ט��@	 (
�ڮ�͘ �Ml2�*���!���i�������
j���z(�����#�l�U4c��j���ǆ?�ۗq���K�6�������l��P�Q�����V��_̕MOaW��+'̅�<��6¸9�V�
��ud�n��.i@�<��tmgx��GH�2���v�K�3��4�H��x���<V"-��c�a)|O���|��a����6$)��S#��5Y�j�{�/��3���Xa:"<��`�-��k;S,�s��/�#O�L��Jh����f͠��^��Ha�~��{|������B�(S��pBhC��\�V�K�J��]J[dף_:t|�o�NJ��ٔRS��\�g��o��K*! �ly��vH��3���tr��4��V[T%Xf���r]e5t��uq����2Tצ�8T�Z���x�9����ig��g�h��
��<C�P+3�`�c���e������*�QF�,�t��`k /�{/���?Κ�W���7��4TB��W D9�r����.Prh�j}�M���9�#��ȸ�f'1ݖ��� q�b+r���(��J|�$)��},r*���Ԝ/XH�n�a].U�F�i���
�{ @*dU����o���w*�Gl5�}dmim���j{U��.NT��$������s6ؙ��$����q%���[�wK~���G�����g��:�� eA���-^O�A;u����9^�I�m�r�����M�$����&��&C.��p�v.�:�$�]���҈a�P>K���^��<t�g�^��{�L�HuP(I�
o��y�:@�4�gFa��^)7^�ţ��R��t�u�w��Ch.Q:���I�e�0t+�(�b
� �KR���{��� N���4~c�v�Z)n��x��緷��]��Q�>�*�B͙������j�F�1�������{_�"�$�j�g�[�r�: 윗���20��)�qx�ǵ �~���aX��*N=_�fo61��\$�?��W{�E,ލe:��V��X�a"�a�]to�{�+1��G��j��R�V=_��V��%�9i9�?�Bc۴��c��m�mo���J��KW2��+2DD�F�3a���ʙT�����!"�U�#���{�<Z���:��ӥ��Q�/
$M(�c�T	�C�l7qQ�[���H�����*������L�	z���oV�2Ha�L��e�nn�TcQ��=��~|OӸ~sY�^����M�a�RcT���"c}����ƀ]�4#\��fܶ�AI&b����O��g��׌���.D�e)�%兝�+�f�����A�vEd&�#�����>��l�d�Qf_���8�xӪ`�p5K�.�Ɯo)�h�Ǆ��?�p��p�5��vE�=ǀ5�M%S�V���1a����M�����
Q����ڱ�=��-�b$�
�4, �d���F�N�k�j_�1��ixڈX��0�l�'H5�������i�r��!�r�$���M(��!�>�W��[tX>��c	4iE>��ͅ��@j*���ʦ3�T��� ��0�-���fd��� >#"�R��7����հ/2F�Ԍ���n�_���H�A�*��$U@\Ͷ���!I,'�Q�SF��5Z86K&fwBc�f��A�MBڃ��%	Qj�mg5�\���PN�Dct�ڇU{K�4	A?���I����ݫXY�SU��p�μ<���DR�"��e�s���J��WGR�|V��k� �\����C���X�@UV�%|�Ƶ�JJ���M�7ъ��(��v��̮��5��e���!�1�p��܅��"�-�K�J�V#�I��ƹ�/B�i�4���)+�&{�ͻ���Lt��>\���h��gLEL�k����C��p�D�<[J����?�1�չ��c>��cy��Ɣ�'�#%!��<�,AiMa�]>H&�p��K��;���g�;�rUl��y��+��=�`���U
�/�"��r���7yn;㻟�M8�c�*�%�3� ��r>Ҵ=��W8��Vy���[��-xu|8� F�4́�>�V#�hN�o�(�Lk;�Ŵ{a��\џ��<���\.D�m��������0�Ր7�o�G9����J��
���Q�[���u��`g�\d7K��wuqn�3�w���#��/|����86�������x=��De�D����_�9d�ώ�	Pu��� f2Ek�,֎c�m���"M�@}!�fTi���3zX`��I�Z�r@T�H���y&lh��{��P��І��`����ܨ��$N x9zCv�����a�?WªZ���u[Yt�� :~�b�@��h��r��p&tɗ3�{ޚ`)���n00��7��5,
,���	.�;7�ƽG�����E��*�B21H���=k��>II�I/t��O�y ^��^j�d��u���Z�u��9bt�m.����L�K���Mm4����!f ���~���B�s�4�l�n�D%h��bj��.i萬��
۴)���fz�E�Df�`44�s�B�Y�*�k���Q�G�5M{Rd59Ko,���].G��3+b��Փڱ3����'$���a)�d?��٢1�Q�k��1���Lo�0܏Sf�����A;���GIu�n���y�E�L�P'�h���/[V/�\��������Hw�����4�FZF_[J�P��0 Q�w�T�<�N�ƵŤ��H�9�%e��8t�u׸�q\=W)NYO�	�;���-J ���R��K�&}V�_�%2��b���� ����Ho�p�ϔ'��<��Z>�=r�7M��q���Ţ��.��������3����kƈ����Xm@Y��nU�ۋK&Ea6S>|AZ���LG�n�m� �v��T��7�m"�8���%tu:������������9k`�c3����AzA��k���͎75U���.8�>9:IkF�r�V
֙@hvd��h�|���{i8g/H�2� Ӏ��e\�'�#��M(����ʁݜ�,�����r�P���
M(7�;�K��8
e�2�&�hW��s5�㓭���<询�t綶_n�$��U�J�mf*��D�����ԍ��|[\�ʘ^������t�!#�֫`���F�e�����!
�w"nS$�u�nQUQ�ew�]�vN�S_�5J�t�6)7���	rX��l�Yհ/A���յ���~7�M�{eg�������M�u[6���:8�Y@��.HJ�ә/��a��^ZfI��gwkR����+��H��|n0�g�^Du�~�܃��E�9�٘�N{�d���EÙ�����>�1�CV_̰�`�_������)� �0t�G�_e��^�;^PH���П�$�aI��7�8ӲQd�p#̝Ր��Kն.�v���(�UNw��Qh�K�gc`�|��9���N�ك3���mO�p��3���Cя���M��D�e�>�Ȧ��
B�����R�}V�P�x�!Ԝ��[z3R���}O��I��L�>?~}B�S���%N��p�s�y;���7��[c��i�M�/�64\����~+����ϊ�6/7B��ST0��2ein43�In{���Ǩ��!��)��� �=�����1�=��X����]q�D�&��y�̽)�G�_�G>��	�e�E�����������D�_����e���:� ���7.w����{_���#̸^ղ���q���	U��z���J�d�8-�.�jG��'��-��ǉ�f�j|�;��.񷬝xpg¥J��(����������@�U���޻�6���=�qp�æ�Q��{�|z��,<�	N,�VA]���i��zs��4�qSK�)yQS�VF��.$�����L[kRv�
�O�7"^��s������'] ��tr ��O�zaU�x�2ɥ���Q����&3��m
�4M(�a�N�""�xv�IU�z���)`;��*1'�����-��$��E�yb^�W*!��.����7�����W���0���ӇU���U})���]P�x�$��������.����bp�Iu�JI��c�s5}wP��=��X���^�W�s&�䊵�\��0x�o2��g��b� UZ�/�&_"r��tI�69uˮ��МG������B$�d;���;,8�V�;��t�.���[r'jB�ŀ^��fR^8~J�=�Q>�~�LC�:�7����~(�8[K�[b/�5�uo٭��g8�T���׺'�e܈�LB*O|
��0���g5�
�o�;�Zn�^軆�=ԙ�q�^mZ�������AT��GL+;��-/�-�, $�T��l�0��s�>Y���;P
Q/:�@ �*f�u&�Io�+���\H���Q~ش��wKx[19�.����!���<��쒩���)2x��U��`:D��,��E���S:�Z���L�GB����l~��t��8Zdjj3��MI
+\�S�;�	�����Kny@�J��'�2`�q�3sQm�0$���)��9��UL�N����IW��tHm���âƣNp�V#G�&2����$�vVʶ'�������֣:O~�b��é�fAk��tR�D�5�͚��p�� m�f]r�%M�*��>�b�
����������ME���|�e׹�g�+�5�|�>������W�~����s�-�m���E�gz��%����L��.%��5��,�$W͹[���PMԶ����Rc���B c���9F�A������Wk�����LE!ԅ��R��)��i�d~.򺋢�����W�$��Jo�F��i��7��K��d��_vi��ďJ	�x+����/æ;��mf����?Y�+s�.*�$Q
�I�v:�B�!v5xD?8�O�g�x|'���AJ蟇�%��U�=�ڴũ����bm@pz�2�n%J�!�,v*|��Yv�5�ͤԗ��A��4%���@ք�Lj�Ņ�y�~%���+UxsŭL.l��*/��/��������p8/�Ic�d(H�f[?��j���R�"�7|�s��ȗݢ��<��0L$|Ĩ����7�~�ϝdܦO7s�|�����c^�7B��F�{�^)���Ww&!IҠ0U��J;���"k(2�}����x.u,(�/�.ЍBf�IƑ�%P[�Wy�����|��yBHG��<~���(�
 邵���W�	��@�b�f��4����#�Om�.�9��ȵ�>��D��Cw�y��rp��C��ظ%޽�lE�ݵ��<�3��"q��iw����#�����X��s�c�{���"]yTTן���Y9�����S	��H������:�5H-Z��`��>�cl�t�C.�Vs倧x����?8�%��G6[6[^�P�}A�m��׀ؘK�:A~�}M��U��f�K�S��
`���=��J�ՃJ<�<t�p�_J��6v&N"pK�H]��+ϛ�xp��9	x>x�ij���*j�0�-�1�4��\��GԘr��B�#�`���ߺsH�5�K�$�Ơ�D��N����QaLR�Ձ!]�_�d!�<B��"m�_.���i��9%�1B�4\%�ie2��q�g�[5K���qbi�jh����k��h.yXU��=�z�� �$���$���.K��LN�bRZ�M���T�@���ق��:	9Q=��`o�T�~lX�"�5���	jD��/R=���Ld��S���5�t`G�_랏qѿh��w��+�t��/�S2e|�3��]$}EE���t{�>�=��.�	\�[��{dY�Ip��_~\���gW	������.�J~��,����M�����9@e��!�`*�Do$�%Ř���[��X�e���ˋAS�	���W����5)��YkǶ������n�DF�`�]\���V-�H�D��e}@��dh1��:? ������ѐU,漹���J�,ٰ#J섣���n�0ɟH{e�]��f�ψ���ӆ66g[��rǜ�d�4F�pu;���[�[��į (�R�1��o��ؿ�ds�^P� �g<��a>���3S����_y8��-:p��N�t�M�%᠎-1���H@��{�҂;Nl�@ R�	-N\���{��X�7���W�ta�8�Z׮\�[����L���+)
���0��2v=�X
?!�w���A�pO�g�ʨ���R���7���ۚ1��y�ف��M��P��mi�288���:�������D�0��/� ��8��1YxLGhP:K3އGh��oB��ol?�j��F!�-qÁ3ig�#&3�S-`ѵ�妬��S�Xb�^9Y�
_��A��u�+�!c�:KM�<�q�<���>�_�F����YL��f�1�	��#V�r�N�d��b �!��h������}!>$#���ʐ�ɴ�7مu�f�1/�����]�qЙ�n���awңߨA�8ז1"
���q�y�.m�將9SFp���:���b�2}��E'�k�ltu��f�/]����l؛5N���Z'���b�&����J���׾�A^J/g�-4���c�q0f���Rדx��{�s!���:�t[4q٧���H�s�9}�C&�k����r�� JC����9JzG��dY;�X	^��9�x�-��ٰ@�HM��W�01��fu6 ʮ�G��3��aia���](�9�3�$�PJ�߱c�����AF����=��LY>����yqOΒ�=�.��[�a�ɀz[)�{no��Q�����>+@���1r"�!<v��2�s@V�QET�^8Yn���T%��� FP�Z�$)x�����F^Sj.�������(D��  ��d�b��	>���[�:�dܖQGF�rL~���N�(Z�����'Ut�c��7&�9gǴ����'�j��K_�,��߮����4kjכ������V��#c ���	���"��K����)¾/v���	�s�B���s�ɮI�/8��5nu�1>.w��
J�vv������Zt����4¼A�"��c�О����S ��:����ws�6�����b
�t}��5i{Ӿ��d���}X�[�T���(��V(��o� ��B����AŬ�zE-'	"�m�F�yۋO��w�,}�J��?nO�D�nh>Y&MbQTΆ�ak�#�R��L Ƥ���@7��27´n�k_��㉏�D:���޻���}c��tP�+�w$�p3�H�`�5��F���q�$�����(/�N��Z�,d�}Ϟ�}qO�Њ㼡�odۗG
J�{���i�ɿ�uē֓
=������5�/�E k;�s�'�z��p��S<�� � �&|��e�包Y뫂�B�:J�a���E*�k����t���k�\���K)+֓��A|��w'ۙ[?�c�.���`�"x'�}Bk�v��V�Vv�t�D�Mm3�����H�'�?u4x:�G�f��k��Ŷ2y��80.��]7c'���� /����
��5��W��ɚ�~6�+����0)����@��A�Z��j��y�5�#a�sN$����,�t^���43�WBn�JgfI�����g��e�<ʵ"��3As��,
{p�>��Y���3�q!�os�հ�9.�I�'�2�6<�A��r
�p��R�Sy쐣��Oq(��A�A�:��2���/��	���(�x� ��Z:�M���+𛒳��d��m�%�������l���r1U J��Ā55��J��WnQ-ǗW���x�#�Q����
�-��[��{2�G�����(�ǽdmɰ4��i�U��.YA����9��]�O����5�x��"]'B�����*�%�;Ұ�'!U����ύ("�"S<��"��h�#a��ƞn(��_P��>e�gסL�����̵:{:����*d�R=y]S��!,��[���r��R���"��K�ǆ�'�8n!��QNF̨u��s;k����\�bjQZ�}��LG�#�a�mk�l���)��CLے`�ǒ�	&��!p�g	`��+��T�a���ML��#����fjC�aG�6�H�͒�f���#9��k�l�x�!1�\T}O,��-+�G֎��3�������r�u՞+W��V;�_x�qW���+F"au��[�ާ���  ��oQ�2�� Va4/a��c@V�o�?�R�]�'���7�� �	r=�2�5�_���gE�~ ��}T'N#)�n�%'J���$܈�`_6_�B��ߤ5Z�����~:p^��L�p�z��R{��-��V_����Q�Dهuٍ�Io�i+a[��Ic{���R"N��]dx����P��c���G���M��Nk����p�̎�2
P�q~O�R-���y���������?ɋ]�LSsH]�"�J�Ԉ���1��t���\�v����&����D����&�)e��{Tl�y�7��u��g6~�����;�1c������p�Y?~���m��\�+l���N�;����=�y�|7t� `4I]>����ȣ�2�� ���E��CO*��7�(aE'�2z$��-pp��D�N��H~#�Q+'�y��2i*�ң�BB z�p�/���.ocZ�.�u�ڥ�g�ˀ&x�5ۭtЕ�/`Q��k6"�!,2���Q�J��z�E��T�K$W���k�M(<�6$r�Gd���Xa鄅 �nH2��ܸ�.H�����¾Ʒ�����X����{P����6ݯ½3C��p16F��/�q�_B�/d��ILerO�u�?��Qap�"_������d�OuKb���ny�nt�X����}�6��M">Q��_?���N�^N�N���*3������0N�.�]F���75�@���2Ah��J�=����3�n�]�'A��T���2=�Z�߿�e0����������9���v݁��'���͙
=��z'�k�O��	�F�W������[��=P�Ji�;X�p����E��b�7SӔ)��o�����ђ�IT���&���ک5���	���� ��͔qj�>�޽�%͝�
$u��2����<^����T3��z�E��}�%���^C݈Ci���ux{*� z�^��"����	���	p������?�3�>��X$�,��z���)$f�أ7��1���;���f��Կ�?U��?�\Oiϭ��/`�uq/�%��[}��S&ݹ��}��Ѐ��AW�.�{������n�<=��ϔ4���7��V���|,?�X�;�li�Z�"�+o5U���J��uPנ��Z����s�׼��p�pDO��E�t�/��V�#�� �!sYU�k��)3���%K�ϸN�k�Bߩl�Y����vs�j���H���J�M$&���/Ī��c�l=��:��%��|ŋswC��K�*>�� ���JMk�#�P��� �oH���r��=�m~->��[���	�3��������b�rT%�u� c�P\'5��L>ƣ07�ȍ����abV7'� �������m�ʯ{��d|erƹZ�f��0U:y!tKْ����K�����(S٬��Z�����bW���x8����oh�ҭ�����a����<��3�2�H���|���B��iJ����/	�!(���Ӌ�Ǜ�1���z��}w̛���=�Z.��ӣ=�F�T"c:��n1��T�#�ЉA�/^?1W�MO��0�(-@(�Gg����n�jkn}޻�ka����4Ů=9�?h�nl��tc�k1r���wݏO�-�8Ǝ��]c$�
�hI��֧JC�q`��L�8��w���Gl�x?�&m��;��H��	̉���r�bj��8�,�!K��B�)�2�?QB��N�~hIl�tl�f����Ug�iz��5���*������I@Nd�r��a���W,�Kټ�0�k&R1ުQ��ss�ܾW�!�]�F�#��˽@1G�ou��i�|>�����F���P̡vo��iw��V7Ӕ�-����B��M^u�f�UZ�sc��Y.q��LG��q��v�{8Ɇ"f9�����\�hӈMf[ǻ+f���;���$Fj�Z*DUI��&�Y��3X��~@%�������+�5��`��H��4NE����n�Oq�E�~�0�g����+�OX%��Da$�@_�}n�[C�CIJ5~�޳LweӲ��0�N\Rth�&�}�6m������u�A7�v�7�A����$��i
�?�-�o�f�DO%"z���n��E�6�
v�Җ-�*���U���@%�Ek�.�,�*Q�#�"�o%�,��4Vc�c���Q��nJ5�Y��p��QK��h�d��ibWq���JK�b���d1��k�7�.ƴ�c0PxHo�P:�Ξ/��Ђ�q~]� ��q�Kо��(��ç�3���M�@���^M�����->B��#��'E�
���;��c�&���.�*�U��K~�(�w}��_��.�/�n�5��U¼t��DȦ��\ubP��"x������G6�m+�g\��$V�v4+��-üX���G��q9,�L�Uɞ�E.J�e� �Jv�	-s���b��"�{B]�	z@�}8!�����q����L��N3��T��� xw�\�Y��՜^\g����`c�DAE��:EQ����J�x��$�
�$�>���7��F�.�o�,j���L`�I�
��
q��?�/��ú�)�U	:��:�	 d���1ƉeO�Z|��ڄ���g��Mg�a�/��M�m�Y��ޚ(ju}���GּNz�WhM�.���(��Aό� �^%����M%����_����RB"dM�gU�p�@�X���^r+Zͳ�`���̔��G3���>B`ޔ���]�O�az�g@wT«���s=��p����[���� �BY	���N}���.$��1�*�p�k�	 �6F��_o�KF�?�)�߸�<Ȥ0�'x~�AJ��A�S׆x�������s�b�D�8~~)ɘf���S*�(��1n�}\�"�x?���ұr�n�B�(Y)�(�Y|^�D�'�]�E2'��� �U�xF���Qs��X/�77�9�m\Lې�@�f�A�5�w���g1t��봲�7�-=������O�1LX����2��*�u��#�h ����~�P��7Y�A�;�P�����Y�G�8�������ߴ�N�^Dg"�dR&m�!��O��>�,Ūt�GH���Ut��ܮ2>Ĉ���Rq]y��y�y�)��C�4�k����B�����i�Ԃ��ʼ�5<�ʨ��:2`�=��cx)��a�W�D߶�"D#Q���u$Y+x��Lp��B(@r^���8��@Nm�$g���ᩳ��AP��>���d��s��8�}�}�O�"���e��J���1F�'2l��M}��jbN��*� ���o�Ĺl��m���`�%/���U���n+���au�4�𲝓�s�Pq휯�I�Qu��n�����7���5�<����JА >�+�R>�gLu�iC�3480s帤�w+��>��H�5���W��?}5���e��vօ~�C��Q*n��ToMT�(���dV�y��r= 7%��0gS�/�,hL�^զ[��vSQQr�jW0��
���b�:�[���X�'��A$y;y��<��~/��/�Mr��T=:�Aʻh}������©d�X��Y\?��x�J�q�g� 5�+��RS�we�f	���Ԗ�gK<�%��Q6\��h�l�H����Bg37`�&�\��^�y ��(��������ɨ`�4h�;\�ӱ����mL��ay[ye���uo�V���Pf����MM�'N(jn[�����l%�Z��<���'�:կE�����6r�3ٷ�elD������o�E_Yo�k� s�|U{ח�9�)�?�԰kbC����7���H��Y~���;��*�ϥ~�$Ǳ(����{���c�>5�s�����L	3v[��(k��X��& n�d!?�3��w=۩L.%��I� ��W�ۅ��!�a���ѐp�����Db%�D{L�� �ԼXG���"�0M�*�wl�$F똧-�ɨ99�O �۟��h��v.��Z�`-]*���m��N��x�v��nl��pf;�y')�ᆧ(J�2�=�w#��ϓ�ʟ�u�5�����+�Pxu�u[�����3y�XF&)���v�h��9�,p9���#�]�iKih�w��Kx�"��Y0x�[1�A�ż�.D}�9���0��w��K} ���	m�pc�����.�ƆM3�C�5�ֶ b*v�)I���w� �,yU�A@c��I��zz�.�?�b�ٜ�����\���>�ƚ�PZ ]
d/u��ӕgp�m���Ӄ�A{�?2C+��jYs�����T�+�f�V
���R� g��I�$]g	�_<I,�v����$�erҒ.5/_I�͏0�պ�?�
1XaR�~�	�Fp(�)��ۼ�Ķ$;�ę; ��0����u!!D�5�Tvlb��`� �c&Ry~�@���4�V�@�tK��3(97��9�\�%7}��-G��c��!�0��mL���V�1���Vq�j
���/JY�"jm?)�;X���2ۯb�8��s/,�@$/�������~f/T����:�S��1�|��B��B��B�J���R���{1kZ
�����#�E�ͻ,b���#�7�9i	�%(2��Rm�\���c�f��Q
b
 :1�̛����Y��ih
�l����.}�^0� ؈r8�Uy��
��h��D��Z~{*�4���8�Pv�H��rbz��cKad��J�EG�jR�9[�K�$ݮ�&�}Ⰾ�h>�( ��r��V��B�-6(�����Ms�z��a�Z1N��#�����GW�:��8s���}6��D|N�YR����ؽ����3ns9���3m�A��u�]�h�EZ��NtA�y�Ҕh���������8p�8B�Bi�5�eU��8A�ꔝL
Щ���M�l�DÍ �.�6 �:��k�����`.�E�)v�.V>���m��������Η2��*�N���Ż�e�f��3{�FJd������Z�e\h�,���u��/K��ʂH���\��:�����V�I;���M������Ì>6�B�9|����8�|,�Ă�����#ŭD	hf�l�5�v;\T7�`�Dl�ګ���[��P��O��)	�}m�����k�6npvN�D�;�z.�*qL0�%�	�c>�b��q��c�?��ho��9����i9���x�<gA�>@l��@ ���/{jh��+��M�F�/h�	�_����0�_`��s��|�<x6�F]x��P)Z�_o#��{S~C�d�p����&\�G�(��Y.U�
��?�^�E��'���D�om�8!ղ� Y�J���sK����v�n{r��ή��L_]u*p&D���n�Х�@Vor�WZ�Ky߮�m�H�ҟ�)�T�m�^!�؏.ڧ�8*���Xpm����0��46��@�u1v ��hr��%�w�.!���׈ϵ�Ӓe�%O�������&@~U�A4͡���/g�������|6A���ݬ�XE�fL">����^�W|ș� �ӕX�;���)\A�d�XI�ٽa�����BR"=��QyS'%1�+<�r�����O����w�b�7�;i"�����w�ҩƿ�QK�~W�0&=�I�"���?Fp��,V.�h��_�$u��)\�r&���8��z+��`�`�ֱC�Z)�c�|Pm�(��|h��\�'L������׎!���|��{��
�1��;��Љ{���)7LT0�6�����o�!Dg���6p��X�[����^��Ϡ
�?Q �!iW���X	�*�ax�E�������H�!U��n�O�5Ipp�-'���pZ@\�L펁K���{���j�]D{'�O�q�7��4z�΁�W��ǹ�fA`���B�)��`�\t�Ȏ��� pt$L�p&�<�xEy\���*���ᐠJ������,���v�wKNt��ew(���W!�玷Y�����1�⭋D�3Qu����T�a�e�I�Z�����m���_2�գ�7m�B�Δ��xV&�%A�d��h�����
�P���]n)@�S��T�qbEO cJ&l�j��#��Z�!�&�1T�d4���g#�/��nB�F��J�����&U_��]j��23t�RQ�-���-��]}�U��O����qH8a[��킍��$���}�>6E�dWu��&>/ثL.�=��V������c4��R����О��`�4KT�5m�tz�X�*lz�}�g�1�pe�D���9Pm����[�g�ҷ�N1P
�EX�3�T]ȅ�e���: uO�����f�
�Q!�[���/2������z�]"�%❬��^�F�����NO��7��5�P������K��PmgTvN��SA*�~�	�.�Z5����.�'1V�����9������  *;M���J�1A��
E�� ZK�  �Oۈ@���ɫFk�y�jXVN)�5,ՅJ5��{s6����\�ô0�d�V��\�^{�>�-+t��
4�.l����bAs�8��2�R�%��rrb
:B�s�{cI-y��ڗ�5�bc�Ҙ$�M�m�����rM�ʚĲ�ve�0����t<.�˸q�}�ve|1���߸�S$�mꪔ�*�w��M�j�,/�O�s �T=��v��6C����\g,'Lg	GH�Xp��q߬��>���3 ��Q�� r��3��ϰ�� ����f��`_vB��2�D���9h��o�>R�|5��{���x*9��&l�8�}�p%�=#3��ʊ���U��6jŨEQ?��?�'[o��xN����-��"��᢭�+ZC]�b�[Y����i�4�#�D+�H�[)k��@��m.0eDK/����C�A�~��
M a�M�%a`�@�*��ʕ�͂�~��`�re׆h�^���h/ڶ]?"0U���GI�K'Ӽq=ѫ�Fx#m�\��oaƐ���@2,����F�z>�X��ꥊ|F�����+�8�����ԏ*�X
���,�\��6! �B�SwJ�#<�|���v~v�9yV�:�O�e�d;x#�ٯ⥘k0�)������bR�ǯ{5�m2L���� y.�"�#��5��VD�1[b1,�.��8���h�l"�%��Pm)N�w�/��Jx�S孒�߾�㫌(��V,5)��Q���utPu��m`�LO�L�=y��A�O�)��h��Bk�/I�M%ք��ͱ�LG>8������Z��0�8�4�Ҁ��[L}6��߶f��S��5;�1ݳ?��"u�ya�C������
��+|jmC+�6f	Z9:j��k:�5'�5�F��x��ȗnlq�aPI#&oК�Vf��N	`Yz��<
>޽��!�k· ZX��Ȭk)_��-�|�E�SL��18ӌ|��G�^t�l~�����?��N.��J�A��(TTp)_��S�s�ϔ� ;��E+%D����mp�9�KEU���t6 ��ӳ8X6��Q?S�B~�os;	��B4j5	�$���_O`�ǁǔp9�>�lb�k�yk�t��z��B�H�S�Q$%j�	4��T��1<�N�E�1���>ԆC>g������y8�Y	�ϋӹ5l�����T��&_�b�lO��&Wd-�̟��ݒ��� �%%���0!�een�ｙ���$,�[݂���8��񃾪��R^aw=(EK��s��H�-T�@EF���.��
XKo*�/���	͡5JBXآ�~��Q�N�_��q���m��ݍ�#�M0�!��
��i�͈�
�"R�d�Z�8}�;�p���e�V`��5�Ǹ�/C�|�Ui"U�����|e>�qO����̗P;>��ſ���4��f�Z<��� �N�u�5JM�&�Id7v�~�-��ـ}&z1?�k}BQBrK���/�L�әzl�A���4}�Q|S�t�`���m[��$�k�:�jja19[��U��F\ؑG�5�3S����y?���R�U#.��AN3���l�`�+��`l�x�1>�\�U��I�ܫ��!�/� ��\3�PtpY��Xp�a��S�O��M7Yl	|ֵ��܌~"$'�%�h�2<���0M-���OK ���,"f����Q��� .H��3�n��cm38�M��S0��k(�[䋌��R�����flPP\�	�v	�ҟ�~�w����9�J`��6~�A_T
'�"��ɝC�I$]�TOV@����Uk�D���O�g��v;��s0lr����x.��I�,k��|��w�ĵ �� J�$��MqsŶOW��+�����6�<O܅]�2@�)!���k��1��#8)v��EjA�%K
��8-�fI֩�#`�p���e��(-	&˿�KL��yɬ�K���3N��6�rP�Y��] :2{��P�i'u�3>�����s��ݢH��6���)�k��gnZ������K�$4��������A�D�!��'�yQ���vSo�:��_���t�	&5�9%b��w���Fm���zc�Çh(����ze��4�U5������"�>nV�7=mV�b�XEY<��h��%���ߞF�����)<e��0q�*�J 1���4��`��q�ò��õ��ͽ�*��S��)���T�d[����(�Wo8����-�\���f�ʤbj�nA�n���z���M�u�O��_pO_Pۑ�����|$�hٽ��6���2UlRd�%8~f6��aI��,����tս�C����]��5�
,Wq�����]<z�t��"��I4���I喣��?��N��!�zs�k�eŶr���s���.��qQ~"=�{�ϔH��ć{�}����?a�?����$�&�J{�T�à�Эb�fwD��e��V�nC�Q����5`�{�Z�| ��2"��e���_g��]��CZg0���?������1�F^�﬒G�L��<Y/幰Ո?g�l����z ��c�4�K�Ⱦ6+�-�Ji�E����>�0J\g���6l�8�X�����
KL��-+�Z�×8v��f�W��g���lS�̽׎���4~�v�Y�[�_���H5����[�ua{�����,���{�75��Z�e�J�b*�"Wŀ뒶}%5�����OT���=Bi#f�f���LW9M�4�^X���u�ND���u]���V��r��<��a����L�Ҕ@��w�÷��Z���#YVD���]g�S�D�I{�!��C]��2��5f��3SC�|�����Ԋ�)�zm�]��ڙm�q7��	hmz&�)S�f��H�0q���#ʝ����"�|�L�t+�:��am�|��t���Ⱦ@��w�2���e��t��5[=�Q��\���2x�S�&G��a�8"����{Xg<��zDdfz�kj��|�����s�!u��dG��mbjо�!ї�n�];
Vow���%p����0|��]y�Q>����9��-�6�a��N�q@�H�	������I��c��3��5��ϰo�9����ߩG�A��3�?��c��c^�$�>�޴U�	N4�ĵ-spA�X���/��=�l� .�@�ɓ�k�G2�������k��81Z�y.��2$mp_XP���5�]��XX>��;�����^��H���9���i
L}��p���� �{Al���"�T�q�++��K�㈟9w�n�ؿ�s�����@L�e�:�*��l������,c�J��+Қv|�Rz+���$Z��m��sP��Tw��h����5F���_�z����7��Xm�È,�w�-0я��lY��Q3�ή����l�N��?v���(_�	��Ǉjs{�J�
+�~,(OƲ�'��]�?,)yA8"X:�m⋦�DI* ��@��q�Ի�<�Q�������AhC:�y�6o(>X���/5�J53�X�	��Kֹ$b�M0��ܹ�&�V@��r�9e��B����E�'��~Ǚyr��&N�ע���Fׇ�NJ�>=Q<�@�ehr��������k���P�Ԏ�!��	��ﺡ���t8���k��b�wez����X�4�aoS\|e-뎾_�rHcx?l�l�Pyg �,��J�۹��'#[��S<$�d�����Aa���c��K�36�ǥ�)��Gv�Q|k�����P��cJ�~d����؄���j�.�M��bO���*�����L��C
H}�|�ߚ����s^C���
��EQB���Q���f�������8*��������g��o��%��Fd\]�P�
���'k���-�DO��ȧ� �c�G����B�,�m��י��L?7p[���5����F��{S<δ)��E��Ӳ��Paҁ+q'�I�����e.�YFQ��	g�~�]�02��>�uɣh�ÿ�(�΢�v��Xy��.e�D��I�+�˨��z	�Y���&E�x�J�hЗ�0�m�� �ZN�͘2��8�;��Qy"9��Hn"i�!�&|D<����%x7v�7�F���f[X�З3������r�4�����Ӻr�@$e6,j�a^^d	�q��SW�D7;���]U;M��Yw4#��HI���L�z�׬�K} *o�����GVJ��mK;d�RMQ 6TU>`N.YLs�d����ָ���h�
jc'0W���u����=g�9y6�o��>�C��;d�;�E�`�ۿoA.�e��w�t�5�s�4��q���L8�*�@�%�\�����������۪'�hӅ��s`v; ��w&���*�`����E�aCU׌lJVD,�ہ��͗��홅�ݏ�1 �	�,�j��&88<)�u�O���:*bu��X�wGF�[�������zH���=�]>�h��^���_7{�\�,�����lު�C����5 �3Jbv?5�m�԰)|ǎ��m T �y����*zM
П�a���]�w'�'{;���v�n�s�A\"_���:��P�[A(�T���E�B��Ľ_��n
��O%��	*Qd��'��֬	�5b���Ԣ�ϭ�� �� S�~��t�f�����>&�)~��Hh��%���T;i��?aM~dT��9dy�^~�LN��߂�䢱nly�V��<�V���,��/�*.F���!Ź�=���1v��fo������}�)�Г�#�Y�I�x7��C$|��8ZYH	F=�[Fk���3���so�n��W��'IC)�>ƞ��+
�Ss����AZ �R8�$����.\~|����tCr�["YǞ�9�A2���{�LE]7b0��"V@�xeF���I_C�����#�p~�K�d�jt�N[5��p�g��P��d����H��@�'�y���6�X��s8��N�}���G�5��T"\�)51�2��-Y����fm�y�\_��ɸy���~,|�#,x��n��q#/0�ԨI�B�fKr�����y��N#C��5?%TF�?�D_�sx�.��s��X�Y�wzfN��P��h�+Ø*?����b8�^wj�PA*��K坳F�� ���{t��V��g����0$�%���5x�H�i����{�b�`��>5OC�im�Ń����V��˳{
(��X˹�s�˒�Ol���C�k*��5}#mn�/UA���uB�u�doIh�f��u��I�;����������t)
��>W�b׃X,@��J_n9*�j�-��loh�3ly�g����p30l�V�)�lJ�*앴C�`�.q�hw�)8Ut�qS@O��\R��ޗ|�	m��Y�@&�����S'�8ֽ�̣j)~Dc�8K��,���6q�75a�2���m`�5���U���}��R��l<V&J�(v��{�� Mu#�#���9�~w��tTL��Ƃ9�O�0�~F��҅�s&:>S0���J$.��C�NPڭ���� E0kR6I`�ɐ$cE��Ghm�
ߠ��qeR휽��?�7�%��c������֩I�<4!����i�C~��X��4�e��.��YZ
Sw;��h~���ht�fs4�hL���h��z5e	�|�h�UFL�>V�{=Q�d�KSU��+��Er���ǖ>>&�9"4�*uAt�ે���<�b�`b�e�ֻU�MňU��WuƗ�_�]E�45��0D"1-�C�^��z��PJl�BP�8)o��.�a�Ǒ_����=[
��|u4'��SH?�p�L��߬Y�/kny|���L��_|v�[e��Ж���g��%�j<�vJM��?��3<;���EǑD�]����!�i�s����n����C�Z![2�AC�dm�H%�
�6�t���G�Ɂy� 9OU�I]��:��ꍽ���9��&�u����A=����2���d���>ۧ\�d>\�D��ߨ孛/��u�g��8G�5��u�Z</�L>��g��6D��3��bݵ�R�O��&9#\��3�NH���r�ٖ�F��(6|kT>��k>���T�ăD�������}���K�^�W�����]�-Xw��Wک�LHD���&*���~�G��)o�(�+#a}��K1��@w���(�Dx͇(`Ҍ��x���P=�0�K��S1�	��i�����p�I�>b�bD]��#5��3w�9cm��!���!�\��8	�:��'CC&�����ְ�1�KƁ��n��#c(d-�@������H�BXN�l���!�K<7Ag56����}�~�3D�yd&
�΂R�n�����"Nv_��G3$K�ئ0�>=�j�� dL�W��Bc���1utj�X"3R�����qo�wG��:��������,P���{��u޾0J�����5'���@u�?_@�ͦ�8�5�D���uP���КS��v�)��?�	�����/�<;	oU�O�l�	����b���ƞ�c��z�TA��ҪH�+-)���#ǔ�0����x��u*�s`�V�E�vn�,��Jjm�T�'I�*[�PS���Pd��s�����,=���kƥ��KiN��5u�m��k�����$Z����F��x>���j�b��k^m�!�5�1����m�̅VM����dF��H�@T�y�Z�
j^��y,f����@j��������>0��ɓ�`+�\�x�?�Fs��ܳA�%�=�Q,�m+�?���	��.��'[P�U�|RTvv��M��%i��m-���+d,4͕q�	��҄�4��Xv��(Cl$8�<�s#��Ya� ](i���bgi�����O��b��"�xÞ>P�Լ����zt����ȏ[�U 4���"���ɏ鶢M�0��W5r-a�¢X�I��%ڈC�z�j�����@�j��u��e�&`���l��0�d���Z�%!F䚈C
��dz����-*N���F������c��?y��hGn~��|�ׄP&�EG�9�g�P��idp���#����x����5�a%%/<�Va�Yj'�����lN�k!��"u������#0�O����+D�Ȋ��/u0���Sн�o�,0����X�y����ͮfj����y��&�t��?�n���#)�9��H��[��`��_q!�,��^��~����� 7�������ֵ��C�9ބ9�zƄ�1�f��F�:Yx����\óNr�)���;�������&�-� �X:����ŹBd�a�V���ՂTL`{�� K"W�BT��ѯnz.ɩ~@V��z�����w��9���SG�>}R]�&���0���D���j��8أX���;�_(pG�����98�{�q�`��z��b̼��(-�'�����j�A�а�*_Rѧ��ߛàh�>��4c�0Ѓ�o�V�l��t�r'⊣c|���:���h��g�����YWS���"�ٽoeY9Q�P��f'8'Z�X?��]�(���h���/�Ǭ�ND����7L�oH��tE_��	z�M*�5� ��@��y3��@L���y���Dz�:5���ߞh�|`�s�F
��8�&�Lp@։Gb| ���[��@��!�l��n�G*��@r&"<E�~/R6|��X���e2�������:9�i�|q΂�����Ün�y��=Y"�̍����v"�3���$m/��cyԣ�&�S�k���^�Q;71Cl��~�hB/��!�$���:ت3��ST������g}�h1�n��Sx��Q�$�䘫�� �y�����FA"���7��n�Q� (��qQg"(���K\�����z���3*���p�k��>�Z=E�}��B�O���qU�i�_�ۯ�&��挍M��+�%Q���Q%^���?�U��й~��$!7Se.VlYB(��9F��z�2X���5Fa�h�-��e�{?�� ���=���YȂw��P��8����Ǌ�U�ҟ��,$@>�Ju��@ˡ��Wm�
	ߠ�~a⩦��l7��ԟ�[��@��T`ŭ�N��c� ��r�U�.�z���s�'��d���F�E�>}+\XX�a��+���AC��=�����H������%ǼZq�d��M.3�Q�UF�����;b䋑T��C�M����{?������	���Q��|���0QH3�tL����h@*��h���̉�sc����E����7�O���\�{,(�?]����A�\�&�NS�l��.��F{�*�i�g��'�>`�qjt����Z�j��YF�'�}�E��s2����4�U/���-o�:�Jx�N#�k�JdlF�':a�-@��m��aGa�X��.P��m�" �޴X��e��v��8���+r��%ݜ*M`���4�]N���5������>�����2p���Nٛ��U�SSi�%2�C�Ru�}:LA7)9�3�Mx�w���O�źz���R����Z�s ?���E(��Z3P�^���D�k��ڡ����~�.дJ�<��[ �<��eh}����'/G_8�԰h�
�Ưͷ#���>zn�=�<��茕$jQ������\B��&z�T��࠺���������#(��{�z��d����u!�㘖N*�=��=��Zd�Q��N���~�L��b7G�eS{Bp[S���d�Q��&X)-�Е��k��B#�OCJ��\��f�0� �v<�L*,��l�+PS���\���x!�S+�..MW����Z������C��)P��D��@�Ƀ�E Z�#�:��ȶ�{���a����3�e�K	W���6�C$ὍB���ݳZ�,��qӵ��V�3��ʹFE���@��~g�50я��f�	zr⤎"�Hm�Hyv=hIg;�(�����������<3|����U�▲�s���4�#���bkV�#�_o� B[o���}�I�YԀZn�aB���`]ד v�`�����L�,������-8%PH^�/����"E�4��%�Fdo[ʠ�D.�i��$!������"���Dr�ٚsO<3/�bx�`��.�
*�M�*�a�Eie�c��L�9g��Un��W�e�0Xհ�žO8]Y2~$9X�(dՀ�N��{�4��q���i��*��6۵��D1��q�,�~Q�9�[.m4Y7�N��0�eA���(�H�S/c-�����f�����S�7���7\���ĳ�d�#v �8yB3���3T�~�C(����`XJ��hA߄^y�Øھ����q �
��Ħ�k�hS��A��{._<v6UeĈ���q&�q��e(N��/N\�GXҦ�@/��1��������`L�fN\�J�+���Ln�9.�DS�۬�e��Ǥ�-�Z���	lɴ=b�a85 �� ���D�h&�9��1S����i��KTƏ$�Tr��x�h`��,���̯T鉋4�`\������~�V~
��Rʉ�H$"9�!9|g�0��tnZ$��{���=1�/�H0������=C`w�]���1����ֲ=�蘡��x �)��T03L���	%>�Λ��3Bu�5࣫Z���@�t��m1"�B3���-2����v4���9�ڽ(]�x������{2�q]���m(|j+��m���Ci��G`mņ(�YX:�ǳ����.����͗($y�3�n����_�=:���
��U�m��ZC��R�Ӝ=1=z�2��Q
y�\�6�4	�gGdE�S��W��n��?�>�yP����̰��ќ�/�`@m�����_�s4|���PV~�Px�0|��R]����c�'�Rث![���ɿ�u�$h?�n�S � �?ƥ��e�ID�Bri�"hUz���lߪ�/�K}g�|�tCX������h�D����!��Ġ�����&)f����t�kӣ�pG���� 	�Z
�$�\aw���eA������/���T�Me>H[��j#
�*CTT�m���]�~d�b�� ��cSX��WF�@e*_��a㰲�vU�т���YV�D/5�N�V�WEU�ޖ�~����5��̱��c;ZQ��8l�=�V�1E������M��5��'ɲ�qa�~X�	\%fي�|���e	}�����1������i�i�#���z�06 /�`%i:2l�{;��r��ଅ��ڒ�\��&$*B�@�r*��`R�pv��Չ���h�E]��S�k�C�(�>��r<�@#�+<��B;/&WԒ9]�&�U8�S��y��/G3����J1�KP6�KI�'̬�iʶ/�_2������9:F 1��'��UEA��KZY�#D�[4\¼*�ȍ�D+���#N�p��YlfҔ�Z�y�U�2y���Z��n=||�1�i�pd��5M�n�Po���R/Qc-�}��fbK����m���$��Mh��>z4�����������8��Q)���Lq���ߦh.�H- j�Mu^�\�Y�۷R�B8��5.[�5�����U���Y��e`������'=�����m�1��A��IXǚ{GF�ȑzgg�З
���/��硺�UK�`�x�`p�BG�?���ˬ���~����wɩ$��K�0w����W�����g]�|�|`vⶖ�*����~sP��g�+Z���-��3�����^�r�һ�mU�;A�q�2��Ʌ�����A��YC�0(H��*���5�ț2n{��1��c1���Ma/QF��w�K�4��̩ӿ��8�.<�"+N��횝�l��t۫���
}�c��
����A6�	�T���#�U��6���֊zJ ੹0���(��KLfhހ���x�z�Z���*ұf1�yf&�y�W��!~[��*a�����85�7����+���J��(�FM)��T1z�a�7`d�� q���)�C���`�n��f3���O�a�kj��9P-BV�5�F-HڶsL�؞��.��E��F��{? /�fp��e9������(���L(���F&`�b�����/��$¢�ڨ��lAM
��j���6�NÇs�-�pڬ��ۯ��`���#�J�~��؂�Gd��<!�_�ҊxfA�u	��;Fe���� �9'�\�p'��'Q��R���zM?9�Q���SסO��/ً2L�����H����x�
�w�8CXk<����D�A���S˔p�&c��<܅dO~&��"m˖�����(�%�ݰ ]�ݥ�j	�k��^�k��&��:L��@��9X(ɐ����M��F����d����H��9�E�	�ɅN�y��+Y�ו��F/g]8�@��y�T�]�v����,���eZc\�&�/�y`��º����lf��yV������P�`��38�#�o�xt���s���?�g��SPקZ�5[G)k�Ñ�¬n���pg\S�f��[vȨ	�p�j$ ��K��օ+m�,f��l��C�:3
��'W�l�4����y*�Qz�N�Z�� s�~�>L'�0�j*����[�|8�Q���N��J�;�,v`T�a���;u�y$�J����a��7�>惄lM�5�(P)�._���n
/�WE")'�)�/R�=�+c��"ɷ��Dc'\X�%�w���\��F���=H��[�P	��㴧`����
�f'����{`��L�#��5�ADzZ�J�\(O'	{U���f�v^�v��oiu��7[���Bm6<��x�]��j���1õ�L4r;���;!U��Zs/ F��%��&8xf�
@�.��C0d�J~~�12�n��>�,*�"
E�2̿]��	�Z
ULa'�Qe�_��w3���L�Q��GS���IsF�F]Y���3�I�j��LG<��}zzPE��O�:��jؒ��(����^����x�G�ZɌ}�׵ʆ��dUi(W�խ���V�u�1�,۰�G@��l�PӁ�:��:?��<����h:��w����+ǣ� ���-"H4j����C�J.��ǝ�+�ݶ�&���->{Q�@n�Q�#k\�(��T���1RpSx�;�� `H�94joi$��-Zs�p��Ze�~��ģ�/��"1/庀	�3l�X��N�B�Q$�*�N=$jc�BaX�u�2��}���-^��6������-�\�+3-`eӎ�(�4x�؝i���&�+C�W�wsX�{I z�3�����]=	�+�a�Uŵ��N	�ϑ��+��e �xt@n����\�a*�^B^S�û����#_��I�{�����4���`��D�����I;W����	��b��.�2.,�ec\R'L!<��͎�%�1Jq?B�0�ɪa0�4Gd�]2M�7�
�%wR9�׷ѻL�E&��^��7���$iz)�q����:�w�A2�ݒ��� YG�G���=W���R�zp��x��>9
ƙk��?0����m��[�o�J�������6y�g�&ZquL���nB���NxY�|!v���`��� �,�O�
zW;щ���iD�#Ḏ�W���şt෮�&Fn5��0KE.?m玄eQ�&5�t�HPM�[t�����Kݵq�F-�$/�+zgtǀF�n���wg�-�4�f�]�\� ��]0��HW�W�D$Ϫ|$?���-Il��}�n�����J��^��.�@���oҟY+T��`*� �����Z��!<�+`�Ƿ�U�ll��\���;����ïW9��DK����Q��m&���KR��%�0���9�$��Lj��$W�J`-L�	�q=O|�c�Χ�>�1wCm,M
�31� ��"WZ���]2��ͧ����5L��DmF){Ps7�x1GeYN���	���*�H^@-^��(ӄ��ЍR�I��y�Z@g��+T��x-���z���\�X[��p0�89�s=)����Ֆ�@��B'���KO�;4��O��MRHE\p��m�j�P���	�%I�H5Scrpuw>O4�{.~+J(+`�q?`uؕ���ol0�[O���>5hF�æS7����Rڦ_"~�M��n��;�qKڏ���|���4�����w^�F�Ӷ� ���6<�dQl�ׅm�Sh��QHP��O�t�Dgſj�m�[��}��hZ�&��[�^w�d;N�E��T~|�C���_�$U�F;�����|�i�T���"Rx��t��::�]�pq ���cd,�������ڧ���ղ��mi洜�TR;R{����8VB�-_\���V��܆���ש���p[j�c%�@��N��9���\�9���t�H�4����n��g�Ն<���v޼BR�F*���� ��s�AI��-�<\��#B�6	*�����~�!�.��z��	m`�A��A���%Ź���͊�/Ð�&�~��|%�X�X�Ӗ�hB"j���>�e�&s�s�b�!S�sUZB��Q2=��_�`9���� ,�E��.(�>	�Q7�^
/i��ς�ˠ���1���Zb��a�(�jzF�F�� ����ňݦ(�3g����(1���iz%~�( �c���@F`m�Wz�H���� �xb�}�V{A�����F�h��L��<*�OR��%�ĶRZ%�������_�,.�-9W.���ci)I ˨�b��B���Dc*,Ї��0a{#�,_�����<���ߜ��궮H�����k7y��E�%~�G�	�!Q�a'O�k޵hI�N|�G%�0�F4U�܅(+ܠ$a��a�j�o��l�>�6���i�)�D���������woN������w
��U�L�d2o?l�o}�KzE���/Fy����+����b��/�6f��{��yC��]}����|�?��^[��8��]�m�k�`���|;&c��:q�aHd����� �!�\�4����Npʻ���֜�S�&��d�V�߅������N�40I3y��u���vG���.�oKi*�˦�f�(�m�����-��B�8�Jڰ��h�"��
K�ܖ���U%��JV�>uW��PA���rv��e{LMȅZ$����fc$�ŝ�{�
�?�
��%��L�+ �����B�K7-�D*��"�8�F�bu��b����W��Yf�`.����Ev�8��\�P�������v[	�!e�.D�(P�Iע�,���Ų�����|�2_M��b��H��0M���-M%�AY-�0��N>��;��sv����0���S�_f�ɕ9��Z�+��=?��[L}�j9�? �/�����Y�=���|���ч>��in��7��[�@��C�Ҍ�`�:��_�&'��'|`��&W�s��5�w�I���v2��F5��D �E��ԚV�P����fq�:��� k�#��3�ϗF��� ����ȇ���<I$]l�p�#�a����C�Գ�����c�cM�-:������Y2a�TW�8w�e1������U�n���?�׸���,L>���%'�'��ր�@d9]|�4�n�6Ѿ$��Ŀ�R��,2|�)�1�������X�"�ڀ� ���qtl>���x�����ڠ��0lӁ��"�]�fo�ڶ���2�^��'�V�|��F}�n���EN���G�?K�C����I��s��M��Ƭ��᷃�e�r�|0D�w^��I�B>�EP{�⢲gI�d��j+TC�ַW���8l끺�i�����7����N�<D&�),( ��ɛ��Z9Z\�\����}��a�[N%)�o%}8);�؏J��v�|@�$T��A�p���]�&����o��.ʲ�O�2�IFA��O�"��:��+��c�.�3���k���^ZL���ZNZta�M�'�;���[-+b&v�e��^#�}ߊJ�sIp&|*�G+��8�9�,�W e��	W0 iV�cL�<�<0D/��hR�Q�۱'��Of�9����N��3��Gs0s~W�I��P���oQGЍi�?�Z��H�Tԉ8\jn�+��1g5f��
�`�Oޓ���3�^X�`�u���m,)ð#���v0�~G��㵟������zQ��4 �*f�w��V����?�uk
1��z���L_�tF��
R֚�Y�*ʩ	㶘
��y_8)T�j�B�#��ё��B���pl��
9!�ۘ^o[����
qksr����}|����gt�b�ǁtȱ�,��;B�"���:�1f	C� o�Q���i'H��ńf!�M'a�CSb�Ը�JJ�H���
D��֐�L6�T]G���%�P��|�5�Vj@�v�ﾤݪ�G�=�\`j��a�D�|k%�SA)�.X��8ɻ�G<��8;KSiUB+x��m�aW/$;����]j�9�|D�Z�0���3p-Qս�Q����[����">��7�{F^��aR���$�#�Ó-�ۖ���||�����
�L1�U��M�sKnyn	}�N�PE�T&9=hO�#�v��_[WFL�J
i�MP����#sc:�����+�4�o�2W�bB�"�k2���X+��T,DI%��uAiK�r_)���j��"�F']�Z��_D��1��N6�w�,���Nt�j���'x��$F3h,t�*�j�뾡ie8�\�@K>]'*�U�Pݕ{'�):�P�;ʴu�SrY%K*�{����'rN>�o���#e�"�R��wH%co��7�B�k	�(���N���_қ�,֪�@��)�T�����Q��Sl�Y}�E�b�m5"��-Ww�R��G�T9Mc����B�~�j�eY/��_�
v@?\	25䉀Q�ڲ�~��'���:,T������[`��r����]�K%�&5$�Q��G[�UD�����7l����{���͓9�s\�SK��ԍj�7O�=�H@���:Xr�T*�D��]��WV�k��ݼ��84E� ���^ْ�Mϫ�)�('�����$m�ߚ3<��S����ߕī�j�s�YSf�֫�1�Wd�N�/i 5u	߹��ᗳ�r�촲<��+13��߮�0Zx��y)Jc"�:)��,%2����Mk��O�q9�ME�K�Su�7��!}��3�ֺ�Lp]"I��'�U���,�% �\�Wcztd���Y�'�&N�vy{��AJM--*%ԸChW���l��'�����t2z���ե"�lë�C�МGS��MU�%$5%��;٨DQ��Oic�== ��kUp�I��M�g��ڝ��!qBӿ(���Yc���5�.�����zm���8� 3�g8c��޾4n�L����j��p+��I�:����aa)0��ū~�z�l�7O{,]#EDސ�����?��}ꃍ�X&F�2�G�f� !�ˏǂi�l���;�~���\&a6��@�3c`|�U&p�s�WN<�'�8ʕ�R��b�v�	�8P�Nm_$E*����(�!A���(p����ӂo�/���R�[��� �c��C��S),%���ҭZ, Ji�V�h�ظh-�lW��$QO��f�(-��Z�r*��kZ��ū�@�`0�f^���XMGOi��<;'ճYk�L�i(������&N���0DF$D��7��@%�|R;?@���3�4�d�H|ҷ�q���|�z��7ӆ�f�cj�`Y�:`�&� ��G����X�XM���V��P�Z�a ��l���H$�u���n�W�zP۶��3&��9�%V���3Y���,��Ns��;j�O��l�Bb�{�qmv���	_�m�;Z��4ҁhߒ�Ҩ�R��tmL����*5����C�=�o(1��L[|�z~̣V}�s�M��x4��ya�mNŵ��w��q�u������c
qT�������Y	������K԰�`+���ä@��R�NM�Bo#�:K-g�Zˡ�J�wr�g�bI�t)06�9���t���bM���N����2
��������P��Z']5w�)��DH�5F1>t�[
8�Sz��,�x��߮�z�V��eM�R���r)� y�|$�d�6������SN�6�}.z�q9�V/R�{ُ
�Y���C �2\�}�G�4&�`77���7~ٰ��K�f�박z����gsC3bV�A�ڼnɻ/��!'��)��x[ꅧ�B@�aזZ��ͻG�x��I�Aq�������{].�����m�=��� �%�~�S/����?�I &������O�zY������Am��{^��?�(?y)6	*QvmCG�Q'{�Ή��,��������蚔%)V��6�����Q �J��I 7f�z��<�:<wb��S��"h���<��YA0�R%� �!9(�e:�:�7�K�N����8��'E��h�>�%N��~�H��7%�� n����(��?~�YŢ�6�OC�Qr�����J�'m2�+H��� 3v!,��`/����yo3'���q�[[Y�|�����Α�"�,R�XH'�c�l\��9@P����N�'�u�:SM!�T���>�[�,WqI���)Z=����`������
�|8�b���#��b|#t�����
2DO��3�7�����:P���G�um�� l[c��7]Apy�z=�����'��\R^���5�5�Y��4�1r��zigPԴ��4F�/���+9F�ls|e?|G-��ӭ=�z�$o�㘻�\��Gf}S���D�T$V&z��<�׏HR�e��K�]2/<�fshLk��O">yȢ;S�.�3 >`:������X�)oOU�i+���}vV�u�W���`�N�5KI�����R�g$WaU��BV��P�$��hR7���}�;|���3 b��q�*2���n�X/�c�E3����q�t�u%�0'/*�`��h}=�ú��vϝ��Dc۴v��m(YU�7�jl���^���%��D�8��P雓u�h	3����9��9�4�����9@x�~T=o�,��K	�J�`�ZB;bY��V����k���V^q-!f��Mݶl:;v�s��m���Y�DO� d�"�&6es.] �k�A϶Vd�`=���G@��d*�Z�q#.�������V���J�4-V[Đ|���}�����+$��B#�Z��CY�kZQl_Pj�����"1ޤ�at�����QS����q���,qJh�p�l�y��ϲ90T����Y�|�\�_����O~��/���V)'�Aԧ�x���� ��.@�/�d����N\D�dK� �����7�0���/�
$鞩�n��f˛ԯ6<٥ܤ)m>���ʙkj�r�6��� yF;����I��8�?�
'��p�ȹ�I��?:��8�˪|l��ۨ���p�:�������a�ׄ��/m��Q�jN�[֠���G��~��b}����4�@^sőf{�_�yb9�W��9yַ��_)f��,���s�I2�v�G�p��s�!\@�c����J)%1�w��v)7J���-���j�Z�r-��2^�������`��������nhmZT�5����ga�S�OP�Y���.�0Œ�c������>�j��6�,_����{3���ݪt�1�%�����d�J�%XM�J��G?�8�XK �.������U�^�%��J�Y�X8S���Am�����'
h+yo�RbC�Y�Y/��_s�W)�E��e�:��/T��\&Z�-���(ù���i����y�l@�#��K�[���Œp�Mg��i>]�����f�{$ssU_�4�^>{k
T�A#�������&/f���qM{��%D�,^/fɜ���p<>�E�X�'| �
+xN�^�$�˽:��Ba{�-��m5g�R�+|��Ɣ������ �~/Y'�>$Oۨ�	���1��95z1��Î*��_��7��1�+�I�Ikz����K1*�����U.o�����������<�L-5<�Z+L`����A�їU�&��V��A<I|M��"�-��SԳ*3ze�wG�/j��l>(����jXC�R&9��qUQ�A�w��s�4�_E����.Ry�3�"�M��%�ұ�E͓bHrQ��CS��@񦫴�]�oZ������js�����|�^��wP��k�ዌ@�s��WM���L�U���n�o�(�}����
:d< ��d� 1�)&�Q����ҁ���� 4�d�U3��_�����>�̝��?�F�q�������/�����P.Bh�Ҕ���m8>��@;����ݒWd�+��<���Hש�K��ۻ ��[ޤĖ3�B7Ŷ�o�����U0|��Fe��h���	V��k6+q�DD�К�����
D��@�|��?���t��o��DwJ��O:�x�0&ԐN��64O�G�oV���D���	�����ߣ��:�vK�<��"�)�^������Eӧf@��D�"��vAo�O��eEYX��9r���P����Y���))޵��P��Y<�Ԅ�3��A������g��x+b���)Ky��$�a����ew�KM�D�rVw7�xV"��(��>p.�:?�mWc�ƱK<aL@fs�( ��VH'p;<^QМI=`BH������9�Z�y�jh� ��uU G��TϚ;� �4�7�a���\s�6>^A�N�,U�De|��4銲	�ҞY:�[m��q�>����1��7ۄ�"�2�d.����m�U��?�. ]�&,��Nd@U�<���!&�S��:�&6$��Y�bˊ#1��H��7CK���.n-g��$nAphoaʻ.<��K�pL͂OE]��m���
��|/�ۉE�t�wJ�5к��:Ĭ�ZJyi%!�[���*���\�3ZVZ�*>��o2e��$_���)S2�g׋���X���)!0���cmX�r� Ny��\��=�Y����4�^ꊲk��P��н�HHq�U~���[��Ο[ Ӳ��eX9.�8�K�,�x�4I��u2&�Q��%��NȞ�s{
�Q��e��ǘ��c�9�_�gLlrֹ╇�2/ج������o��s�䃅�z��%����q-;�9e��7j�%$Cu���nt�##��ժ��>�Ⲯ
!;�Q��X2G�m�e�t�F{�c4ȚG�4�k���!�{h�����C�O��e�O_��6�+�o�Ȫ+l�^��-��7s�ud�n{�%L$,�i5+����3����`�Fr��S�������~��
��%�p���T��R�gx ոض�ٖ�l����7V˫�P���!�G��M��v��7,`ҭ�&�f�#��BkTS\�w֗�H���oh��O^޻6�Ŝ�lVt��Le���5S��"�����cb��Av��}g�67��	�_�C1,��<���yc�.��t:�_��!���j���cv���6g��}^��ps�ƀ�E��H$�=�[��Bٝ;�K'g�U� ����+�+��G6��a��xj	��(������
2bS�n�?5�L?�-�q�5-�oލ϶���r/���no!���m��7�'��S�PPq��,�Ҏ��%�����%$CwV�W�$�J�t��{�����Ex{��+E�	c.H��b?^puE���d��Q�>DK�U��?FnѥZ=؟Hj.�nP4UP��^���4��;`��K�7�\MN��6X�jE�[��/� `E0���L��V�3��JQ JF=��_YХ$8�\��]�Z�m�<y	����ב���"��-����K��>O�����
����C��[�߽I�>� ��Jy_�)���L].� ��8��X��3wa;��5d�7���F�ne:PϮ>���/��:� ��ј�ad�/=�PW��R�h�?v�)�5�ċT�%�z�ܲ�8�U��Fܿ�s�o)�3~轭N��*-626:T��ҏem*J	���I�z�ݺ�7v�I
7ޗ m��*娹p��O0(�Ap� �f#9笂�1g6��xcD ���l���D4�Ha�IIF�kOV.�Q}L\�=�5K�E#^S�������īzW�:�)��iN��ઐS�#i�Ihݦ^/�V+��E����^M ��[f��_�$�������FY��=\�1~�P���e���fr0��<'$o)��Wl�{�~���+�F3����܂]D�/9q[5�?�N*�X
�:fMd�1���!���v�St@N���	g���U��tr��ה�N���� s���~�#w�$.���C�QF�kC&u�-���ok�og��JX�iN�ܩCw�Fl��Jr�#�8j���>�	���M�C ��:?	@2�J݂�Z�������O�~�Ͻ�rI� ��c�R�9�nW�U>ooL��U�b;�'@f��j�#ńw�ح6����Y�f��yv��w�~�&�A�{�Z����z�ޜŅ`�9Eo�A��(�m�?�B��mn�S�'� ��;P)��3t��T����G�M���e�TqnXy���tL�C&�EK5����#�{�x�� ԕ5�"���A�"@D͔��>�.���L����tB��,�8��w�^��J�H�޸|H�;�i��֏�9n��K>����T�H��0N-�e��*�ei;K�O�Q}8_�F�"nc��ƣ#ܙ��M�>9/ч^�)��|����s�h��i��X�����NK�u��j$�1��Do&@�̾��|��XHߘW��=���˚i�.�_q�G-(�`���o����I�?`k�X�$�����jv�٠������)w�V���:8X�t�
���%�wH-[g��B-!��~*�L��&J�凉����R^�B�pa�_v@X�IҪM��-��=�^�lvO�gd���_׉��qR�-$��[AY<D��EQ��Q���Ns$��'LqǡY�8��HX��F�o�K���c&Ūץp��Y����.�f{/a�N�eI��G�Dk�5��c���4�l7qԠ�Ć�@�Dd���%3k	��!�$���9׷�`�u ��ւ��oO�Av��V~��:h��k.���+d�a����~=]Z��{��6�U�m7c&���y�5j<.��|�����8�u�,s�����X5;�?1��^ ~F���
֪���E����=�/�#��qu��Z�E����j'�ȦD�갌�Y8vr��iv����ؠ������M՟������t��d
_�!w�߼FA)��,�g�Wd���p��}��:1.�˓/���i�D���P�).YVK�>:8P#���5�-�%�V��6����z:^5џ)�P�T����A��D�'��5l0�( �X��D�������vVQ���%����:O��@w:��J[)��>Ȑ�*�_��f�:���W��9$y�J�U9����#4���=��@Q�<��+�Σw�e�Y+
8c)>��N�z䒟�:Gh���*����eJ+C�_��Npa�"�B�pvG�u\h�)],(�wKh����:6rˣШ6��*��ٴ(1P��v�9E�|�J�K@�#C׽,Y��(�}��i��Y �^Q\�%�Ä���6#$�*W��l��hy�PT�����X�KU�JE�#���h����V<�w� ��/w�i�m/����׀�su����Ԩǁ������q�T.�[�	�s:��]/:7����٦�BV!�6�"a'#	�y>�.lh�-4��X�7i�r�-���yNM�^�b|_˺���r}�n�m�����W��\�c-�{��:kHބS��m� ��g���C��Cv��X/�Fy��K����_��p�x��<<���R���)}�qP��g��O��7Ԏ�(]ڧ�%4�1Y{��x�me�6"G�8�+����t�"���E&��G�!-�G�i��8�Xjf�\��B<����p����3U����f���s5��0`�v�Z��6<�������_���� =UsiM(�t��VdB�#�>S��+_*�F�\�wJW��@�6y"�*?�nC��K/�_� �=��Z������Op�Cb�X���������&��;�\c���TΉ�����1.l�&�����]
������֗b;�T�2�3<�@�\p(�M��_�v���M��R�[P��j7�G���R���z9���p���u"6��� �� �B�\��3�w)np8
��R����|̮�A���c�:eo�pF`b�R��ۅ����{�)��Q>f_�2�rڠ�����|,´��Ir���*A?���1��Q�~��r�`3WޟC���]^�J�E��E�SG�9�>U�:�`�{�n�}�3��}�[o�Q>؝�q�X[^�������R;#:f�CS00�.�>� (�x�ʗ%�Hw����y�8��vGxX��ѐ��&.�e�:�[���'Ԓ�k3y���+���ш"�#�2�A��vn ́@���k��s�,��w�g@�<��G)��� C�<g��[��jp�H*�(7��� �0��{>�x9G�x��u�J	m=�q�,-ݕ���:/���D�H�_��"D!
7tr��ڀ�k�{�N}c}�w�h%��͎np��H��	��6z��m�ո��r���ůn��7�t��~��O��o�0��H:���N��+E��K�L
���>��oFpT�oq��4�YWs
bbF-���"�Z �FiV}8�Ӎ��yS����oY�G�������RL��;�ǅ�E�<iخF�1�K5���;����z^�G,)qυ��j��R
n�$my(����5��E೘�ɧ@k��K���Bm�?h�R��&cR<9H�ˀ���+������|*Ȩ���>�Ui����Pgq�|+��l'`$�ͦ+Q>$(�<7������J6��LΙ5+��=�.��1 ��(� �����R��*���k,8�ۿ)7��C<&��u�@�!bJ(b��,���;�׻�}Y�������_���
\���=.uO�`~�&3����O � ջ���U����3��y~�?�!b�Oۜk�ʛ����}H��S!p�C�A^<��0u񮕚�"S�wZ�\�
�����װ�iXzaZz/��0
��P�ha��7�������@n���#~Hy�m�Ă�c&7_�اCXaU�>#wՐ�;����y$�+Zo��v<+f nb?��G۽��"��|���ʩa��nz�l��4��Z�ti�`?/��^�{�hFn��&cߑ�HnQ�����u",c	hkʮ�}�4ʞd@=9�)!ϒ+�g:)�Υ��h	���������>�&Xa�I�o�Z�CԊ�T3]><ն�Xm�m9�5�%�̍s~vV�Q�E���K��v�Ԯ-.����@iت�2g*��2�e��o�@VϺ��ϵ?��h!S�a�f�YK�HF�J42���WH<t��0rۋJ;qZ�\
�g߄_밲�ә�3X]	J��$��o-\�~c�P�a�>�w��"�_*G��Q�$h�����ɨ�䦮�c�t�����z9T2���e�Z�eD��|Wy�Ke�F'^�,͟Dʋ�A�A�����e;z^��eۡ�R�����,�c���wp�o�wP/bI&�����"28E��.zp� �����O�>N\X�QP�q���lO��_PU!�P���>뼦�����e��~U�����U��%���ad�z�R7�P��W��f�r�]h��Q�5������
ׯ4TyR�Uf�dG�۔��qF`����Ӓ�������&�xxB�}�~G���r\��14·`��-��mߑNSê��B��	���T[�}s�Nh��.�0<I�6�;��6#����*A��]|��d���e�qW|��;�F�&qeL��s�$��tI:s��x�k�β�u����H[�/��p��p�y3XJN�L�2�V������vE3�^�~n�r� S����W������&6���!�b�8k��u��6�k�r��dmga����Ģl<��J�ޖ�� �����r��_�؄�� S��[���9��Mp$�U�j��	�6� �s�TU�F`:�VP����\��A��+=�ʈ�0��rD�:�������y�Gz�jM���{149��a9��>CY�W�ߔ�3����w]��S��k�[X�lk<�!�R�V!3ul�		���v��e4M~
����������U��f��R����Gs�*��F4��wn��ֿ�_�3w'��F�#�i��Dp�n���ܾ��@�\���7�/�I�8����ľ-�%oQRnv�<F�����ɠ,��|MME��o��'�����]1�H{�+.���i��2�1�>���Eኌ���Xy�.�/vp�B�\8�k�2��烝���a:|& ��)L�P?�
]�����}�d�/x�"?�v�j��@�,݉n+��ǍP�?�%�w�Bz��4����8��K��V�t���d��������G��=ȳ��.3<������Μ�~2�P��G;;F��)���#��D#�*!������,���<�W���I�!�6Z��!x�B���A(m�d:!Y�̶�1*y�4u<�R=�D�|��}�;����Z���L-�IѺGv�vj�LZ��㧑3! Ό�$��� =�W�����@�m늶��u&�7zDso��5�S�{�tLs ޜM����I��h��1C��[>K;/�<݋,ʴۑ�Pm�y��a�~����pw'�V�X@�<��kY/���<��(������q�����x�a����}cxںMDz���ٹG���po�є���Alr��`�}d(��{��ۥg'�VS�k�De�ձ�K�DD�K15�DcKC��Lelu	��l���Yi�4bc�t�C~�&N�r�o�K^}"Xě뇩�&?�z�P\�O/����b*��f�O�~��X�+K X��TnT�y����%?A&��K\׌���CHw1��7*�l������.�-�~Z}��'���%������b��Rn51Y����7���i3^1IN-?�#���T�"x�@�e0�J?|#RO�6�y�P�D�bm���k��S�Ψ��h��ނ<`�Qo2�u���P`L�D�{|��>��}��7�9o ���1�����1@שT*х�|���:!�����|ȳך��z�[�?�: ������vH�P�m_�2�T����d�(h?���='蚄BW�K)� V��ͧ{�"~��|��Dq~������L�yF��!�1��6��p[U-��C�qx1�3���V�_�'��6Y����a0g�l�E��h�KH��w�L�&���*��4C:A��jJ�U��Y�憨zF��+�Y�L�!�5�\��z�!�^���2"���QJ����<��O��;����ZB6^�H�1�$D���_S����L�(2�w�h8N.eTq���@�*�����&�`�ם��띳	Nh��*>t,)�x�����8F~^t�&�/��L��0g��4�5�,E9��	�:��WLr������6��U8h�`cS{�� 3A9��?�y��WL�Z.T��v2�=V&!���S��l �ҫѸ�fAs�@��ra��;2m���}HE�aD��(F��?3�A��Fⱅ��"�J�a���$�����`}]C?�d*L��#Y��=U��������_|�lwFo谜~Z��E�ҞA�$֦],��u�{�f�!�ؒA�/̀8j�Rk*40Z(��<`Յ�p��T�A�ݵ�͗�.ƛ>��f��'�8�r�����-�Ô(ϸE�ڧ��1�$�Py���諗�JپtE�J��1�a�ʕŁo���4ٺޏ:cGJ��h�ȺZ���S�aJ��{ �g��B��}�I$(ს$A�:Xj2�V�(��i�T�n�%��A��o��O~[b˒� �1ώ��V��N����Tbv1�Ğ� ��h�Y���;
�E^�%?jO�r�1��,ڸ��ͦN�Da�e)OZ��:�8d7$��i�	��q�_���$������r�>�'Mb�ö���KY�v�q�l������V�Xm�\:4��B悏*�����%��i=�l��'y�tsq�AC�5��KR�W)�;bV��L�)"��kq8b(��􁎬�e��P�Nj�Xmq|��Q��O�υ��I&ͱ�umB�'<Z�Ű��f¨|�T)D1���bQ��ѝ�V��{�"|����x�ɂ�D᳊+k׊B���%�go��ʜ�s����,D� �8���5�e��a�������e�<��RU�F1�%&Q��}`_���4�
̘��$���.ӏ��~-�#Z�ʢ���ن�ʿ|�x��d�;�����b"��u��z4u��WPO{	��+]�Q6�7+z~Cf2X��%I�BW�5п�w�H9}��Y���8`�/�BH�Ι��Q��I\e&W��流�Q~� ǲ&2����|pFՖ`�oZ��A�\���4�������iQ�D\����(*���d��L+���*����5�-���<5l�#�^�}��F�-��$!�w���N��̸���)j�lz��-ş`�����6ƿ�j�y/�2����M��g)i�K'@'��t9f�6�I'G?[MB��GF��ëT����@a:`�$5��A�K߉�z���I�<��>�d��'Cx*� "h]�����2uOe����#CJ6Q���r�r���6Z���R����+��>4��l�[��S�������V��$��h�;$S��?q��0�n������a�u��q�Z<� �T8e�[�*^�O�o��ӮTj
3�wS�Z�B�WQ��_W9r{;�)�֐��h��n��K��*YL��k�����_nN<��RH��� oTb'�_K蹫т:������b�94A4@#�k��p����F�|��S�;~V��^a�(��I����>����?V����c#}X49�%T�b!�|���#6!��e����C�g(2 ��8��)���l�2�J7��m��,M�L�5ݍ���]��������1�h�E�]UX��h��r�q��y%3�	�ܲNǱ�)���{�r�kv
)s��%��e3h�6�He�qsށ��O�WW�T.��uG	Y�U�͇l��<e��.��k�զ���O>�
�b�#�)KO� ]m>۞��
"
q��� �NFMV.g7������Ǌ����l]ĺ�lC��o;�I�Mny�S�[�F�Aa���#j�l��P�O��!���9K��q����w�ƬzmĢ��ߌ�c:�0>�vw���*T(�.4���9:�w�`NǞ�ID�� HD6�@�
���A���Y���ek�<�&Sm)��p�)T�I��i,7��zI[a�Hhjo�ڕ�ܡ����J�<��S��h֗��0~~Ky��b/b��U�	.V-?�$lpD�Fcr�Цd�c�~~*ܹV4��R����[}6T�Y��$�u�w���n��t"��bk��y]\�˚���OPS�kA_	�P���P͸d�09:����5h���ق�W԰�D�M���P�n�Y���h�q�oU�V���2Ն3� j��8	�-�
��鞢��@/�hk}Yo:39����$��c�<�g�t�N��M������6�
`eN���_R�M)���Vnr���]���,��ql��,b�R`I{���/�]$�_��-+�h_��pV�uȗ���N�,��K��.f%�Ŭj����uȐ0�?��lmX
T���J��Y��ɖ�f�*ӈ�@�Iؒ�w��`���������A�D�� ;����z�h����+���aH%v�?8U��G[����M���S=N�Z�sH�;ք��8�K%
- E��P�N�V���I��(�'�@��&z+�� ��䨯��ζ���7u}�0�E�}��k̻A?�� aߌ-��f� �P��6e�ǵ[��4�?:E���5~��F�Į�su�ĵ�ff���rG���4ذ��8�i�����h�5���7��qc����5 #y�5��«Ӡt�o���,bѧP��f}��Kp5�p���-lC���±�6��wg.*�����\�ӷL�d
�ҁ�̓����c.1��	�\�+�x���$VҖ��5�����|S��U��n������,�K/}��������.��nX���@9s�3�k8Fr� 5����k>�4���K� �t6+Q��>d;A1Ht�2[F��8?�yA����wZ�!�e.'/�i�PwZh)]L'�U*��	^H������حǃ���Q�栯�(u99j�c��CL`蓿<3��y#���߳r�ޟ�K�]��#��L�3�Y����GYA��Σ/],0��+�=,�6�"�ɭ%'�HQ����Q��h�@��*�:�@���o̯EЏ���h���~�qY/θ��v`��t��\^,Ǘ-����X�l�T!V�+q�p�Ӧo{��āŕ28��ts�,� �m ��Z?��"%�q&��<�lYKjoņ�&w�����X�,34�l�Rs�l�+�ɋ���Ē�Bs�}��V�"�e�%�øu���	
#*��*{�s]|��r"FAW��jx`p���bwο�����"�D��&D�K�1��R&�dHfZ�p�qYcF=Iw�K����;|%�a;��c�˭Z�gS�T�D=���/~�$|Q�)�}�k}���V����^�w���gE�t���kYa��;�\�~�U���U��hT������l��Hx��
v��u��v��$�|����9^灇/5&f���~xpw��#���1g�.-��&��xd�v�?}��a��F�E�;��]�$W�!��G����J�Y5���XO6ͮke�,WX��y���mֹ?*�ݪ��& H��My�m�o5?7S$��q�lV���8��o��U
���n(�'��v��=����%l���Ǖx��k������Db{h�ۣI{#��+�i�!�jj�ޓsi�� ?��+����:5J6m��a��p�����ײ� ���m����쪓�0����2�b�)���7��Mf��_��`�����{bvy;M6+C7,4����'����Ѩ�Ľ��cp�n�K�FJxZv�p���>�p��-"�9���e;�;X۞C�>��%�k��[�$�����n�|��I-L�@MٖdɷU�O�u"ehvf��V#&�MO���@�g�U*��A����,p�k8�4�@|���cb8Q�3
��m��0fW��/�U�e�:=�N�3"��z��װ��Q���e���d�GH	p9/��:K/�Y/��h��1k�.ӀP�������4�!�w���D�i�ʠ	�O�pʜܰ�с��� AY��·���^I��T	h&�)��\�(prz��i�w&���X�\{+Q���!j��*W����3a6��Ua�?�EF^2䴲
הėU_�Ē��7�K,@�5��ګ��]ཾ��G�Xɇ���c�*d��ua�dub+�g<G��!E2�-I25��w���I�i]�!j�F����$ŵ��A�Au�u4NW��V����`UL����W`שMнD��=�5к�OET����h�Ma���E9ȏ
2���`������f=�d�q؏)$���z��#^6�ͥ;I?�=�;&�.���e	ȼK�ј���;k�5���Vc����V�$��߶Y ���f!?C�~F꘾�  ��!�#$G��'��]��ky�.j����ަ0p�ʩw��޲P<�fgg�ǧҰ��E3�˗�Bk!�hC�K��_��+Y�kS�7߬�d^837�+�Ns�Z���+�U�B�� �s(�U���p��`�B\�oVB9O�`���ӺM�\<TQ>�q03�L��%��"#C,A�M�ik������<ѳ��XG�clm�[�}Ӈ�����RHo�/L�E���78I�
�-:��j��,2o?�G�p��K���c���tY�d�PN�@��?��-��_[f�LP}ɰ�;%8k*�n;�jN�!����� �A?p��s�D�d�D�.�C��N�)����c��nxNZ��������Y(Xlн��t��*����V�v�
��N�iZ\��D�-��$����*�w�{!%�2��=ψ���I,E;Lhէ=��A�/�����x���#u���%:\[y^�����R�e�(��%�lD����BͲ.�R֛�Jm����<�T���~����V��+�c�U1񃥉����T���8�ٙnw۠;d�D�n��{J�����bԀg�Vf���uA�m-Z�ن���O��7�K���fh�ȕ^�ﲫ�� 9ӤE�:�=�b>t�Z�l�l=@��Lx�u#Lm{q�u��'{|B O��D`R�r�b-r��1����ʦ��&�+�~��a�U�����\�]���@N�:L��g;��P����������廄@��Hz�l���ޭ81����$���[�-�Y���v�8������&��Ђ����*Ђ�Z?��������O�Y�"��)H�<���	L�k�ҋ~8 �d���>���"[|:R�»��=M����~ơ�C�<�6b��B*9n�m*�s8�5�c�n�jKb���no?�3�߶y3�z�N��\v	5��z����D�X���NR�=��A��%F{X~� ���;�|�6\�5"� N�Kjd��'�X�%�v{)NwШ!���E�v��\�z�%���lȊ�N��y�O=�hR��91]���)g�'���5�r�p��_�rX���c����P#��Qu��L._֌˨� �B�6�͊<�3����-��Z�Bə����gi[J�3+8ڳdX�R�;�igcI3�n���+!Ԡ�;K���5!�`6wW�M+nwGA��)!�+9�I �2΀��6��1%�I|����j`��b��8�a�5�# .]J�ZnB�'��!��4��j&M3d9��� �Bp�%@��K=�G� y_�K4���P��nK��6Xۻ�w�e[�4Y����s��y'J�cg�|v�蓿m�b��\��fC��F��d"�r��Y�lZj@��DJ�`��, �r��g�Ya���6G���*{��/��>���`v��)^ޢ����=eݻ�2��ʓ�v����>j���iDU�]��������>-��-�<��3zQԊ+(>>0�����2&ۮt8_�s�#�"�r/;��96F�����S��֗7!�	�{���b���ucΐ�f��}�2ń�8�3�F�}4��
������&u���$����`v���I �o� ���L<A9Φ�9c	�����{ê��v0s3����@<�u���m��q<�(-6~	t�v��D�3K��߻f�`���I�ـ_XwP�i�ɹҗ����U"KwTv�K��.��^�fT5v�:��av�{f�Wgo1r�R�@�?��E�R6��p����.Ū�O�)�;�8M�#�n��cܓ�x5t���A��
q. �K��D��9U�7r^P�0}~ˉ�t�N&d�L���N�݉iޫy+�W�,�Ł�9e�K���:�+����cT�1�����el�������,u:z��A�'P�J1A�WoE�#��T8ߖ���\�
�GQ� �L]��l�w��Ol�0�۪�V��;��҉̩7�b
�V����s=�->�#�%�+��"«��9�,t�o��JA����x���|u�����J���Ψ��Y�@��Y�&��/mN��a��v���A�;*o����󋠶�x�p��U[:�����h�t�h q����B4��"=��4��{��� /ֲi"0��z1-��5��)���(P�V&b�0�NjPGt��l�[N���ǩ�$�UFnف�2=��%y ;=�Co9xn�m��$��&+ ��KV�Ti��~����-6�`a8ˑ�9b��L�p|Tj�{�>"ی�:D)�SM��<��a�nv�jr:pV�L�l^�f;���4���ĵȤn��}�:�';��R��ߚK3�y�{R;���q�]C[/֢�:�RI�&(,�����-�d�Q�)HV	V�WP�:�3�=mx��S4�k�uR�آ�C�c8���e��ŵY:0�h���ГBs�iԈ��`�u~�1�~CI�P��1�K�$�O+o��-�j�W���>e���s��n�|Um��V�L�
x�F̼U05-և[?U)�ɩHj�����=�y����8�D)ӹ�~�Ӿ[�_�V�M��/��D����g�ЊD�[��dx�IFt}�|���=p^cB��R��Z�pj�:�XNz� m��[�3oq� �Bv�є���Q�0�!��YD��s�J���c�a�_8���n�2�W�n�k�N�@�F��+8��J�]��c�$5���uVÞ ��z��,-$0s�u� w�J�{걥
�r��E���M�'���$߃N6oZ�Y���z�[C��iUf���	����/4�vI�"�Ju���ȼ[?N���<"�HRs���o	�K=����щP$j�����PFe��?��2\�\����>Ǆ�t��*�/:��`�%r�")T�ڃ�*:�6����JI�~��,K6�����a: p}�����-%/l��黒h")=���,���P�t2 
����x�
Ϣ��m~��\����}[U��+;�D��qǊrbr�[9"f�r��gң6ǥ$�wEU�qt��-f�����}�At/GʔxW��$%ie��y�9�٤gI-�\�0������;���M�|ħF�]�WX�Q�lP�r>S�!��u�Q�����§�t?:�^)�hE�"̟��B0(m��?;��2ia�.�D}��D!��P&3�Z����L!��%h�b�(����ՙ�Х��@8�:s-'ĭ�;�JT�C��Xvi#h�Ǫ���Γ�ѓ�?w f�*?pY��`z��e�$(tǌz�q�Ħd(�$�>�ba���9����@L����0�O���]G����\��rWfDt1�uߪ�
5Nz�Q�����aV��c���o	�$��P�o5���MJg@a,��>���B;]n��^�$f�&�*�Z^n�*���Zँ�~/6���h�P*�?\�+�� �P@��~+R��ZC]O/p�C9��v;+Lu��6���5<���c��@}Weܙ?��gӎ��Lw��$2g�$
_�����O\��o���hl�٪��d�zc��()�dQɯA���Sf��^W#%D}�����,���rR��T��ȿkk��D�*oU�-�9�l7Vៀ ���-RF�
�e�k�P96Xmti�&ă��dD� ��+;��DՒ�Y������C��>څ�~����w%�tFB8�� ���=�+n���e�| �@g���+���Q�(R��걔3f��>���	�%��������rO%W��mia�Q)8����uQ[#J��7|-V�@}jf�To-&r�O�#��^ͽ;H4)�oLK�X�ĸ�������M�*]L'P'+.��>�Ye�I4P����<�f�H�$x(�e�G
2E6K&��mF��YOҜ_�Elj!�������G�?1�(��@cڏj�/i�ZV�w$�F%u�Z�c�
=H��!b�����&�mh�}*��?׎6���7N�i������וv����~D�T��j@�. ���z�;K��-@ӂ�>��]5���,�I|d�����A	�Q����I����rI�]�S�"]�z�?�p��6u\���їY��X�H�t�+w�[���/�l�k�DT ��Ta^>'���L&��V��v��fRZ�8{K��/�oB��ץ��]�i���L8:�Zibiav:�OɅ�.��^r����Y�kH/����� k��2������&��gn���Ia���=�ԵQE�7�}�7f�F%�E�8�mʦ��;�`D�G���=�&o�m�9$j8K/�	h�*nM�-�ܺ��`�D"}���*���yaV�y~�a�Χ�,b`����)�|Z�=�Ӹ���w�/LϣA)�a�L���V�.S/���ϒTr�9xJ'ȱ�](�����.\�����7���?�*����)xP�'��B�^=�;eAs�����{�j�F�u��%�4벥��'�o*l��,j(FD�M��o�M�����c�+�9�鿥���/!��_���7��
����]���M�iop�������8|�{^�l�t�%��⬷87���S�GbM�0a�R��CL��A�hypy-�F��{:��a�g�#
��ͤȼQ�~���
a���Ň�RZ�I8�M?#���f)���<Y�`\�\�(�~�q�}�P�,��Qe�M���=B�ir��}|�l�t�j�~%��X�h�s�d�&��!ͬ i&���BF'#Hg�i�H~-n7�+���ѣ�����U��ě_Ls��{7��@�@�`M�-n�1?Y9��헧x@�N8�'�b���e&_,�+��W+t�a�Д�yF(�=�"I"p�:�``�A`��������AE��y��va������v�~Fm��+���\I�ӧ�u�1�r�y�r�2�e�m �����b�N�.�R�&"���Q4�[?9�ǜ�`.upɗ��Y	��ۭ�̄�����"z�΍�6����>T�s���vኦ�Z��6�#����Qd�~p�ͮP�?\|9u3ڝBcGU$'7h�W&.xVB���`���0�J������+��5ω�"3cGe�&���W�vC2�	�n72�܃�|�e���}���Qq����p��@9���>��Ev�8�5M�u	��Y���,����K�ŉ!��.�*�V��Oq�"?�,��8�`�>Ą��~E��nm�3=�U?D��_���7���j2�U�����������j�pQ�����{3�Lrﻜ��lÃ��K� �]�vS9)V�!�a�.�驋��Dʢ�����8��9"�g�y��~Mb(����7���KTc_��<�Ֆ+^�@L�$e%�1��߮L)S���-z^� ƿ"��cA-���b�4���- �\Et�T�j��|�^��bXl.�b60��͂��<2TYT��WJZ������^V���O\�0���,��H�:�?���[�Čn��f�+A�@���v�"7�K��|Lr	�я����r���IPHT��-������P������T�aT,t���-
Ѥo�b��Y����R�:�w^���."��-.��4P�[�,���XTQ�C�W �\!���^R�U�Or���Dh���^�W�������<� � �y���>^ȃ��Ob��Ef�A��\Z3�(z�gV|7\�4� �,X��[��L6��{�D�Y`�����wլ���Gz5�%���"��Y��<Y��\�	�R���?D��1���0��x_�T��+D������J_di�c���	���&������2L��dD�s�eʺXgA�	�|�wړ�p�%V�M�+�2_��"h	��@=���;�,Sf�����QZ��?���J$�9� �
�{.���J�%�#bBP��~v��[�|�G��c祎edf�M�-ۊ�Ըq�4
�4}+��ϖA{�]�!�\��)��"����hs�"_�C3|�}|�I3_��s�pF�����%�8�W4EU��q"G���05�Ï�r]��4���տ���v��hq�E�����v��uf2�3���	���X���"g�]@J^�\���v���E�U+��j�f`%C��P{�ݹ��ȵF��s�^"�m�'�f`�z���ɚ��W�9�IkH�o4{,��g/�*�^���&,�8�U;x4�Y��t��zzgh*�����9��H��u'd�%�]��f܍y�C�j<g�m>��$��z��&j��G&-'i��6<�b9��1�[��oA0Ԫ��t5F�����%U�X�]�Epv�+��%>�]���K�V�ѯD�&E�)zD�����3N6.a�u&�iQ�,�L�.0����Mm�-%Çd��K�D�����MVz�G�:�c��`��l��B'a�LW_��j^e﫡�nȡ W߉[z9a�0^"����X3ć��xYc��+
��gB���/["o�M��y��k������D�) ����:L'ʈp7*���%��(�N:���ϥ6��;�૝s�����.R����F��C�΁ΫD�����0��_�ۆ�V���W*FӬ�Q󩋤������%��E4��4���ԗ8��4����o�mrqJBޮn�h�]���$��Fe�t����[E���h,=�$M��4����0�H�ڃ��a�Uao�7�n7�������N��<��[c�}�	'�~q����`y]�\�'��D$'38BSz�q��O��D`2��0/yI
�i3��g$�2�3���aq�mB�/��o�0J�p��J�>�tak��[��%|&��֫\v!V;&�;<�B�`Ҧ��ĘB�K��R ���Aq��r�x��m�E}�w��]�{ȳ(֧	�D��x-��/{,��0d J�|�K&y��D��������7�/�ٝ�����U ���hf�W�����o�xB�E�S9�׺���k �8O�Tn��1��t�8��b��8D����}9�م�\�ы��16��H�2u�#s�p<�d�_+��Oܓߝ�R��Ly�
,�Ѵ��A,˓��<�7�)�ű硷o���Q�a�H�׋G�zM"�8(�"�h��_�6�ހ�����{.�	��ʻ
�k<��G�:���Zp���(m�+�gw��wd��{�����Z�R
/��E%$2���2�T2�D�"o;�����C�o�/)iՉ�nϼ�����q�n�m��Bn��6#���~y�X k�.���\���$H�9��*i����@�0���G�c����Ή�Utw<dS���U:�T*��Z,��s���f�"t��7D0a�p�+��1A�#�I�e@p"p?�U�/�U��i��.��8O0�9���ޥ�9y�\W�cKq|�>�W��vT;wz�%>h������D�B ���P��PEb:V�H������5�g��%E�U���ֿ2L�`sc%;d8����><5���|�)�8Qc
9�|�.��V31���6���h���N�n�Q&3x+�ǥ�  ���(@��7������װf#�mBK�Y��\������Yh59�6%�����W7>�w�o�EIѢ_�P�߶�ݠ*[��v�>�N�L,�'G&Cgl2��k�;m�Aoz�|���l��r+!ȶ[��z��o�5�n���Tk��xւ���:5�����F;{͞S�����T���YLtWK��<�L�Nl��/��c=�1�K�nR��6}��<�o��������H۹$���Ir�g�?U�t^���`�?��Z��96j��·�2��T�+�30�˰�w䉙�r�A򟺫���L[�ز.�z[�U��Ϲ #�q*��F���F=�Qt~�g����XOi�=���k}uc���׃��:�U����{�5.C�d��y(�_)]j��z~%�Z��bu渫�f��|e��	�0ӟ _�P��o����W��8REΐ!x2�!�jd��v6n{�?�K&�Bc��	�ME�ͬ���=hL=A�d��,6M�Hm��_ݜ2�f+-��pv�C���*y�'��+��f�6�P>�����?l�*	l��*�#J�6�g�e�yb&)��D V1[��^:<&�X�S��f���[R��[G���K�E�1���PE庴�u�9w���pLR��f�v�c���!�[\�ͷ��,|��y��0�:�y��Z���'����<l(���0�	���Zj�wbE�H�@�nr�Y3�@�
<�Wm/}�K�j�(����3�g��OW
N�����q jxD:ug�~���Z���	��k�rD��t�ZW.�v~�+�^�-.�=�0X�kFwYgAV�jc���{a�~I�2��v.3�l�ȧP�#�T�37��{��
U�'�ii��$��Z���H��������;�>�"Ը�0�>[]{���W��(dS=�����uy	8
hx���i�uj�!����j�u|���(r7��E��O��qZ+Sϲ"eR���!�(A(���������I^�%/�(���ymSv��
.��s�!A���_��D�>7�9[woe2�T&�j��+��?�2�Ċ����^J��X�*��-��be|g!�i�~�R��o�$��N���Ne�!��T�փ����{a������K]�4~^D[�/s����O:[?B�eu7:������Zx?�$j��sU�2T0���&-�C���W޵����:~�QI��a��b�q��	�)6F�(k���Hj��v��D��]����h'�ؘ�p��K���Z|�I��Zg����}�ކ!D�x\�.PA�����PWϢ]�E��1�*}�NъMVy5�q���
2P.��Yޛ+U����v�઒�7]�
$ё���&�\���d�-/�3hUd���;�q;|W��ɩ5�,�l��jcb�Bz|y���'�4����\��n.{=�s������ bQ�G�GDX+��#�Ld{�Ln�?�w�9���ngaW���R����7��NJ'5=�&��P����I��TH���Y�+�������9�I�ې�42�N�&�a��6����Re
�����-	=	*j�Z����:3A0{�2{��\����B�����d�T��r�"��jB�o�a:qim�=G�r%�"���p�Ap������Ll� 뀦�����Y�x�������Q����3�d>|D� ��Su�c�h~��a��r~�u�[xv���݃�Ȯ�62��мD扪�w�|&�?e�Q�;��n��n�כ��ek߿~����?��پ^����6�����V��EC��r�����S�G��� ��|i�����K:� ��kW��}8zB��# �$Ц<R��65�z	1a�h�~���R���<��&����L=�jyz�O��V��b[��*/�����'=vA	���u���J�
�����M�N#op��l
��A�eL�O�����E��p0&��.̔
YB4M��ǃ2�ژ�q�v7���@�ػ�sZ/��������Ɔp��> 򭂝��XRK��U�T/F�%cI�b����) @�j���<q�\���ǼE����a���ї��e�0o<˒�R6�9��Sѧ�U�e߆sz�z�5g
40�R�ip�WF�����%y��yoЊc�Լz"D��d(5�?��!�_o8n�r�}�r��M�X����6W�E������_u3���Z�¢{�tF"��n1�S#�ս���-�N��O�^�������V�͜v �*���ZI\,"�(�SQW�
eٰ��fH���RF�2@n>Wܘp�x�^k����)�(#��s�>_� ��d�)D*� 6���R H�D)�	V�i�*�Z��7�pU��)*���~P�!-�l��+�����_�ƾ4�u՟ʵݭ�7�3��6Ʒ��s���Ts�F�����B�"�ޕ��+.���=�S>4��A}�GmB�=�惼 �I��`e�\s �:p��Jɦx�����\^����.�@R?+[^꘼
�%%��Xu=d����W�>�S.
(���������2���y�Xؗ����;b�� ���n~��ӯ�Nٺb�E	���OYG<�#B���o^��E�5X�j3X��V��A�XR��)+���!?v3�d���eמ��w̞)��S�O���va�Y�@h��-j� ��M_�֜2j�ݼ �k|KH�9�P��9���-�֙�V�bY�ڑ(7��.vϊ^���������U�Jrn��W��;=4�JXg��a��H���e�2\�1�+s
F��v����
 �I���7��m�ڴ�܇�Ċ�8���Ӝ?�"�t�}zj��P	r���\�<�$lfE(.+���$pj�g��J��2`��<^����^ -Ӛ"@\�x~��#�#���� ��$��v�RD5uS��N�15$��w��S�Pd8��Mn�*�8Z�Z�=�#�0��m��4�f¯�%�X�釱FUH.b�!�:x���EPN����yi_���L�"��/��&UI�{��mj]ɡ����D�R�u�T�˛dhszjv�iJ=��Es�B��%W�����4aY����%���jΆ3���7=�ԕ0�l��Ǯ{Xzg�
��򿩕i�C�t�Մe����ׇD��YP�H�-�.�'A�;�^<�+�J
:�k��~b̡�7�)Y�N�D�ǘ��i�@�����Gl�F�R�zU���=%O���RqS/��Ld;l��t*SA�	��	��56�盰����;�<TŅZ�M�s�R���U�3}1H^�`~7�1�3��$��+�
j��r@)#� z��Q�b�`d1�|x��� C��
f����xqr���,N*����>�A���97�@ޘS��|����4�^��9��wq�)���C�҄��v�p�}{����Ր��0�d�����4TI���Ti1.����L��'+0+8:1��Y\���,����;'2�N�<��(*���"��]U{��Rܵ�8�x���j�W��CY�%���|k�����6%;�C��9C]E�$�.d`?����S��4��Ipʭr�%�x击s�,1�@u9�l���BcJ�8Ig�c�2���e���*b�!s%��S�[���?�j��aCz�0!+v�W"V��Y����V&ƪ���[�SQ{G[�\XJu�,0*�6�$���A-�X{yv.�NY���]>�~��6;
��@)l�>z���k��֜.�'�=�W���hD���f %���-����6�o���S t�U%?���HN�$��p�2�B��`�&�֪�p����Q�ʐڹ	�lG�-��C�kþ�!�e�Ĝ[�w��Q;,�#�hLME�5��ZN���u��	V���l�X�.�ih�ю�2E�J�/ǒW��[L���8��2�f�"s�V�r9w/S�]�(/{�as���R*����S�`$��K��C\n�B�n��"��F4��A5�
c+n#����^p2D�-0�P��Q������'ܮeΫ���K;p�����)�K����P��?(I����#��f�/��=�@�tw���nO�g66���.շ��#�2jSn��V�K�KR ���%�y�Ӟ
�xJW���`J�xhr/���|�o,z����[]I��Qc$'����+�Z?���t�������ÍU���-ǘ~���A�����$�e���.qf��w�*F�<��#�d��z!���2,�)F6��|�L{��=lZ��}���� i]} �q��8<Y�l�'�kz�g�+(���:�7�c�������r3C��^Q��|�T)�/7�Vn~��ɿ��8W���m@��P��G:�0��#��^��=껾����xM��Hb�#,B�� M�e�eG`��94��`�WޝD5��U��I"ul���>U ��v(o�a�V�t+�ݿ]�F��P��8c�/�����C3��*��w�h^�r5ϻ{����9��X�p8oU��S]a
8��:"�6��W��u&4�,�1'��3ZU�Lk��C�Q3o qcb�����fԘ���.�z������D�4eK�n r3X�" ��a�OO���"��	���'���J=��|��
��q:��h��n��eQ�r�Ʉv;�p!��A �7T�oTQ?��K!�����Z��� �o{���O�z���h�z6�0Ĝ�T������T��z��!�-���A�ot(���^i���9���Xp�󋁥�W�E�"�V�S8h�����H^j��Rƒ�('�*8�Je�B���0 z������Q�||��z��|+��?-���}���/PF��2�k�ߢ�TO��ƐqV����f��^r3�Q�!��`���|/�Y�u�c���k�� �j�{��Ѿ�F��\�1�5x�Y�{Z�!�y�����o�d�%��y��^(e�w��	C*���#݄Z{x�g��)���Y����Ɠӂ	�R��
{%e+e2��;�tZ��%����`�I���&f;�38��w?�!~�#9���N�o/�Z��WU`k]��1�y9�����?'zr�fj�b�x�A�}q�ky��l��&]�o�o�������vB�΢���	��䷙�|L�>��6��}׫���2���r[���٤qJ�}��ݣ�bM�fa�P�	���:o���x���ɼ�=�w�C�7�8
^����q���Q��$��2s��%S�o"D���5z��+)�3�����>,�@�%�nٸf����.�;��$��6�N	����X�H0$�	�i�Q��qIu�6�AY�i?����n�)DG�'��Nph!~Z�/KY�^L�,)��lw�(B{s�:��.6����/���bi\͟���Q�&^�L���$��HLQv7�mk�蔑�.�#=�sK/�߉��5oՖUm��m|&O;�K�B=�h�#*��.���/4��y�'���M�е�BL�o��X��D��HlD@	-�5������*����N߳>�M)��/��vj��65��nAl�r�7��NݽB���T-³qXq�)
�b���7��[���u��Z1�',� O�NJ���7"����y<�|w�KW�vD|�݌��5:�W��.��y����hZ�c^ �~b��@R��C`�>�:�������$������$����~:��<i��B�X{#��<^��hL\&V����Yu�.��)��FI-9������-��,YgM���ݸgX�yS�}9{�q���OTഠ���Ւ�"^7eTȕG�w� o�D��8����c�Re7P=��"�x=��F�Φ�D�M	�K��G�y�B�c�t�YEÏ�(LY��x`�
�����[v z������Fha�O['�}'&�����C���'�A�(�m�v�=�-jR9�Ԥ4~�5b%觾	�.�4zι%��{j�%�t1!�У��|
�_�����RT:>8w��(+,1kT��V6S�����b8� �{�¦J����Cd^t�'�����t���/(���R����`kK`������	R��1����r��b<+��H-�&���C�J���x>�="�ánV�miu�@�4a�����	����"��aIì��L��|�׾BT�9�d�Z9�Y���&��p�ѩPD躒�9�h��0��odiL�\�V���+�����:Fa������pi>��\�u�9�N��?'9,�#�t���,�t����79U3���?���]���e+����oU^Cr/����1��=��Z����q��$/����e�Ev�Sݏ�DiD\�8����rJ�#_6ON��;��,�����.����56�<#��S��Y��[���%��������;�jaH�uI�����y��Şп7˪'���o�B��,��r�(xp���"�)�
hiM�&��F�z�{�����*7�R����tRp�E��<7U�tdu_=�8�Ⱦ�@د��c�"ϋ�����a|�O�nX���܍�Ui��b[D0E���_����,���j!J�EP���.g����*����<���Bl�KVo�t���)7�%r��p���[���C\��q�B�n����: ��j #*ߟ��U?ha]!���NS~�.^��R��j�6��a�J���͋TP��/��{�`.�-����z=�f��LF?S�2N"	=�]/�r٥�N�:����L����5�]�i��w@v�Unv}��CQ�R)��|�PX��;&OQE u���%7�Z�v�Ї56u� �q��;7�ͧG���U)? ����A��y6f�h[5�<aÀ���?8�!ԚP�8r?��\m�sf��o���jnE*�݇��H�9 ��#
n\�J=X���M��)�jz��A�Ɩb����>��8��H��:���#��.XG�2�� [U�\����=���xO��C�^;�s�)a�ُ2���±A�_�X�&�\�#�4۲��rxK�W����IM��y�o�J*fT����l���K�'�.���FG$�=��B~����_�%�sF�9� �ʶJ?��s!?���~5rߤ�� {�ZW3ڲ�b>�ζ֍�'@�&���J�q��􅿪��<����u�9�j�6�2�ʥ�O���%�N>������1��z�=�/���)IQ�}������C&�����~��� WAX�-��	���d�UMz���"�F�	.N>#���7X��P2�[��D�ټ=��q�C2mG K�c��̟��f�Ah���t��an�����!Uu�&/�T��w�D$�R%����ͣnM8��+��5_K��
�I��kѪD�MI�t��o%%�����
���c�M�$d�b��\�"jQ�!j�qGn^х3�ex��#b%�9i�����%�}{AX���+NxH�Mj�-T�C<�X"�vW����Ȕ �BR�[���k_����ɋmGK	��m�+��)�^@��-b����G(���pu�C�A`q�f���D����@���)Bsu��0]1fC�"�}"g���tUg�\&I
��-�D����#L�%�7��[`>!.�(�`I�^Yz*m���|J3
�!!��M�N��-T3��x��]�lI4���2%?��gm4@C����Ǌ����]ռ�y%��]m�� ��*^`X�
H���R¼�EY6��5Y��PĒ�����ʘO�y��ID��|�+�j��N�ߍ�H�^���q;v����|�/7�K(nB�a����O���o+�1]���堳ܓҙ��lMTN;q�\�%{CP��,��H����u�<��T�,`u���E��b�~h��繲[t=��5��fb��Β%sg�.Ua��CR�����L�"j-x����R�V{���?��:��~W!��U��ˍD6�m��e�B5�	�k}p�',H�
�<>�8�x�Aڵ�f�	ℜ�T(C�|���~�C=]�@�g��&���+�e�E#>JHu<��Ru+�x|f8ُ�.k�G�YI������͕,��2�~��J�����&���ju���s'�w����ȧM�j+.Z�{,ǟ� ٹ-u_ U����WR����� �*'���Jce+�	��?)q�Js��lB��#v�r�=�GW��A&����NL�Tt�R���t�"�0afO��g�e���hP/�0�L�0�\:���ji����&B�^c���O\��Zɰ=�^=�ґ`����ltɇ��i�]�1��!���K�Fy�2��r��Q�����+T׈����W��R�|�����K�d�G�nQ~��M��V��X﯊:6R�F��/[�PI�w��7v�S\G�����5r1Ӑ�ʅwB��EbVr�y��'�ᐬ��)����d�]���^H�Y���ŕ�⺍<'Ҟ{�5��_-��]g>�{`�Ei�q����4Tw;<J[Db�5��$"mL*�І��]����L���r�^J|��,��c�_Z#��Q�x�A/Ti��3����,%�r�0ޑ�p�$�GW����^���0��H�A!������lԀ}jv�qQ�>ֽ3��_�N�|o���F�KG�Y�Ѿs��V��<�P��&����X�0�(Ug)�K��k�ҹ���������H&	�����Y[O|L�Ф��I� X��r6�N3��ds�5M򷣌�$�6��^u3�j�l��1��^�Ru*dウ�2aG���Yc|���ǈ /��8��}&�Ǜ���Ƕy��Y��5*�7����N
-��ĺd}z��,��"�(���y�������J3����#x�6�rN��J/�bWy��\d߈��H�4�!F�j.��MQN�7�G�̭W�Uq qW��$�����1q_���^��r�fW_m���!h_����Rv�i��H􉰐�;�Km��{������$Vf�ۑB��4�Bpm�
䨻b�����3����S\�ڼ��i���i�W-R���H�uU>�Hȸ}��	x��S�.��*6����@S��(�_�����ϸL|љ�8Jƴ8����@�!Z�?�=��<��CHmy�,�028bSE��̻;B�w�@d�P̪W(�Üm��8?�ϮQu�)��	������\ b�Y�o�	��W���0�eھJ����
�W��Z�'_G��ȱ_6D�r����E�ǆ���7��^j��Ԅ�Z�y)�9����F�`��2b;�N�� _Ї��d��_V�:�#I�'��k��Q�벇�ch��h�Zu5b�jE2[ǏG4j��G*���G%�A�e2�y-ξl�(5_�s�.�9��3銒�#�:j�Ϳv��w7	�����䩯ɅZ���fJB�A�֒��W�����|��*H)��Q3�6ӳ� �`?����4�����Oi�Ss��b�)拹`R�s
U��W�P'�0�U)�D�ȡ�z��g�" �k]Ѫ�@ђk|�GD�%������Oc�X���\O]���}��3�--�mB-�Bǧ�������Y�+�^���m�����KM&`���������Q)xϓz;�C1�N$���ɌAx�]��p�?��hD,�Y��џ�)��􍴐H?�3ұ�j�u5���jj��K��2ޓ�C��������ԡډ�G�_��T�MJ\����b�,u[���U�������vw�o�1��yW�~tH�/��_�n�i�uA�|ļ��.A�����<��ؐy�EJ�ѕ(��/ ��j������vy�\��=���`�@͙ne��ϵ��������A���4n�e�f~���?�̇Eb'�ꤿ�B���8��7��dV��ҫ�b�<������ð���D͋Pu�89
�w�oA:ex�%B!q���Z8Jo�(�7"�Pj���*������
z@��ܷG(dk�,2��JK���~��_�쯣+
S�PZ�},��}[��qv�A]�N{��U���:��l-K�e�C��V��&D�G��$ڄ���]X�6ۅ�? ��eT�U�r6MI�u�Q z�7a���D����W�Pe �N�OV��)��CV˃G$?�ҳ�����Z����>\�L6�6�cFa�K�1�pLr�e��^iMU�9�%�������f�?� �l����uF?���b��5?w�/�NH�uJ�VKuĽ�]i���b�����'٬���0�Y����3rA�����[L(�`/;(3뒗��Ǥb�ǔ���:��`Q+[A/�����J����O�� y:���g��^��f�k�XgN�q��Kc�h�B�޺�t;�������cKq��{\��0�_��Ug�y�3\S7�~�w�v����� R�����ư٥wϬ~p_�r�����̃vt
ܩ�!Ζ62٫1�E��Ib�p�2_�t	ҿ �F��7&W[0�5p��~my\��m�Q5�fS!���V&=6��あ<�j�[G{$v2i���<��A5�I�_L���~���e��ř�^MK�p�g�:�����g����р��V�^_̷�'=@����=�M��n_'� 8r]R�&��lVU\=��H�pBnJ1GY�bw�>�
4��"�b�=>4�1򓻥������Ϥ��c���t��h���.L�@؆W
:{�� o�/�U��\������r�k�c��I�ډ�{6���"��!�"��P��>Ȏ�k�D�/����f�G�E�����?1վ�F`_c ��{�����1}��¤rPf
�l�Xm��wc.~���4o���>��V$��b��#U	H����uNu�՚�����
AVP�6!א!��v�=�@O�#�G�#����)g��u���a��T��b�W��g����؈y��v��mz��=��D(5'4�b�o���P����"ׅ���� 'j��
�m�R��F#>����f_��*���~�kFs��5e�-�"~�������qu&gVV�3�#g驊i�)����H�H�&߼\,��D�&'uU��B�z�/ֽ���(r�G �c��5g?ׅ/LeΌ����SŹO���=�7;��Ex���#�U:���t�+���m����D���>~��lz�o�Wԁ�mk���_�^u��Y�Z�O�Yf��7v�������븾,�K��
���������>��Cxɛ'�xŻ��i��;�K�B�fY��S2���u����������rLgj��l���RS�Qܦ�&�x~�im��,��Ͻ �D�6A�N&�iZi^6{����D�,I83�w2�Z.�}3��UzD�^�i��8D�*�ɭ�Ǜg�i��e[�N݌�x��nۏ�G����-����;}�EI�Q\�Hs�lalbYI�@q�<�	AYŘ�i�싣(&8ܡYF��u>��,>��L��j@��}M񹃻�AV:V��?u�#�/��hkSzr>�� {�u\(9�T�)�$i��̌N(n�jc���Jɪg7�"��;�Gs=�0>[�Jg���:#M!��"�����s���s�ww����W3K�l3� !FjL&(t�u��9w#�)Z��Mk ��p�&Fw�E�3ј18��x�sO��I0Z��BȾ�K��aF"��-���0@�-��w]�c�u7L�j�X��q(&R:���@��C�a;�l�M���7R`-����������jH�P$�*��V��=`��8��6vXJ#�t�u�j���z��.��ɟ���
����Φ�As���U�K̦�L�DRQ��5RU� ��� &<�:����R������dκ[�g$_xI�ht<F��!�B�6欖=�/�5�"o��i�?Ԭk�Xiy>�!�=<�=M]6_
��ǭ=5�RR�'�����V�Қ�S�BCO�4�>{8���% )믆jS�[���Z��]WТRMk�3�YU>��|�����Ε&`C�ͺ��h�ʋ�iyYA6]�^}&��u{֖��nce�T:�?,�F���*	:�8W�K3S��:��~V�r�y�"��v�����(� B�Y ,���'��ƽ�3Q��vTEH�Ը� yGL	��B�n4��L9��J� M�$^�����F��}A�l�SK�<��X�[��oh���a�[��"��O�[5	��X�+���������(8d�e���.}��~��^K��Z��r�!�`0bt�1ZwJk����OZ� ^����.9-�;���Ə��X�Ȕ�/ud�!<i\A_�g��J��Xyy6h@o�&D@�	�w����U���E�&X��ɑ��E���{�����x�r��~sN� �ޯ*�$�^�li��>��ˆ:	"�D����R	�ee�~I�ղ�y�(�gu��B�X*�ݷ|�6S�\/�+ɏ~��D>H�c���8xN�8�W|�S?JP�����-��0)�T4��\#�Z�@N��F�d�����rW�&���<|%b��<K��X���^:Bm�B�=���zt
�*x�`���a��̧���t��ԞZ��ۮBT�ވ��:�@p� X[Ƽ"T�¹�3u�A?�!�(�=y
�-G��\:j_5��@)G�Nm��ӓ����ޮ��&��*C�z��ސ�u����b&�������l�ϐ�,��X�w�2a2��<���6IB'���rz���˫N��=��֞�)-r��j���S���*ֶ��H��9i������aEǯ)��@�,ܐه�F��|Bt�q�a|�0}0�&!185~��[�S�Q�}b��̳�Ѹ
�(�1�׎�����N�NUy��w.젮�M�u�ؖ��2L}	�e�iUe��aB�90	��&� Uvq�кC=
��
������B�4_oS��2��gق�;��x׬8JDx�Cq�)B�~��͞$o <����C;���)7�o�N��4��l՞C^���U�@.��{��7���;>��,�"b�Ⱬ�{���`+X]��h���ө�k.�9~?AXQ�# U��C�U�{h�FZ_�,���5�}`�&�G��ʥ_{E���a�Ѡ�g{B��Al~%#��v�
[�ߑ��#u8�/��D��u��=v�3Z	�gz��0�'��c�r�1n�����hS���߯�L�Y�"K�ӷ��(^�Z3_%��}�hC8�+j�ͦ��I.���0Txd1$��8�����O����(�V�.��	8�^����n}!��^X�O�\4�kvI����},���Y�j����ٙ�
��9�F[&!�)3����OD1ň�7tЋ����d�����=Z�`�6Cr��f�>��AX�#	紳�ci#RжA�@˹�eݒ��Ӥ���'n!�b����`e�ǉ����}/�Z��>���a֪0:A�eܢ`��z.ye�
F��7�?�.�;k���"m�M��Ri�!��uT�.1�����(��g��o/!����j�h��$���T�sJ'{�ۮAe�ܰ8@{W=�����������/��x��͍m���Z8?�d�Cb��$mΡ�Y��T�S$�;����U����@����]���>iG޺�L�m-/y����:%o�4�JA�j ����2E1��yuV�C���Aq�X�a'쓚�=����S��[Nj��P���*�o��Z~���wv��d�i�D9�i��l�f�_���T�b!FvG�bZ��pvI}פՠ�E��m/�� �g�X	��?�ܷ��|����D���B�9{Mz�����в]����t����nx�N�fT�g �o��z�,;u��4s�սzl�1�"ݝ��`??�HF�{�P�2�t-z������k��.H�o&h쵲  3��w�b�y��x���z�B��.u>c�]�u�P����K����_�Ԩ�l�G��,�9/��Q�
�E����� "�	U��Nbݮ� Ok�]@7,udK'�c*[����v��)[֖g�O�J�?�u�N<Y<�<�l���\�'�=�vg�'?��Cx;%|�Θ�D�r??���P5�/AVS��6PM��ɮ�$eA�#i��%]X��KN��?;�c��Bw�	��ld�����l
����(�U��O4�u�Fn��6�٢oLE]�{2�����w�4��q8�$H����6���f��%�´�V�Y#"�Q?�"��Q��gPi5)F�<s��a�G5�7ã>g3������@�?f��� ʛ�shq�Q�]�JI��22�WF�T�,=�Ch
�sVL���n:C�X������?�Z��	c�,�6V"i�������΄q)m�C.'���@��4����q�c/��M��̕+�T�-s�k7�_��1p�� ���֗q<	��d7/ �\�(�L�O�����/ciP��$*D�O�˵��r����ɰ6%do�]a�6ʦ��N�Z�p0Wt:�Z$������ܔ{6\�_Q����9DP�̚&1@�����r�S����	��kAQ��ʂ��LF�r�K�([�r�0T�1.氢?�.t��Ve&�{��w��-�E�ʠj�MV����������x�[^h�bgK"�U0&�Fm�B1�N���iLj���Td�����w2��MyH�p��ԉ�Mt��!B��n�즇Uyi�]��!.��F��1%,��դ�` ��T�Jݼ��7�t�5yr�vIVO~I�����Ys�����ib���	�q!�:�p�(�٢-BL�p^��؁��8`����� {��%M5!��fGL?p�k��� �>���Ly,vJMxˇ���Ic��7�q�q3g�j����PHw~�� H�����D�H��ت�Y�u�0%-��%��_~�@��[�><��&�bnD%��=u�{b��Ko�O��>��:9}�����6@p紃�{�n�d������r�͏����0h"{���yHw�m� ��a]������S(��_,G�*�ԩd'�-���ayP�ԋ�n�X�Ā?����*�qH��Դ�_�4�N�q�X��&t�����=�)��VO�!���ć>�W���*1������r�;�C���LV����z$d;�Ɩ��4L'�����ӻ�U�LЗ���ݨ.��bIn���垕������{���P�����#n���9@�����g�Ķ�-<��wb���j���b |��Y����D����� �{��$0� �
~U������LZH��$���u�I�W�2����Y�o��&E`��_&�ꊻ�菡�-c�����sk���H����{Ӱ������/Ϗ+��J�ԖnԴ6�J�I�T,7��G5�*���QZ�eF�{��Tl)��+k��,X�=�ӑ�[>�I�v�1?g4�:u�q�T1�l�������ŏ�EPܥ���cY�O&:b=�}=��I��yN�3��"�M^vf3��o�]���e8��C�%�>��@@w.�;��e%qKK���!  ���W)�[h��ͯ������h���'�a�7���a&`'.��̴�?�*������)��b�&�X�������ԉھ���pzVK���I����\����<�t��Н7�ȩ��ٸ��"3�t�v:�����������mB/���D�]�'�~�z�ΚPi��<N|�p�/"c
il���Q�p"��vz���#�HFDө�jmBbg���H�F{�y�[ڙ�E���W��A�q�	H���i�VӖ�� !^�6���J�z��oVRI�il@*ҟ�j�~�R�+��ᇣ���yj0n��m8EC�� O���C�~�*������e-Y�)���D��b����hV��G?3N�%e���*}H
ۚV�-8�w>.��
R�`[%U��f����L�gH5p�W�qD�gb�Z���eE�JA&����c���1u(|=jb R/�;A�%.P�}�X�^����|�<n�ki*"�����/�́����
��ѓ��0 KMI�R���41��M�M�Y,`�B�l%�y^��� L�7.�z�f��n������x�')��D)����c0wN6)J����>���M�X�_�DW�~��7w ��,�7rk��'���-��@����~2�����>�+;��K��S�z����_�V(�_��w"���ܿ��5���'J��5j1��������zn�����	�gO�K����X�/�7���A��069G9_��:-}F�'��A��������hE�QF�M$7���Y_�?�ʰ~ʭM�� �YEȗ:�����2�.28Hv9���GM�ĳ� c� ��?)I~Wya,��cB�q\|�[Q]R�o^�|��	�ZP�y���9�����~��{��)��)ٽ��W��b1��LbxyWaיЉ�`�@ �������v�S�v��6���g=�S�0g7g��֐�0;�wx�y�_��j��5!�ٜ"U�ĝ�PVw$ͧq���t�k���&y��&�W�nb���X��d � ����+��m�����0�jx}���y�eU�PC4-�bl�`� )���<��Fp4�z'���b#�z����?�����=�Δ-�k9�fA�~�v'{�"or�&r9L�Y
��7I�z��U���B����ށ��䃖{�I&��FJC�>W7!$_$g�c�O)J!qds��Rˍ)��?����`��r��e�Ka!�	1�H3�_=	ݢ�i��_�X���q^�1�Tn��h�R:<{���|Щ/��A��Yƈ��bu�i���R�$v1�&Oޔ%DH�%V��ϕ�>j��;
�ʔ<98���ٛ������G�Xdl^ʋ�ͅ�����P&w�P��xś�T�9^|���Ѽ��/����p�6���sӯټ�|��=�V�T�9g{=��d����3�O�_�1�f�%��������l���� G����D�C��3K�g��c�� #�_��=G�#-u�p�aހ���a8�����ߛ{1z�^Y6_,�< @�7�	�����j�8�������ٍMt:�v� �g_����]���%�bU&A�f�/S�+po�V�3c��6��˕�f�:1����$\�"� T�0���'�[9�J�"�b'�
 T����xhA�>��K��������&mK}0�Hf�?kBaA�J�{Υ��M��I��wU�`�5�Drw�}*{T�`�ax��Ȳ�P���qyD���*����㐾|�U��+z4�n�i�e]K͗�P��S���\*�4��R��']�?��a2�ue�d��ϛx�{����M�kGbn����\)���,?��r��y�;VX���ǳ��D-X]����K"{e:� ���~{�U�z���VZ������}�������>���B�=w���;)��x��s�zx%Ns�����)c�������]ȴ�F� �U�u�w�G�!����Q:�,[�m@@#~�{E�G)��9����m4s��Wؽ����u(���^27KY����_�\
�-.��V���=_T�z}7f�b�X��JS��8h�ɫ̟�=��������Y[\;�ވ۝��t'1���1�<C����J���7~�ml*[��C�)��&�>"�ZϻY\'1�J!�1D(n���͝L��٨ ���s^��D~ ݴ�O�ueHZ����-��,��d�Wm��R}�n��c��$�M-�l�^&�r��"�m{����J��5���������P`�`q$��oʃ�>3d2E��'f	Q�u͔+f;���3b�$#��
�-k��,U�;����BҞvy �
3^=�f$�XYxg�s��h���ߦ�Y"	oYxړ|���Ȼ���y͐��q�K�����"��VzO�ٞ�$���$Hm:�fN!A�""|�����v��
s9dj�\�犆9��47]Z�o���KB�p��"��=~᧏����Ҟ1#K�Ȟ��%mЫx�ڕ�58����-h{��ˁ^Y�?�>	E��96l�)Y?�^� �;�<�x�|Eų���%.��#z�#��ϼԼ#��	�|��"~�7.�K����>=G"�˧Y��NY�<R�4~q�O؝�����ը������Y54�!О���e��]ya"f�h�_��$y@�Rê��Z��yT\��p���K���s@���\��ɥņ�Cp-R�h[R���	�Ѫ2A,��Tm9y�ȝg�4��ً ����LUu�Ξ+�:�A.c5U�IP�8�ܳs��t�*����BJ�.ɦ����ԩn�6��2<��Q���NM~ o�ӿ�ɟZ6���H�d��D���4�Ө)�� H+RY�����l�:ެ?wF#ΚX���56,�:e�W� S�]-�o���0c�K-�A��}�V�f��\������Od�۪q݌� ډj)5�$�+^���K�X"��V.���?����]9�gF0�Fk�B-�VsE+��Zs��dՉ�8s�F<�LA�O��$+p����@�q}�? �^2���<�{F�um�K�ë�v���<V�������	zKO�$!|a(�������#~!�5�>r���N��s��!� �ⵚ$MSi�o����P��Y ��l,����B���N׍Bi�4]�Gop}�;*~=��ǐ^SPۅ�b��sz'�6<L&�A�^R��}��1��''�k�S��G_>�\�dH2lr>��-���*�-\���	��;�TCk�Ѭm���x��:��@���#�6ņқ�5YA���œ������Q���Q��Di�w"2��X�h`�9.�}ʅ1K�_����7'�Ve�������ՔN��\z��z���(jd�?p�y?ܮ��=y��ڂq_,�
;)b���*�C!���>�����P�.Fv㑎5v��� D�%���9(��V5P�����z�j{�R�����&0bW��)J���*%�+�Ho&��^}	��lN��\���In��s�P u��mS�׆u-�w��QV*�[n힕7���xmV}�J%�9�����A.�aﳗ��b]=5t3��H�@8��������W4� e��������u@hA��X��o�����l;r����K�ikfn,C�wl��\��6	@�j��)%�IM�9${�E��:���*��7��oZ6�f3��Ylp�P���z$t�
�Z�_y���	\f��O�u��c��%��_��;o2=�����d�^0|cݻ,�g�Ǔ���I���3|���R�8X�9�C��衴��������d+;|�6����] 1�~�k�ł#�%O�%�}N�䢨!�m� ��RB�|�!/a�Pf%�Z�-��DH��c|�W� p*���~�M~Z�{��Ҿ	�4���S�-O;=E(Ϟ�a�~��h�9�͒_�Oؐ�OF�ϱ �m\#Ԃ�����y���]Ǆ������3J��.?G���̸���� ~'�������B���>P�	��>��8�<,t���%��"t���D#�0r�j=�5��㠚�g/-h�g���1"q���?�F~<�bPMU�!����"|c��Z=��]�L Ⱦ [�u.�@j�&}P�n��Iq�'�!��&�L���Ԍ.=�z�e2z��.�/`��}����d � �e�0%m����vu���q��=�=(h~�Z���.�^����@��8d�]i*��"=cJ���q�*F����AC"���x���ӌ�aqnj^]h���h?��4t���;;&��A����Pˣ���X�� !=������&�B�%3���2�;Zgk<�~��9��K�����!��%Ќ�0}��ė� ���U,�pr�,(�2�2]/���&�{ק�a����X�*�H#��@Kk�M����{k�Kpte����h����Ч��6���/\�S��=�7��Bq1j}mfJ�o�[��U�r�mF�5��X�R�I�e�����Uyp�gf�̼d�`��]��� �&>��O{�i(E�^�=[%&�(eĺ��NC��#$� �*������6�Kß`�A&u�s@0��85C"�U��l9�|<�+ޮKV��Ν�=�r���\��H�ꆽ�#�۲y@1����x=����3���A�/���i�4��כ��&;�z�L��o�F�A���!A��� �9��5��Ƥ��~���+�:�O���}3TU���|/�b/�x�̈����%��m��e��ו�3{��kg9�7_Hٜ˴o�c�٭$�NX2�����"[,�N�PS7�:�;�.I�.8��1>��-�1��e�D8('Ƴ�%�4��X��%l����v�.�4HAIv�ˬ���Rk�,#��NȰI�Ucڧa�K"_�ݎ7&��Fqp\.N���b��`��r>$�z.��<�<PE2��c�x�!z�@pU�}����ƣ�0u�0�S���P=Xߖ2
��t�p�(N����]f�SIɉ���)���zz�y��+�1��L>����� ���f�r���+A�5~�G��8;��V쟆�\JZ�jh�5mhΟ����	KM� ��|Al�E�Ӿ�9+Z�8��і��ؚ���`�?~[��%�%�%K<�TH۱��X�qed{�4��r}��?fX̣�V]�pY{)��`�-�ړ{ū���-����Fq��g��JQR�!_�
�8��~��yG��i������T$� ��/��/���7�q��2�X��?�3.�?������	��f2�]�\�{T�=	7�(z��= G7*���
�s���ӛs�({��h�"?�-|R))pӢtN����/'�.6�֓/~�,�Y�6�x�*WZ%G�L�b~�8Gq�������:cڲ&�I��C��E�����s?��]��n�{��R��ǹs�C�uߥ﫞�������z=w.YZ1bxBɪ����+N�M>{;/���[=S�/�+�g��̽�0��	�QO��)�-��Y��|��)����
L�i���l�x�
i�R���[b1u��<���_&2$�t<��:iu�n������K��[�̚��6� ո��� 6�X�p+\�"��=?S��Z+í��"W+�r5��Z����3*��և`�xY#��!E��KA������qq}G߉�2$�4a�	��a�6�m}�	I⇫�h���L���|�a�P£�������tiEr��f|�6Ȇ}%��i��z�p�rW6�gV� -����$�(x���8�x�ބ�l��p�CLaZ��N��h�k2B-�A3cx,��Ѻ]�?(��|xW�+b�9�������P�dxk ȕB���.���[2���t]8s����$��'_i��CE�LF����.�ȫ�;����P)Ɏ�F�]�����А�SQ�S\đ���V=,�	j�G��gg!��ޗ5#	��;��Yɢ�Zuk�Z%��5�}SO uɮ���>֌M�6����\� �^���X�L�өwX��	8���7,Ǜ����i�	4��<gİO����3C��ScOi�rx[ǫ���<_������t v��D��A�K��~�P��#��?�9)-��C�q"�p/0(c��o^����I�W�(��EeK��V�������ڀ۩G��1ٞvȜ������6÷s��C�P�A B�����0����f1?T�=���&�c����v}Ju�x��,&\v��JHZ�E�)zN����2TSp�eZ;���Ta�_D�&b��[)5�c�b{�v9l��"2_UR+�����0�ߢR~�^a�2�j����ҵ�/v���DD�jc�$AgSг�	R�ϣ�K����g�!0rާ\����D�w����p�Y�x֑�M�M,��sO>C�^j͙at��io�����a[�mL/���s�x�V�#��k��[RI��?�y�J'1\��G����I�3J�K�h��|e�Vq��i��;�~�kXzMt\��H0Vi�����ұ��Һ�G�㹋��Ou?�Z܆��oz]�%���;��^�)=�u�)|���_�F2���B�HV�B��y4���2��� �k�YI]e�R|�C���gX�C,�ƍ�}T����9(�h6>������;܀ǻܿ_C�Y�����V���&�$Jm���q�wy[;\���Ku!�������	��*�?�t=A)�&�݇H	Ji���w���KpNH�-E�pIz���<V��΃��o�H�T&�
HrJn�آ���"��Z9���R9=v��ȶ�>j�w` ��*���	W���3ϵ�_�']��S����e����b���o�5�au<��"K�xL,�Vԍk;����
*�F��!"	w�s��`�����4:FЯ�!ԡ�t�Z��B7K;N�>ѳ���x��g#ł����j�����3���\�<�H����p�C���|=�@��R�x$(�~��3�t�Y׻ߜ���i�b7*�����b����>t�5b<�%H�cj� EisS�E}�>&a�#l� x�*���^�_�Xh��5*I^h��|��I^P�G����{֟$�L���~���D��A��p��a0t���q�Ɂ�t��`��"�fи�0!mǨ5Zq�&��o�p�.�Q�E�x��w��BTX�yZH|b*���_�l��� CAxj�2'�d��~��,SગH$i���~�	�Sd�/6�t���4Mkc!amk��ӪR`RBo�ws%0���C
�qX�3?�l71+�s���a��aw���Þ�B� K^��F46��I��Z�%�p�c���(��'��s�uXzȪ���ۤVn�;u���\��g�
@��+��80�C����G�3صR0�Cf��O����h�0�;��l���A�K;�&���"�e�܈���e��j7]��L�a܎ "���S���u��1>w��$a�)���T�B���"Bc"�]������TWu��XR����#��������>���t��1+����P���,9@�JxI??���2���K�g2�(��������<p��1@�֗�L���w
��_U�VT�����HmWܤL�p���uˌ� oC��Ba�xI:����և�P���ޡF��K�q*ժa0s�()N�WCzC⊲���{VM
*e}�?2f���@H�G�B� ���PrG����R(A^_�����4{�*?a��g8�9������O����*�VF�'�B��v����M�l&�o�"��KT��	d�&4f�-[F���`���*Ҁ_S2u�@��f\W�p���A�nwcSǹLj�L��>a�N�-�U�q�l����{!�bF��oQV�)�mz�>�P"�V�8�LU��O��h���z=���~��9��i��z���~���D�V��ˁ,��r}�]@Y�3Q�H���,F�N��!Y�%F�ܷ����p(uJ^6�C��i[.3��+�RB3��Qve�:��۝�D0�ۂ�t�\\1����*܂Y�r�]��>����V9PR�ս�,���KM����ȥ�Ad|�t�h�L��V�`X�qS���>d���O�t祦��h5�99����w�GR�p��g�cĩ��Ÿ��@���[uEj6"v1pH���R6�yr���zS��ʃ�p�D|�[����7��+dk��2�P�� A�IBBI�U�/,����H����H���P��/�C꫅��� �F}�g5����;�6�fOL�\��5�XK���n���V5�;.����5�f�ߎ������0{x��^|j���8;B�O���&��W�	%�bP.MM�y�g�.F��jD�oԗ���Pzp
��-0��Z�c����':Һ���,B�|�Un�1�}�3��YQNߔ����Od��p`���KvuRڂ�`�3�:2�K{5��m� �ͥ�FId�wC+ԄT�pE��g�ё�h�v����7���sB��'�o��^k�5/��^!Ձ+��)�}���ԣc���م��[*��,|�6y�:����s3�����rY�~D���� �R˳b��c��e�ȹ��ܼ��+��,w OCE���<�I��0�	ŕ��#1h�w~7.�DsIW���_1t:<ez��8�j�6;ތ�����<|�x\��`q������ǧ�'\�\��{l׮.dJo԰/ʚj�5��_[\�y�Y�(��nD���ȱ�w���$��2c��W5<� .(x��K�G�J�j5��k��^2jO�G둱Bh��B8���rA48��S�l�VT����8��!R^�Cw��_��I��l(C�/}s,8�.�8�>�*�>�=S����MP-W�3�X�	*q$��/}�Bێ�UՖ���*KO:S{0:�{��Lg�a�d�8^���<-������[�k�ʋ[�6K�a�v
I�Ll
�ȪB=��$s��v.
�H�0!��<Z��B�< �6��r�w8eM�'O��� @A��:є��*�����9
���A���˾�l"(�s�O)��3������T�W>ߜ������#�VC�A����jI�+ڵƿ�8�o����@h���ь�s��)1��(�b#��3jCI�I2p�sK�p���гu8�F�^��C!i�V�Hl���:����6�zԶ��T��"�|�vb��{�(RV���FY8<�s�=MS��03;��\����� �Y,�B�h'Vv��;�5��z�f��`m��A�E��G��l	�wFG9�V��J�#1&,��fw��Im>T�-�X��G��	����BP�!�j�*$|FE�-�ۮ��������[Hye��D����ܵ�ZpN����k��v�l�#�tJ�������v�؁���#�O�^c���kf�0$jz�u��\3�n����ک�rjg^��vt��-zd� x�����a� ����J�Ub#��M��S>J5n�����(�C��u�����/��tp�vJ��ϰ�0�Y �����������ĸ���٠9��N�$�G�~@��=��@H�@�4����;S�m(�kU~R�Xjbu/��20<�e�V���̈1(T���	:�Bj4;�e�^���sS���OH9Ch_��k�ߡZ$a�6f�[��s�]5:Z+�Lh}O*Ӫ�QZG��E��c������+�V� ��?���⤣M�7�D��M_�;*�&Lij�Edּ� ����=0�3�'���c�u8;�����-lk`}#�������H�il,�>�!��{�l�W +�'��2JT��t�A.�������]��J��b�1���8/ܦ=W���5rR�Kk�$p�O������d����P�
^ҧ��f������i�k��T�<�˘�'�X�ޢ�4�5���?�n��n��K��p ���Ğ�M	�
�)OTk{����~����ӧ�u������\���:y�Ԙ��j�W�[$P<�ֲ�=��F��+�v�Ա��#��moi#Ym�V��xO�پl5F&rZstv��9cÒ�^_4D��� k�f�-��Zek��O���w.���8�V=�̼0�Ī!�׽�W���#�}R">)S�Z��D���!�≮NA�B��IU���v��\#���cL �u���:%���GS?�/�0�W��'�Ң�lb�$y�T�a�d�:qkB14���[,���Ԅ��l �m����oV�m�P�MMZR#I"�&��8EMѠ��kp��"#�F�8CC��/5�9L��ǥ�XC$(@��g�6���9���U:���A��X�P�)�U��U ��:M�Ga���K%�E�Cwv� �����v��i�kS��/0�t��5*V�)�����A�%`�I�i�ѯ�[a�ن�|D�� �{䮱'�h���l�]���0z���I���@��[i�9V�[YB=h����������Mh�a_��/A����Rh��.6H��i� � �.v�V9p���C���NSh깈��.ݶH��Ab&��&���!��9����MD��x����,Zs�s&ȴ�)�c�g���BĨ�fD�%%:�&!�F�����1�|��M� P8FcW�P�\�d�N��������B�z�'�n<]��Ӂ�փH��*)����V�Vz�qi��e�`���,޵�TU�P�*��Խ������@�)�B�+���eX���o�L�z"�M�q0�yX���H*�#S�E���D������0
��|[zD�/�����IZ�OQ�ۀ��z�Q���O ��_�P@��9�&1�n������ݓxL����cv	�s��-E���S:r/w��r�@j�q9�����ր��t��BK���"*�|���v��©l@��T���i�ȃ�Z���6� ��j!�?���(S��?eq��wLMe�W��$SA�=0�c����J�|_v�{��p'T7�F;0�^������K��l���+�4?/�����Jr��
����JK�h,�<ﭪ�������H����T0o�_,SR�U��̔���ܗ��S�j�9!�G �5��:oN���Y�D�����l�S�5�<���3[��R#J�V6%\�k�x+�{����\�Q]���0��p��*���h]��)�F�*9����-��wr�-��O�ǵ�[ ?�!Gm���$\?5��-ؓ��G
���HքQ�5l������u���(��t-�e�=Q�$��S�vkJ��%�s���0�T��Q��&@if�vC���$SK֒4���N�~�]޺�ѐ(��]�hOY�YՁ�W��BX�j��gl�Pq,#���ir
V{L?��*����R�����꺉� ���	JS\�8)'��_��W�h���b܍O���D��a�2
���&o�����ޠ+��A���I�6�mC��8�(�Z8�z����>W<�(�_�qĹ����#PQ��o�v���`wPB�q�l����B�����҇��v�7�e���[+Q��!�~ax�_,-��ˉ�@�D�OϾ���4��ྒྷ��~n\_�q���h~(��fx��6���h���(#�Y��2�0�R�ed��#�������@/n�j���r�D����)[�a*� +�q���vDm�d��Wؒ�`FtR����Pq��[�X�Kd>;~$�s(�!w���]�*Rױ������͖���M3�(ș�
��PdR��q����,q~cM����)Vg�Ӧ22ebzzy-��s$��Qj��D
�:@�O(���$81/K.��ŵѽB`�M�-	�>�8{�K���Q��.�]�e�B\ϛ���&g%�)��mUp������-���L_�����R���=@,��.R���.�h����Bx)(��T���{���Jl��\����\���b���g�pri(���7v���;�� j�5��1aBù����a�<B2'�½I񇬻� �ͣ�7	� �/�~Nq4c�lPmiHO��T�D���ӜD=1f3�=V�2�yZJ_cި
�X�SO���d���ƶ`(�F�S�̄'���I~�$R�xhy�F G��*c9-��,����Z$�5�M WK�i�����r��ҿ� iܒ�o�q]��5Qv���P��U�I4������B��+�[_>v_DѦ��l�e��(v��E���Ko�Z���2AT���rJ�1�,,Pj,�u̿�҂EN�{�y�)�)yu�e(D��y�z�5�aLƃ���P�jC���:��F&��<^2|�g�e9���O�mK�}�����*�G�5u���Y�t�(�n�"bT������l9k5	�4А�m�`g���O���>Z�v߭i��
��_,N���x|���u�f�Ը* �?����s�� S��Cx�����4l&��X��>u��wb�sP����z����,�l�G����	��i#�H��j:����h��!n�=0=B�g{��嘙�}U�Nδ�M�!b"������]���C#E	"���_�� v@k=ϟ��GE;�|��@�EgkN�����Z1M�E���m
��zf���2��)�6ݶoBX��I�+�.�R����������#���l�p.��Y|�3[\��n��]7��'��)������.�����˼��ĝ����S������@M�?���6���:�8կ�9?���eJ�m��=�/�5���~�t]�{$������j�cr-�aHׄ������*w���{zV+���u�P�u��ʡH��((7���|�c��=|����{�%���l&�\�@�I������#gr�cg��G�X^��-���+����\�!�E"�>�L��"�
=3�"逢+b�w�*���X���i8E>*���b�yX�iq���6A��G�Țv�l��r���%�_���P,�{L��9u�Bz��t.\$��3��Jn�N�dWA��-{e>>0�q��=��ȰВ�k���m�*4�?���T#����O|�-����B��/w5�������e%���^�;!�J��F�柬R�u��*���������#���f��;`g�5`�X�'�nvu�Q��@�&�5��Ps�eTd�ا�������w��ӏ��a���ؼS�L�_t����(O)��k*��?/�=d���@�y���`,�.��b�O���`��.�1������T�&D������S�`��qH'����r+���w��Lb��Gg�=�8�`%����D�N�	���ɓo�t�#�����b�n�=p���#6��t����P42}�bxvl��}��G��v�`�.�-ȼ��8uɝdC�7G��	��M6�{�� ������xP?�k�^��S���ەX)��o�E�m��
�5U��3oI���j�0�.r��U^��[r�;��V���n|f�Q����yi�5v~��b���7R?�F��K+&]�e��Xv ��������♊x'@l�B�.P��\���|�f!��y��؆SY����n߭*��H�Aƙ��C��W��H��E����j5Hƛp�w�=�h�Zo0��偷�+	uzӠ��j�$i��s5?H*��	V{�]�H���}�rt��vX��<ն�ca�THM�7���n:��W�9�+ui���ᑼoN�]��O���j~��|��^�x����v��i�@��cB��߃F�N��:k}��F�]�#P����3 6�M����b����<@N����Tl1���4�o���{�@J�l3$5�O�[�7d~�����}�����൳�� ��z({Q�@�N�(S`0h�41�?)JAi�"��W.A�M�����WT���P[�'3�d��O��M( )(��ޖ��k��Q^�Aw�L�BlE�`���8�)��C�H~6p���?^!�ߑ�wG@0�u%��瞫����!�
j�U�ՠ����H�hkk�H8s=�-�8,ܸ���H���d��i��ص���|/�'�@�u��x�\�<�����t8h�h�f���jd�1T���(����jy��7�\�?o��G*�x�k�&o�H����
�2�0��!G�?�՚M{�h��F��`��gɛܣ���fNڄD��×�9���S�<�Wzskw�v̙�\���f�d#�gܓX�D�ɆN��<�L����^��m�u���v_�r��J���K]�q&�&ƍg�&�y��
G}�Z�/Ό+4tE���Ij�i\Ђ�A��%K��D�[ԍo�]�8Y��WjC�'�λTw4pDIC��d�IL�
:���8����X�O�S�Llo����*?T򉋡��o�$U�r2���i#����5y~����]�(�������q�{*�Ø~�E�?
��Kj���!�Q��aUQ�ͽ�_�;����fx΋<#�r3Ψ�л�$@�CZ�4Vg�m��,���"l4�U_�l�����_3i�-@�8lX�=)B*J�}�Q_����X47�sRO��?{R*_�_��QwT�:<���9�]���8��b9��R�l��DcuA-�w�VsF7.{u�G9�({�+��M��{z]�@y��;��iO�J���#N�1�
���$� ?��7�{�[o0KX@5���gJ׼�6C<s���j��GMT�c*Q
�9"��H�|���g��[���FQ�����4�7��=��
:�;�ED�M>s�֣�8`�9��7J�ɯ�t�~�tB:���ͯ�y���➙���U�n��u@��o��P�;b9��$R��]k:XL=��'4��n
ղ�1�����zp�L��(a�k����Rr�ш�Pf|���EE1���	:ԭ�ֱũ�65�!�R���&?��'{��{Mڭ�}�%��{��S!-���Z��Q�JWӈwľ�8��6��Wĥ7�U.����4ܤU�S	�G�wR�4r�,f��J��!h�P��v�xv@��D��Y�7 �it���\.F�#��3����)�`�{$�ԯ�H���=�}T�|�\���"�c�D]���6��s,@k�� .�#�~�%��5��/�sY�&��k�h		���&�kC�W��T}�)Qi��А$H@���w�83"VY�B�ΞVx��?��;߁�|."f�5n���l�a���X���A[#o]7h�r���W��l�pG�i����D��<n�HR��Re$~��:q#\�z��4�u���r�0��&P��m�.�.W���,`	��"�DZ�_7;Ε�Ө�m�1N-?о����0���ʽ��M�|]�hk�"�����{}OAF�P�Z�V:��4R��s4��o��	A�7�}$�Q�ex<�Fmt��j� A<[5���3���Ӕ�DJ�b�3��G��&�*n���f=���zNS������؂#<�{N�G\������逫ۈ3�cΜ��		19q�G�dA�Dr!���(��xD`V�];]MC:f~3F���B��b�ڜ�� �����#]a4C)���sa�Uk}#0�f�v����G�I:xф^s䷎U<�Zx�a��%��<V|��O���`�Y��Ph2�ʝD����8�H���Nu�������U��h��_�eX[#�]�W�F��4�Wt��D��	K�],�������� ��a��z.?�:/x�څm���b�pE��CO����\+n�\���~���nq�z0*�7T��E���;�;v�W��&
L�k �k�x\����8s�Qf�� 7"�~�̼TQ]��{�R��{wG�. vuEP8C���Dw=Ei_�?T��tS�Gh�G˺��,��"���9^�:�A^�ܷ���s��G�.%�|��̼7%K����?��F����Q'i�i�K���U�A���U MG�w�$���	�S�'`�o���Ϟo�h5�ѮQ�]�*��x�è��jTA�����U��>"��k�k�{�m����h'��'�> i3lY;]��7	�#�6���ԩ
Ъ$̖D�lV]c��6u��ҳv��W%a���2�[�_m[O���%�MP7���'f��'�<U����BPݿ]�Ϲ�}�|�l�@,S �8��g�ac����l3'}7x-�%6K�����k~?j'��qJ8�RB���֔ 65 ������e+�D�5bOQ��	�{/�)YM��R3��ƽ�,�s�Bz�zT��O��ۈXn��2$���U�ܡt��Kq��&�o!�DWBP�A���j�V����v�v����C��N*��14�hLr����V��5���^kԤ�]l�ݎU��X4��&��cRuڬ�p_���2-��OvNI��}����B��/��k7�����D-ɉ����5i����CU�9s��[X���:�k0T/x�FT�G|��+sY�8@���}5�s�ۭ��� x�����Ԩ��U�����ct����������7�+q!5<�'���J#(�#*��œ��e�L�ޜɢ�0������6�3�awh�ҕ���r{L���
��!6�ǃVc��u��A_ΏLol���~�S�>�����͐�d��Ŏ[A� g����;s=v[�����ژƽ��(����x�#㒄�ը�\I� ��A�D�Xt��Uiܭ#�MeB1�2�H�*}5%>����N�bN/�W�!�ǽR?F�ǆZ��Ie6��o����i��l�W<�r\���h+�:KX�y�=��-ΐ�"lV:����BΏο��U���Q���t���t�i���I��3�a���\���M[��v�f�=]~ZP��ɍ�"����=A92�g�Ű.�4�|]9bt8��D-�U���	���7"e2�a�-ĥ0`�ʒ��/%e���A�3'���
�e$f1> M �W�-���� �@��E娽ʫ�vUpI���qN���K��آp�e�b��d)����t˔7}]
�C��0��>'V�$.]C� {I�����EH"/�U���\qu��!�y�����/�=P��>27�1PS�"P7����~G[�Npի�P�-3�ϵ��%�=�ݦO���c�&�Y�J��v�sg�V�, *�1�d�
��x	� Q�9e�Ŀ�O��򂏂	�Y��\�y��h��ǝ�������t)�G�emU]��9��Zc�@�AMR(S24��M�k������5&�<?[��|D,y���g�����Q	738�����Ut���C���8f�B��+6qΩ΁^�������p6�aųKA��f�����E��6�����L�9��/yykD��[�g�M�Nq�;�`*q���^�ZɈ�㔔�w����5}�#��!���U��T�y;Q�������a[!���×��s�=�d��[��9���I�̔��rs�g�i��өe�sl6�cOLU�cSə3p��7��������X)���ux\hlW��7�0��K{e�/u��jc�e�Ỷ5�E�r=-=qr+��f��i��xEz�,9ÑӺM��/�%��y���'�qލK��Z?sdGG����S���ۥ�z�:?�(�}�e_�*/���q���M|���/Cr�OM /k;؎�G OC6U��@���P����[�_���-_�3��l�4CR�|��U�jg�$Qq5�(a|�d��i�T�rXs�\�b�|Y�r[�Sp ��m'�G�S�?�>t�w���@�@7����p�`!w4�]����;�H�����~�V��zX}�r}?��>�Cs�o4-
̩��۷����KO9
0���N-w����� �(�կ.Ă����z�� �_��q��6D� }ץr�>�cFy��[H�/�5�Z�m|�Ʋ�R�/h�-0N��7������4E���^��ۣ�D{�NjgT�Eo~䱨�9��ˁAl>��%��ġӉ��A�����<�IbxZ�������V�)\( ��SRT(�Ƴv~9<#L�ؿw��z��������8l}#Ӿ�9J��^�č/Ek;vlv����"�%g?οoFSq��!��"W�S;"+P�Q`�Yx���=������E��)Yӎ%�rd�}&�&�U'��%���q���g�^R�y�W�p���+7��(/�,��l2`$�8���H�-��"���󬃯Жe�,�G�J�^��g`��{�x��sÒ�?6[�E��[zE'���x�K�
O�~��ФV+nK
 $�<t�1xU�f/-����	ޡ��εx�|��?�V
L��N�W�\t[Ժl��o�q��=ߎ%�!o�k(�C�#D�R�+�u��ŌtG�h�P�Qz"��O�4JK9y�δ����;��A���*�����_wStzp�[Zb>�H΄��B.�K���gk�uI��n��/9����G��q� �{��A߹�y���*Ǵ���zg�JuZ;}�~2�s&��3Ŷ�'u�uB�[�6FE��s��9��:fqa) .>e�i�뾞+D�3������Qm�Z���"�I0���mY
��^=j��vJ����|ya�eֲ�I�pW��ݡU�S�����#�AP�8�b��B�3)n9����n�)���	nu&���Z�s>�%}j�gze _EK�6e!WK����A)�~d���B����(.� ��h5�[��fp�����u^_�y�G.Ւ��geM3\>.��z�x�����Lc�
=*�@�}sy68v���S��/w�w�2*�8� 8�F�{�7�����Nt<�;4'Yj�m�`�"u���K�XDf�<��r�'5����M}�v$M:n䯿pl���L=�6�'5��R�Hlhm�p�4 �0Լ�|��dùl銗L|q�X�Y :~�󧱃O~r��1��c�}k|�}���k^�<�mB���,!q��8��E��V$?]ڼM1�L����ڄ뒗�?���+���Aa�>��N��K]��s&ן�jY[|�>@��b� AdXxoZ�sN��q8%��7��Y�M�d/3I�@͆�8J0f�u���-Y��F�.�Lr�2�b2N4Em����(���)3d��i��1�.�Nw�0r�,�#6lb��/q�	��da�ZF3J0�OR<�!�B�8���,SE�l���P�o�j�Ɂ�}�>0F ��/��_�� +�B�h�C>���h��\���~p=0p1�	��n��]'�N�U��/^wYz�2s8�*����	Gs��MsP��UER��Б8N����Zž�Q�5�=�{�D�W�ˏֻɡ
�ҠaSZ�s���BI�����q��[u�q�A�a��":y�P����������yY�m�������>����\�w�q�DGx��7&��3���ц�����]cy�Aa��(�Bh 2�YwW%<�L��ψ���.Jd�������ޖ���Z{�eS_� ��X}fTӻ�ȻfζM��6�g|�F{f¼�d��L���� $�(@?�@�s$w���^����_I5�����i�o�_Ph'�wx:7<IO�̡v}�''���Gev�8XIg�{���	h����|���Q1ܱYq�J�J�b,�m_����������7�f�FA���j��'hOY�G�p=8�\�T��-�O�z�&w�+bY`\�yc�aA^91Aq����Ѐ��u
#e+��Z�i�܃��^;Y�����G�{:_��O�}�*|�sx�a��Z4E�kM�y�C�T茧g��bBW���1\�,L��� Jv��7�IC������W>B����`�Z�7���%�� �~��l+�����
��-��;�자�*ɑ[��\^�$a�������[ˢޥ5k�>*3�Z��4Df` Pp���T�9D�_p����!��c�]��(x@�%6p����[Cl���cV-���j�-9+�����3���d�6�������#Ko��O��U��g�ÂQqL��l�w���$�Z@cP����$s��+J<��f E�˚@M��Qp(~p�<\�ߖ��dh�*��5te]�H�ME\ۂ�ȱ#��zK�`���+�u�8R�8J�k
4�D�hZ�)e��Ji��KE��Y!+pzN�9�V�/cj�����44�L�5n�F�n���6	�"��$�_3 ����_��C�381n�� ��|� ��Q�v���NB����m��Y�!�[���/)�� �aUΈ��r�#�>���aꢑ|Fx��S���4UL����K`�񇞗1�hQ�(�n���a^�J��I�7IOC)��5�~����x�ݺ�Y��.��Z.����`��h�.|B�g���)V��`�3��[ץv*�sF������ō���q\��1���$��&_EH��m`6'I>��P�����6+;��d_t7���7V� ���*�E6�Y��0�C�K P�~t� ���
��h��A�� �#���@��ǫY���ڮh�f���A)}d��cP�<+���AP����Nu�o�G�8F��ڍ�ϡy��l�.�r�k���0�w}�q������I�I� �3��GLX��|cD�U�J��bi��֊t!Q����&��n+�X�b��/,o�xE�-X�"�3�$�n���*�v��;�'�N�cʗ���(�Gc]o^j <^z�)���f,��"��⧅G���U$�9�#F�#�֒�Dj�@v��a.�x-HE��*�I�A�M�z!��6m����:�tk���ˀ�[A
eW�,E�j=?-{�m-�o�����js[�L�����=�@�D	�LA���Sv�SX��$���&��:┅pS�G�^ {ZY-kˈ^�LM]�w*�M�~�ȹ���L	;�����b/D��LX\݅��aBe+�1����ἦ �t�1��"Irxk��q��Z�\C�о��,_x
x �pB�ӝ�dZ?׻��K"��~�%�N�(2u��]4Ȉ�Fm��b��k�C�J;!���L���{Dn3a�)��7b�$����Is�`U'u6�i��ٳz��f&����] �n���\!1�2�"!���BKa�14�&w7����[ek��\�����cZ��`�>@g��+��6�s��oaU��[���3��fR�h:>��]��d$w@h`�YM��=�`���|b)��l��­��G�%y"�����4�dD:�#8r�XacRP���>���醐X�MY��Fy���P>�"�q%n�EmJ+$�!`�z�Bopf��d��[[�@?BO<�������rg�j�g@/kwU�������j�U���V�1Z�y��Hg��ln<\ݚ@�������Z|�9%�m�P(�X��Z����<:XI$�Y	���V}pF�T��%�Ҍ�^	��I�4[|�-x�>�n��gu8�,��}��{�������qv��mz1�R�����p�W}SR��_^����G��&���i��1��	S��Z�57���"7@�0�}z����R�N� us٤y2	���m㵽S���������i��JgG�:�¾��tv+۠�p�r�E�	�l,B�n�)	�0����ԙo����v˫�4�v���ZsK=v��f�K\��1��r��<�]>O�ӧ���2�e>/��Q��U���w�	-�?�J7f�*aM�M�D����<���&�^�U�˭�ʗ^�o�N��Lu+���c��+'C����o0�SZí��<xu�;��	�7��d9�� �᝿R��`�� r(e�"������I�L��W18e�	ڴ�>_��T���Wլe���P�C�/��d�Q����}��6M���z5�����1vTi ЏBS�uwNˤFВX��9ċ�@��qR9p!��١48iAz��d��e_(r��y��`�>��T��.��jk"D@��3��$h��[KH)��|��ד�)4Y<W��ZKQb��Z������7҃r�yPs�k��&ka���l�p��A���h��Nt��rO�����z��U�9I)�-��<�Й\Y�(�z�����2�[���.�3ӟڣ%Zx>7�V��Z���3*�J�Gϐ��D��Ϗ��Pv�(�.���[]���J�0R�h��~���F[(M�B��H��O;x���4PϿ@$��rd�^���eSj6�aS�
�N���b���u�,i�p�^cV'�KJܻ�6�h�[�4yr<|&iW_��l�J�C��k\c���������R�О�$���%����R���*�����"^��Z��a�u!Z4@U��0�(K��)��ȟ
<b.�S�e��r<kw�+�wR�&��&��,��A9IP�i�C�����*O�c���PH��lW���T[`�����7P�<�� ��r�7^�C�x���@~3���<���_Άo�İ����]*%IQ�_��^vRXꨮ;|���u*\�v֬;�=;�Y�yt�(�M����(vZ�Uo��3V�.��Q��cY��B|k���+�}�r6��
(�q�X�F����G`�m;-G�ڷA�Ħ�PUS��f��A}��ykV^0x��צ񊋥���E����28�;
��������qJ�k��^�p�bL�^1L+f���̦�����M��^"/d2gg�!�3�N�5ʽ̈́tbG�d�f���J=�Յh�.�hg��Gw]n�vǑ9��(���X��6v`w����FE^��0Y���)"�HZ;˶�����ɨE׆ʪ$^�k�R�/ߠ`�V0�"r4��3���e�t��x��l���a�>�H/�?'�J�hy}��B"�y_)��T����t��)�(HcP�C�_���jh@���J9�8�#�}��j��
4���O�.#T;8��g!r�>o��\[B�ӈ���rve	g,|���:G	Z���&_O�2G#�:<��)���$W�7j�w�����IY�:��5/`�+��H�dg��B�R�<BZ�甮�A�/��~��PyE�]^�q�=*?��i�^v!��F�$�$��%հ�7a����w�#�5�b��ːΘK��mv`| R�a-�~O����P�k�:ˌxA���F���9uߣ��E���x�7�N�=׊�yL7��ￍ]�^V��vF�L`~��mˠ�$�2r1m9��fjZ��u�øT���!��X�'U�!��ٙ+Eɛ��<�J�
���|��y�ymQ�}�@w�{oWeR�NQk�Rm���~B����|�ی�D=T�F(�����?���8M,&ŕ�o��>���� ��7^|�����J�$~MWN�2��F�΃W�scJج��M�2��x�6�����f1;�>��/���*�1�<<P��Nf�8�,����R��J��}���R���B�J��?\�]Ɨ��y�v�t7�I��Jf��Hl��f����xQ8R�jS%C���e�� &�=�2H$��G�'�.ɩ>I���<H����_Ը�4�K�-1m¬���ecP��Jynm�<����X��#z���̤H����ұ���u0��� /��Pg����͘���rm"���(�h�m����
�+^�'�4J>�u�Τ�XFo��H��ý�-�O�6,�,�]�\k��dy���.��vt	�*�n�m�1(3�[�Q�!s�9qAdy�ߌ��:��+P���7����#p��3٪�	(�� ���߃'�ϗ�;6����LE~�=�O(���$gͭS�� �̼O�ŋ&��?W!��N�0���JE��u� ���6k�9i#�RY�)���ؼI�yF�`]�~�H�*���'���aR��h +!������u�b
_@ex$$�m?�Y`�k��!C�?Tݞ��HF���S��gr�#�џA�>d4{��էR E'r3���)�[�&=An�K`��ٔ�Z��W5oü��7�<��ݸ���ˍqe��l�o�����D�r���h$��G/D-�;���"��I�)���]�k��䈾|�A�R|��U�3�!���rq*�iC{fL�VQܫi��4(�r.�D�mkk�XE�Ah�#���q���f�㽲r�KR���N����eMj�AG3�CW����muA�����*#>���R��v��Dn� y��>I�����!�� ��<a<�{Wd�\,�Jl��ړہ�2{P��/bl>%�8Ш�*"�򨹔ד�]L#�����y�
-*�������g��Q.�Ҭ*���,�/P<����C��<�-sH��3.���?d�M^&a'd�/��>䎩h��L�s���y�<���K�[b�h��j2������F����R�w�#(��1Mw ������$Qk���U��C���|W�{�K~��ϴ��y�qE�gNF9���fIS���|��f���l�����ء�d9���g:*J�7�zz�DJ�B&V^}v���4��F퓻���7G+!5��Ow�c��X1&�_fu�4����b
�2`V�r����kɯ�\�T����C����1S�GM�����H�������s��&�&�MM�Ҵ�Tu�_.�9�K0o/�Z��oਠ
H��Hَ;�P�[�<��g�Ҥ8>��ڑZϛ���?!U���P��o�Nq����NA��Q�'~|�
�F�ri�@�K)|t��N�9`�ֻ�`-+llr�E��'1p�N�n������8
��I��r�� ��s��L���R�6`ܑW�{+q���x�Au�}�ú6��@Ρ��B1�������+���Bk��z|+���=���-�bi�K�s��{cr���ɶ�KLƈ�V�1�`T*�lVʭ�P�l�\���"�0�<:�Z��]F�BHO?�Q��#��o[��&�`-J�I&���ֆ�FG"m��r� �t�h��@��{(n�j����6��N��Ɠ���U���(�V���F��g�!qd�*cн��,0�bk��B/��5��|4c;1(��kӽ���U~W���!�<��}>��Qu/i�A�������X����L�(�U ���~���F�[#�% �g�5ȃ�
�0]�6�=��vo��:�
iS�k�������V�8?�(�Im��8�v�����_<B֨4����&C��R dG4 �s�b]�A���bn�b�ʬ�"���_Ȃ+�:�r�8��M_<om����Um����b)��?��l���u���	.G�Yr�����~ɟE��׏]�T���J���c@�SfXwj���@���Ϗ"Ux��!F85&\��,�	U��/�ˏ���j4�$�۶�w)�D��O�ywC��Nsp��|�U�X$FJ����]�0a����EtzQ#����eYC�$�?9Z������P�MF�7��o#�%B[YM�dF�=��{2ۘ}�y�6�:%ϓ/-�բ�]O3;t96Re�Vſ+P?U�p�4H�F���#�A�X��z�@L�7�!n�_�9���O���{ 9����z��fr�Wŀ�΅GZL����p�}��w��?3[_@�l>ڂ{�%�ڛ#�b8�^/���@ۡ&�N~�B�U}_O�i�$*!�l���F��:})��1�$@v1Ź��W�-�َO�0��]�?�w�����b��ޤ���G�<t q��ST}�)�4���s
�y� BW��A��R$p�����\cV@��F����7�����-��\��BJZ�D�$�F��Jn,��_b7�p�0�G�X�PP�DB�b |�8I�F �Jk����-����/�J�JU��"Ѣ�8���h�h�-0���$�s��?������7��~���#*��������9���?���X��������-���}�{5,ڹg�؇T}�^��VlE�tjE\�P��r�x��S����m�UW��#
�yl|�Ǡ3t� }�N�>����%�����@x��ـ63"�P�4�ܞ��?V?��`�f�wHY:����V?X��ϼfſ��� %^}A���2v���|��i��A��)b����I�?�{���;��EMD���u\1hp7' (�s�B�� �fɩ}���I�ջ�yG��nߋ��>5ס�qͷ�~��A���+U��7O��^b���S�E��٠�b��Q�m]BgD<�1.[T~dRk.�	�>�f`? �K����u8��˦�r�$km	j��'�����5��֭��B�(��E'�~���'��v>z:���!��!�r��J�>����ܧPw�wJ�yvcw�:�|A�B�)-K}~>�����E�Z�yA ��}v�`�`�z<(2t�֐�-����H���Gx�M���ߦ/MX�;'�M�9�[���5m����5�;�K�7LT�d�߯��$�I��Z��CŇ(��1���s^y�M��?���;��h	�s2����h���>M"3Ʒ||��X ^6�:��b�It��[����&2���}���2�8��`;���N.�p!��-"�y�
5r���K�C]����I��Ǘ��R�(�B��4�Zrl�)n׶d$�یi9�t�iƨ"��U�Zռ�+�Y�t6C?��Ȇ���+���(��)�J�G˂�b4]��Z#rD���\�ry-.�?Y�{
e|�����m��E\�}���T�韑M~�IC����Y(�|r��<%��g��lr�K������-�΍"+B}zn�a_d͆r�^l���{z��f���	ٚ�B)�T��Z�a�O��5wD49��x���`2(�R�>5g�z]�W?4�|eD����`C��������4n���*�z~��,��T�P|�D.�B��GV�0ՙ�)�x}NU�LEk���Ј�;?D�/���a�w�x�˥j��$�E���,� �M����V�WU�eL�U�������������1մ�p�P�Z��Ƣ���,:�X'�Q��w�B/�Jh�I��'��ئ8,�8p���	�e�zp�)":<Q��X������d�N��s�D2�w�>F��i9�{Lq�ů��8��n�˲�)�0�m�*�ě8��4�~Y u;���h���ҷ
E;I9�=�av~���ۇȪ[�#��;��ߕ�����/xITBL����ެ:*��S���-����BY�c��ɂ?���������ag�oq��h S���.{2�d��ȼu�(F*i��2� �3>�KG{~��'�э:��$�LY9
*�(Y%�\]��Ft�ˬ�7��u� �hE�}�F�L�%�~�]|��Y!��zD���u�����<n��k���4N[Zu���O�U��5�0
r	C�O
�{kyG�{!�	ò�'7�m�"����������"��W�%e�k:t�j(>w� �5�O"g*K��[h�]�:���,��`��T0�EK�en7_(�dO���7��x�S�f�wJk���l���(���7w�#����ۿBT* ��O��ة5�Jq���.t"QTۍ�+�-M� Ci�;� ]�f?��y��du_(t� ds����x��4h�'��c���KSɷ���v�����p3t�>�d�Ò�PQ��:��SIO�H��C�g	���
����f�� ��DR䝎�R�֣ߚi�h�7{&ͥ�6�"Ծ�Z�]L��V���1~���������D�I�Uv�_��
Bb��i�]ɔ{���w�;{oY�mr�}H�.AͰ(1������0��򍻄r9N�$Y�O$��n�����E��h1`�����1�;%�XV�k���?u�ὤ�T������hw	
��&+��f�ӫSn��ON�{ݱJ
3I��D�A���!�1#�~����vǩ�Mh��d���Q������)鰌N:E�W����-Q���o�`��n��'��� �Zi@��=�]:IB��w�{t��1Bb_P�0��9�������i�%Y�"�3ٰC�j�y��[NJo۪�d�����pPv�����D��jx1�O�˟�7��%��3{)����ķW�;�Bܭ���ܣ,%�MGN"?3L�
� ��Ȧ�I�O�����V�����R0-�#^*��I9���0ԁ�'�<I[��ʟQn���S0^h@�W2�T��tQm��{2%0������9��q� >>H��O�D/�ܩfY6<z��z��� S���D
��vtŇJii�>�ؗ02#�y��AN�PU���lu�o����%�O�}j��j��M�bp�_�]�������t+�|̵��f�/����r���N��u�?'���~C�����U�mV2h �hp�������������ы-NJ�kd]��:�.�ψ�hN�-�<+Zj�_�����(9P��+�p��α��?�)XЖӵL��?��q��\\a����ĵ���+�^r��#^��2k
�c�g:�P�����ڧc��y�UES��#����S?�*����c��l�2t_I�^�Қ�$,��f:�)�F���u}B���N�1�~ /��s*k}4�y�OI�2�u�U2�0�I#K+0;묌�m�>&
�n�U�g�9��N.LSwƘÆ;eJ�-�;T�a	�����Z�=.��s���S�29J�����l��%G�S�'D���D	V>7K�S���V��-z5.�>�v�+*�@��-S�#�A�	[Ɉ>�e$�g�|z *Yd��&F|�~cc��b�<�&�1��G��!�г��eqEb�7u���S@����t�#����}(J�^=�Fv"��NE�n?��a��K�Ie:���dɩ��Z�a��
��s�O�C{��_�jO��l��]wg1���S۬�w&	:�̅�$�x2����!�-.�Q���M�ADTS:�l?���L4��p�x*G(rK��<��ɮ�U�MB�S"$H�Ŀ�Y�7^����i4ia׸��f��zM=�x�4TNф�o?���}�\�L��j�C������=�x�,�)���ØI�&�`����B�H���\�T���ư�w�t�*~
��P\�\�t���Ҋ�5i�@��c�3I��ؑ$i|�Ÿ������"�'G�i�N��kU3!��ٶ���c���%�3�~[x9̥T�,Z�弤�"]�0�Gӓ{7G�/Wpu�h+��})_��x'U���d)y�/��9��kE���0�ҵ�.�~�g>�������u�6����G%[M�C�7p���xuLfPX�*�7B���Tb����e#Ͼ^��!�����n6'�d���{&�@�X�b��&�s-����W��j5V;�H�8����`;�h٢�L�2Op�2F4�' 2Z���'��H�qˋ��s�������{��&&�6�~��.�O%4�L.�QP4kMF�ڄ�d{(���
���57݊y_�U=�b̪I_CS�`���H#���i���ˉ��L37[��U<J��.��V6�1��,�ғ��b�*��8����4>�?;�A7o�\�L_�c`ؿ"�0�� \4������H�Z��zt@rs�� �R~����,7�`��ZE�L{�R��&��:Jc%:y5�h�-G�����a��v�h���䋣{�& ������T]p��.��"NFШ�QK��*z��QuE���������p{������p�ԕ�̕�
ci��naT_�V�MY��\�2������8��>vG3�u���MB��L��]B�%]�l�rx�ן��d8��>�E��'�����D[[u`���)���C%���uӪ��c>�-8��C%
��⢭qj�^�Vh۲�'e/M� 2湏Σ���wɄс�@ͻ)��_滘2��w��o��<���Ƞ���񯊊c��(�y�p�?���7��qC���xDK���xjϷe��&���*C���t
%7��TW�ɞ�,��K³����g�f���EB�I�_��f�p��W������ ���[#��a�n'LMQ�a;�kf�'Ti���xW��fr�2�u}a��f�0��v&SIӗ�X)$�8���QHX:{�x r��,�X���2�Xx��q�˄KÞ��V\ h|���D�Y����eU���N��Q�8 ���'ٞ��xF��*��zO-&�H�L�cB8�̆Z^λ|~�Z�]��O��$�v
��<Ro�$�nzx!7�fD�Ɗă�N�j����oԉ/����ǁ{cl�
���Nw�<��ߢ)x��?�1{�Ӳ���b����Wqq]���%w���;��P>�lR�������l��v�S%'�p}��I�p�dh�k�^��V���`9 �bD����~\c-3��\�l�\�AC!�5J�>�F1v3�9E�n����>�>.]��vg��^�0Z�v�������em��Q����P���w���v㵱������4-��g��U(Z�Y�q*�G����.�+����x�i/�<���o�!0=���! y�?p�дlj0��x+��/�u�<���m�Ճ�o��]�al�EK���gKs-��):��C��8��������r��%�[̣t�(�L��ö��b��o�ܴ�(��75k�4��0�*�
��K�P,&�{̘8>0� �L����;�EF�����s����6;2W���57�ȫ^�G��� �|�]�s����p%�D{��7�yam�f�!O�,��A0mD�@�
�S�tm9'�P-��n��ދ�&m_Rڎ�֮���A5��W�.�\~�7��l�fb��LW��"�ߴ��`�B���X����k;G	�+�[9�	a�7�Z����aX$��g~�!k���|�"|2�H�����\jh��5� /���(k�h��u�&�`__IU��t(�lpL���2m-��{22;p2`���A�;��?�o����=,P/2'��͙f	�.�/�,qXI��f
�a�n��'n���;x|����/���XжM�=%�$E�����0��U���r,ޟ��O_z�aM���SΥ�r���Tw<�P�:��N�s�6
fZq�B�E>��g\�����)ّ�L`4i5K�>ZFg�}Y�a�g��6E\���EH�6����`�"bN0)Ptt����0a��?����R��C���Az����>�o&)�,Уe��#L�8�{~�9�(������	�w;	)~\�,�ƽ�f۷�(A)l�C
��<�g]�^*�Љ�-�T�b@g56vי�)��2ɩӹ�����[��MN!�R�� x�%�s��#�X��ɹ����LH�Rz7��������V��s�l${4I��.[b�� �X�O� R��Z(*hZ{���G�p��[�?^�[��&�;�W���Km���<2~�ۦZ�_-P��H�
�����5��M�E��S��A�C���X�}N�k�70s�\Tu�4�
�)��$�5X��
{��>��2��-��}Z��m�L�u����cu�W7}��cjh܂r"Ym�l��Z ���nft�5�t�"�W��<���{�F<҅�1�E��0G$��]y��I�Y���|t����^hkqa\n� ��$ 5�6��i�x��J�{R�(E~�#�n����N�Lx����{��	Sh� ���k�b�5��٬���j<}Ǎ�l�2���}u��{�㣾��2�r7��S�y�5�WA����B����D���y��I���9!ӊ2�n���_J�iyu���q���.���E��[���]���9�R��ZP��3�^�>�+���0Hٙ��7[ȡ�������ۙH�$�W[?����7�dU�^�[��̐+ﲪ�����nn���1��dvƣ0}9tr��v0�f���A����ҡX;8�p�[@�c�:�;_M���la�wχ�t�_\K=l�����0����x��;O��-�`h�ݫ���t)8��N҉!�t����O':@�5�e��u�D���,�"��B��������v�����/N�FE�[{9��s�a*,{"cU��K^/�����;��M�d���Fz1f:�%G?Y���(��R����S"e��Y�`���kt�q^��#�-�/Wn1{ÊJ���Lb� Gw/�E�����p:q�E����1\��Ӽ�TT�9�݇��]��g���m�9�)�F����ԚOLz�',<"6���G��<Z�7��xIU�1�x���7�S,�"Q��.��9`3A�ep��&�:�tЫؽ�r���<�[p�u���vf6�3�q+�:�`K�a(��J@*\�;5ԟ>���=��W�N�c��*	�
r�i؇%�wX�zx�:�#m��u����'���Azz�A��_�n^7@���g&/D��Nu��8}�S��ˡ�#�&6�n]Y�������!r/�_����Y�yQ1�27�528���F�B�b��܈�-�,X.��䲶Y���Gn^����ī�?u (;�12�P#Ž�P1�w�[�/Iΐ�*���u�A1%� -�D�V���x�#�hr�?W>�ZII-~��e�Z_����^���k:�����w��A䤨�Y�B#�i�d��ȉ������-f�|�׷?�3��9��T��}1S����Ni��ja��Hё��ނ�&	�<���Jί�\ܩ�����f0UB�|
sl�+3����ٌPfB� k��'�N{��n�61��u�N�xV$��őu�b��X2u��ɷY|�&oK���h�Im	���D|�+M��"����M���
�� �2Dy~N-���w���!MgI���A�*
�rR�(����xL����a�v�5[���s��9}�m�S�O|�\z��j9����5��)��p��2�ҝ���NaG^y�^�[��Ν�m�^9�&k��M▖Y���-�~�ȥ�}50���[�##���@�e�"%S{P�'�s� 8"ğ��ɶL�
O�
7vz���h?1�r]�Oxg�~1jk���Yx4��8I�Ԡ��|~<�>(-�tt"t�����N���6M;��+ n�5JZ.mdD<��di�|J|�wx4���$�^��纠E�9�e�ހ.�C�-�X�X���O�g���Wq;�O�e̘0�S5���h�<�k���ij	M��[z4�sc֬�n�܁��n����ge��#�,�t#���
����u�c[��&��v��J�58v��E�%g7������8&:I��m{�`�1#tb��ҀD�� F�*�l@":	��Ħt��@�)9�N]�+���X�C)�ׅ>���h=B�F�x��\�]���\y���G9��9{Mμa5C<:��s�GD���ԇ*�3Gk�7ԓ����ӳޭ���&��/�}�9 ^Bxц�u�o�����F��d��`oΩXw7���G767B�rU_N������Y�y$S�b!\�?�}uEZ�%��y�3��T$�q���-�ƫvx��\��b�rӧ���,m<�� �eh����"� ����tD]l��o>4��+6�q�&v
R�6g�R��S�X���a�'���?�Y�y����Y�t�N�ŵL�R��}L�uv�dP��7���
���g�����ܥ9��c��ʵ�Bf.<�w��t��t��>�Ϙ�����^ukZ�Hw�ҧɭ[�8�Y;4��ђM-,��O��â�%˃yr���Vwu� ӣV�nJ8z�V&��sLa�f�N����դ1�4��&%��|�r��#����D�$9md�lx�ݗ��hR��#�M;�O'a��$�z�O�;�k���n�{W�IaХ���"����nWڵ�Aq*8Vr:~�zݟy�U�Km�H�0s�V�+��
�7���\c6nu�f�<
��GO��1��LƸrT�w��P�[b7i�{RA��~�l)q�
�=p��ހ�
l����V��U�P(���ɢ����}۹�F*����FNn�˗�r����f�T+�x�FL����F�J2��X�3	JA�� Zq��3�I�_Ǥ�n�^C7�3�i�9J��{�
��.χ��%6@�����"pϠ~BU��[AN��z�rjV,G�0�H�@��/��V�s+�l��_��(��/Ej�`�'�&�������u�!_%�hK�i����`;-g���Ԁ'?�_�y���ƄM]��<}�<
sR������'�b;��Gg�UJ�.��
c� Y�X� Q6qVq����vJ(ә�_|����������8v*�����c��j�8������֯�S}@�c�X��ځ��:~��1��J�Z�7�H��oh�2�M>Q�oK���a�
��)r���b�r���3/޾n$k����R^�X�Sp�q� ��5U1��!�{M~�q���(%!��f��~��D5qeX�Z����`%�S�����av��R<K]W�T %Ґ#�j��_Jc`���=E�BQ�f���L%�qu�^s�Ľ��.7��\�n)��z�D�8�rc����lѶ��q��Ͼ��;D��NΒ�Rh]�x|!Y9�I3�.\�Q�F���b��_AÆBo GDNT�H�2[l�_/Ɵ�?�g�@��_=;*%���v��G�8NFc��68{�!�D��3N�)�N��'9{h0r�^�J�c19,�QM�FI�-�A�9B���po������aZ�K}�}���}]3��R|���.�֜�c�9��V��+���G4�u�h��gU�BM�-�cϵ�O)�6�hs�Z�M���U$��_*�O�>b����;!����g�t�NP8y�t�"�S�4�*��eU���
�v�pR�߹׸ �4X7�Ț���C�t}��l�ԍ���a��W �:�k��u�ğ/����y�=D����]���3��B�S�[�NG�yI|��j��K�GQ��,�,���g�!����\����9�۶�ue�ag*pV�+:��q����\���������!{�"jG�Bs�����[�H�P�nYt9�*��k��vR�����i�XػV�geͦ@Ό��n��d��P�P�7����&;��F6�>��!�w"���.OM�ˀ�����4�2+���;l9�I0���Ÿz��?9ڴb��t^	�d_�*3�i	�$�]'T�Z�詪2�4����ʆ���F<G��&��s��T3S��pr-�C�d��Tt8/����^�2�(��$��6#���?!�u8��?EՖ �:r�����y� ����]�d	S�2x��n7�3g��m�E������*fQ�����XݕP��hҪ�����m_�p$2�t��`�(��U-=��U��*?�ϟ�Ap� ����.3��$qNB3t�o
g�'ò��&V3�Y˞�H��K@:����Mi�\��-"�W��H�c�%����{
����*�;��ؓ4v��,�񽿲��;TygGb	W��T�	m%����� 1U=k����ҭ�G6��R��yoV��v"��Z+S�dRƾ/㻘?K�Gjy�t?n#�\�(yx�"��m7�+Cݾ�*�!Wz*������#"��Ś��88 tTQ{89�\r�n���#�� ��D�n6F�&�0�ٺ:�6�p���Y�9Z��<�m���HG�b90>ڨ�&�ԗ˙�,�a��$ ])��e�Uh)YW���59	A ��m��Ӽ��o<�Lj1��	ď_��]��$�͔��'��lv����� �@��傈DGu��Hd0:�;V��jW\u.�wT�`B�W©c�Ϲ������d��hoW��OY�A�/�DO����$�!7���_>�#]�a�,_<	������I[�A��p.W)���PT��
��7\ݐ$q���S��I>-��m+@��w�Fb���B#��6������s��V�h��|�fZ� u<�YJ1ߎ�T_o�J�c>krH2z/��'*ɯ�b_܊�o�$詻%s��=�(��h��;Q�D\�S[�ؽF���gwK����w�᜴�"n���/�S��t���Ll�l�|m0z��'����!�U(M����,2[� ��!�.X��G�v� ��>����.�{3*���g���7#5cwq	����d�$��ԟI���C$czK�`Ԧ��k\�'n\����8�?��J/୼R��z�a~n���[���4�C��&S{�h@C���;A��Nڻ��$}a�-&��>T��.Ʊ����E�饈�pKJ��I^�],�W_�3@�"�C�Xz�D'�a��Z¢
���c4��[:�Og�����s=yW�P��j�0�9Rz�ر�1���-3�ئq?:�fd��x�@7�����Nk.��S8ɆL��wlVP�H�
m���i�K+��[�����֖r�	!Ŭ)ߕ/��0���?pK�ϗ`Qp���Iq��OJ�x"���X���5��5A��s!��{�3����
B)p0���V	>&��u����>��ƛ0`dy�w���,���A����A,�Y*��ɣ�\�[�� ���T�L������~�2W��ܿ3�������*���(�u�q/����ˢ�r禞����wѭE��W~�2nb�?�5���gG�f*���j���J�n���,1Au�'x?D9�#^`gJ����+T�6�P�z����Kq��|��_�}�A�M���*���Ӥ����$U*Z�N��$z���$�Zx�UՃc%�f.q��p�q�oMʕ�.�i0�\�S�I�7F��Yƍه�x�ϾOEփa+�
\̭YC�`�|z^���S&��=	�=l���Ba��:7b>7˽@���J�K'�Yo����ö��bi�5,��U�FBb�6�6�҄�f��H�O�^�e\0|�A�!$�Y���#u`:�P��z5�Y��p��4�4�xh@��d���֧)-���s���F�C����{�$A4V/Ҡ��t�)5��2�"��R��.i��'��ԥ�����_��Ac�?Oð�N�Q֊�Uo�$t��l�D[�8W2	�3�o�-��-@~&�y���t�t
k�L�~=ők������ذ[��
���Z(@E�3W�~�-2����1��!|���t�(�n3I�u�lͣΔ�.U[ƛpC�e�8��
	��Y]��}Yڐ���g�`�?�V������J�c�'զ�b8~�K�-/�������4�Wc��qV=���t����Ψ�Q��N�Ys��{���J[s`l�u9�	[	+)���1~����2M	(�G{$LM��~���%u��pۈ��eH]�Iʊ���D�C'=��î�I�J�RC1���O��O��ς�����������(���f%�:rYV=�H�\�^�)9��嶋Z�ߟ�U?�����#m֔��[�l��!�ޙ���{S��<ϋL	W<�"�_�^Ge|�O����rw�+�\c�T���![K�7��I�M����_�r����>Ħ�$F��p4��7�o���VX��\��[��[�['��\�`Y�
fD=��� �h��8@m�<�JN�9�T�t���^�\�/��R��삣�(bv�q@�w���y�K�`F)ͻ�՝{�e�"��P�E5Ӷ�� W{�t�vS� ���r�Z�D��$?��C���f���=ۣ����f�ս0�dݪ�C��,��Y�"c=����;;��U��5�8iW��ҡ3wW��M��<����m,���e��[Ϣ8F]s��c��VD�'P�6m���#���,����!��nԩrj#�[�L�s��f�W�m���We� �t$�N���јS"�
wҏ!S�G,.���e���H���>���&�0ѳ�*�(;��]W��+��Z;*J6ߝ�T��ܼ��C�"f� ��v�22c%J�C'P��I�X�k ��{���n6:��'<s�x�u�v�IZ��ɹ'���B���3��F�ܓ�]:���X��!�^��kѧV(�7��,4��%<�B��/�P��vp43��
2�{�sY�>w)��Qڥ%-�U���X-���;��ȁ���JPm����K�p C��z��R�G�I�
�8�"�#��s@����`�=*�'�XA�46eي�7����F�!���	-����
����9�`��f���fs�焰o�f>u<�_�~��3!�{H���	qs;�.L��B�UU1�[�5�!y�m�	�\��� (�2�.@�o�r��=��@��nV�D������d��kW%J�����MoG�'S+|�� ��&��,�c�c�/sY����X�~*e��8�m�=%���o-��4����J�K�����s��e 9�kM���M���"3��Ao�<�����¼�хf�o�	q*9-d����l�A0?�\;"eٱG�+ܗ�������$K��9�N`c�����\��0�$�=ye��'�G���RŁv4�_}ž��"�}Jj�k��%���ەʜ5�*�A�NsQ�Sڃ�y�a���"D���)V�5v����ͭ��𤨁� Y�P�����2�E��g�։��=��j�K~i���6E��5�rJ8euձ8w�s+O!ƕ��-�t��>\-��N�@ ��D��-;��G��푕�hNkT�tM)���08���S�0hj��*�ՙ�L�����@���hh��5�>�'3&W��}^?�V�:�#�W);8X�&��oH�و��o��'Щ�`�ѿ�B=9�D�x%u��mo�&D-e�,h��O��Ճ#�߁�5{��3���,�
�2�	|�q��;�3�uZe�[�^���d���Ǌ��	���.$vY[�xn�a�7���W�g_9�]Ϯ̒�F�ܾ���a���$a����q[�YzX-��H��N�Sv�8NI�Ja��1y��� �#�͒ͅFǳ[�ep�J�dF����jgھ���B9��~�U�dc�NO�Aƕ��6h��[���RB��Oܣ���'��gR���V�6̈́n�tX�����%����J���9���d��B~-B+�@�W���I�����3$�M4@Z����N)��\���Ei\�'ނ^Y�߫NQ^������X ���]�������7�V�F]�S���v,�Ȩ�`�K:�EQOc T,������P�Y�hE'̜�aW<��F���Ti����}��:��N�pBH�r0:Mr�Qs�E�?�4��gsv �aP�AV_@��-p@-ˠ�6"�>�������׎r�F���i�;����x�ӛ]�\_��b�Ƒ���K�O�O���M�u=V���0X�������|���@t���@Ǒ�o���{����W��,e�y�Q1�Ǯ�܀�rv����h��r�T��+
�����z\e�d(	�7*o�t��󰣽qc\�=ḱ��Ft\����{o�3�wԟ�E<�����
@������S$��d��Ӡ�>R���D����-]�s�Oֹ
?��x�}ll$玼JY�k��y4@ ���q���#=���i2���,r|���Ţ�%�T�d\-�(��?�G�B��#D���v��8*�Y�h�ӕ�'nn$�w��D�p�:�
��(<��7�A�=L�lVm���'hq���9O��Đ�1��Ɵ���+76��4�R#�eG@wE��e?N��g�b�nЌ͹��ܶ���gP��>.��w?#������B�Λ�;�tNuF�4b��3�b1���evM냯q�鷛@�� �s��=�-7�]��Qlc��VSf�<��#��TQ~���]A��x�LV���W+�R(9޳���k���P3��ﷶ|�&�@��)�����PM�X���e���x�ƴ��	�����q����Z>!���/\ ���vy���C�I�a{ ���2�Ͱ�?�4�����U,�|t��/�^RF�!'ҁ C��t}r�Y�WS6@�o�-o�S�jpG8���1�yš�l	�x�L�ɬO�6E��:�"r� "�(�θ�/y�v�4�Q� N8�\yg�����?n-�a���|>�����wT	َܸ���0��d}�T�	�����3����X��q��록�'������82f*�������'��U��T/m�2��u�F�XԨm��<��!���z�y���>e��S'��8zw83%Z/�O��N,�h�W�?zSa���mpk4�Ub�+������T��Z��H6k9������Î�+%Zh7M.J${������an���nb��C�K�t�x�\��C��m҅p���M�xJ࿂���ò��k�2/�=<�*�i7�NE*,E؇�B��($I�.*�\�MQ��R6Z?�ە D�����r�\��S�<|���I�b��.�mG-�>&+��Э�*�*v�]��T�G�����}
G�U�Q�O�$'�@���:�d1B���с!eɔ�[D�A���RnH��%_^9�j�.E�T�����,���G0�L܆[���B �$��@n���T<�爤:%#����~W㧎�-L�U���}&��^[����h���H���q�0����P�����i��f;@������d��*)����H�1Y%
W�>���.Ö���T1�`<��+���#^4�7;E�D����T(Ux�y|�G�-?�8�� �@���{�J!��#�W�ʿ��)=�D�HM�s�D8�d��؉x.�S�����B�,������~��
�h���BÆ��k9s�(ɣ�F<� �$H���.o��Ӗ���9���c���G\g�tv0���� �؆��B� ~m���eCӷ� D��f�JP2���L 6��s֧��`g��ǌj��0i�п<�&�~� �*=w1�Ng�Z���u^M��ǆ.3��|&
�j�R��S`PGA�����c��qMGQ��MJ��kb�|2������Ӕ�iŉr��Z���7C��?�R�S���6:��7�/^ܐ<��e�3��2����~-����g��v�O݊�(�&I p�%g-0��ڡ�F��b !-r`w��}#q0qGBh_�l��Þg1����02Gj'#y����E�LI�]u�������6�]VÅ"U5�p��jwP�3�R�=�nx릏p�g�����q�;��|	{�gjŲw���F ���A|e`F툰�(ɥ��`q~�d�t��iZ0KNR�}�Dv<��Ȓ���2�	 	w��Z��r�����kʏ�Y�������`�{��� �	cCV1_b�ǄqZ�������V�wQ�$���]����R�d+!������:��q��ڤ�0آn�o��c���a�[T�$��´Ia/�W��Aq�(�9��~�V��������{��i];D��y/��@ܪ�/s��ԇ|�� k�>���=�pҳ�_椡���и_=`��t"V�9��&�T���'@	�)��q�#^�m�(�۵�9�f	��yg��?�{N;�~Y�� �c�U��cIa���#�����3
`�����5��bL�̌v@���J[�L����'.�[gK�I�%�bgP�H��z�Z�}桐�AkJߏ���
Sj7��m��'2�fy��]I<�˗��U��F|@��d��-aD���zJ>,H�o�JT>kh:�#0RT�0���eQR�9�?�9�Đ"���;�ٓ�M���Y������G�tqa�g4��V���x�s4�鳥G[��^�s�E]����ڢZ��7H����[���ÿ_+~�щM������g��e��T��+>Da]�SJ����!�mF��n�:b�h+b����}�[�a6ޛA/�EWx��ckT��N��
<^j��X��ћyJ3��N�DN�@&�?H��W}lu�ù(g��Ӎ2��8P���<��t�]Z�(̿#T�	����x��s��q�w����Eo
�E���>���a�_�!5�tI�����U�R��'�ԅ�#޿����,
#���<Ҵ��BUUJ���<i:�����T�p�<��.0���m���b3�^����~Q1<M���k��W��ҳ��m��)�#Ga�T`@��p&���j�۽4�@�90i{��g�~,�|;{H��i��=w7i�n���61F@���$���'����#�vZ�:|t})�����cox�]��~FV����x��ՙ��]+"%c C�Zd� ���k�)@8����pD[��L�DA�<`.K��`�����@4���(����V&:��61p��r���� �vZ�0���M��iI?�+v[���rW��NE��
�kj�}�����X�P������5'^r��e��*��L��~��.J*g?P0]�[��1(Þ}s��ըm��,2&�ŕ	��tyБ�$u'A�?m�~� ���gʳ�be���]s������w�ᭊ��d�%V�$]��/\u���WCf�c��?�"�#����U��ږ'٧�w��ǯ'��?��A8e��d]�l��I��t*w��Okv���+�G��	���dF�<�''���u;�Tri(s^�CXub0Z��!@o�a�=%#��ӴU)u�������ź�D�*��i�[E C �'Tg1]�;�f�&wA���`��,��Evy!cL�%k�
Sf��{Y�V�����=ܢ��b��:��� 3�N�\7�a,�D�{��畬��UN�0'����Is>K�0�*f��t�)S��i�7H/��D��y�3aŦ��t2� ۙ2lh �df����R.�id]3���v~���q8��q�"�����/��R���L�8�u�$��'���`~��ԔQ�QYQ�%�E|} -q��4��D""s0���x%��z�>�T�)�B��2���Qyfˇ����:�M��b=�����p�5��܉c.��vT�R�>b�:Isoѵ��.��
a���s�G'����ʠ������v=�v/�f1�>1�
��X�2.v�b{�Swp�X�Hy%���ۥ�g�V�ʥ����������(�k���b�wn�H��@�_͕v���6C�)�Nk��;Gk��=qԒ�����U$�Bz3T���w*l��O�������mt���;��3:J#UR�G�#�����,B�4Q%�t��/-�pc$��!�z�����P�����L?LQtyJ�G߄-u\�²TU���C/��"7�b��Q��
\�y9m�G՜�!��Z1XG9>;��i��b�9\�P�|~����ַS�K9�����Zf&�\�d�LR�v�B�ۙDº���9/x'��w��k
�������7	6O�����'�D�B�.wC=��O)�b�FoO*j�g�F�$�;ϰ�����!C�� �P�+E��e+yr}�çVEII�סrG�h���=��j!#[�b'��ǰ�)d�u�x�լ}�g�ou0��J�.���%�W?�=W����]H�p��&����RTW!9��t��8��
�%�qC����V��}��sT�0��O?�p33�a�+�j�l�xj�V�m�m`�DO��O��G٨W�؇Q�Q�?�����%�O��5�W�k���a���tOW^�u�B�J�D�}�X{��Ie���b��N�8:���!�,4F��;���T�'H�(��B"b�K�HJ�{�|�\\���h��"�u<Q�1����2�2��0���u/��ě�ޠ�pA�_V�oϸ��yM��.JT=&ԺZ��k�,�u�
^P�C>����L���G�Ҹ�
�6��P��(���VS�뚸�c*L�_�\<�|�⣶	��,�9Q���V7���,��)N�d孿�[�h�ɪ�{�'�H�����>�Uf)���5%��|���_�"�V)�M���˪�`͇k���p�=��Ō!��Oca]Fv0��hj�\4Z��=�F����}����`�Z�h��<�Z�U V��q����^�=Pd{�K�����x8�����ç*����:�x���x9�A��*7���)8+�R��Jɐ���8I_A�f��vhN&��F���P�n��&�x�v9��Egm5#�������SJ��w<_��+�y���@-�th0��{��3��Nrj���_�~�`��J��Q�)��<g8�g�B5%��SͿ=��]y�0j��#��/�PFҠ��)ˑ�u��V,��1������.�ڗNw+z���m+�X@�WVv�۫�,S�A��O���\����,�H���4��5_(�.��/�19�A�K�3��5$Hw�F�C'�;6�p|�@Z҄�0r8��5�r�1~���+-.~7��;�8�4*G?y<0y���X�rH�dI����[X6�B'�}�wXߒ9?�����	F�W�n@�	��H��J���!ʭ�J�7��D�&�qWo��W��ϕ��be�gAp��b����[��y��b��]rYw��Z�e{ሁ�p�w�a)7���|���Ҝ-yf��'� �V�2��b��p5sI�S���ڿp_���~���G�i��)�d�tG�h��I^����ip/n�J?�RVBsc�v���S�"�#�<��g��I���쥆�����"l���Уk�Qt);}�v��ν�	�M_:|J� k�uv����w	Z��ܓ��QP�����z��~�OĆ�Q�l����?jC�z��ҫ����2᪽W8<�<^K�0Q��5�12�N�}s��tw�P��Bx�ӌ�u�� 6�L�He�ӂ��w�+;QaY|��
l�WS�!?t� �m1Y�N
����E��5(��/X�L\>kw�x4=�h�e�	u�վ��aE�1�Ƀ-*?�t��_���0N½]������Gz�3��J�:�V���z�錼���-2�"�55���;BHOЉ���W�� ��z�T�5p;��@����pI�Ͷ�f����s��$#�T�ɾe�� y��:�؜����˧��^0��t�7;M���&��=(Y��h�V8�{`�uΠ�9��Q��J;��T����D�����?�����] �vlfgi��������]ώ1�r���᫺��Rˍ�{l<@c���3�rR��[#LҌ���@G�BW��e�(��04�&3���q��� ��/j�_i �4��;�
;w�.�,=�,`H\���<^�=8���z�Vb�[t���N"=��|?[�8GZJs��4P@������QI[�F[#�~ �Ǝ�$c�^�p��"��2����B�.˻K2��j���?�BC;�>�`�K^���S��D��ᄼ��>��pD�M� @�A��	*�d�e�6��O<ƪ���s\��g�գ���'������<-�J�j �Un�Fȑ
�ٛh#_̏X4J
�����(!5�1BZ����c=�z/v`-��UL�R"t�����P8��1r�dh�N�:��`�n4��s��݄ M��C�OF)gg���U�R�S��$ee�8�aW�/��%�/�h_�d��m����������W[�}�TG3>8��K�z�K�w
DX� �f;�2�9��"��j��O%��8F
.�)���XИ�s!�G;w1/b��јϢ')k���^��S��D1�ʆS���
g�z�ق3�yEu�:"!���F6�p/X8~�6���A`��^�^�}m�����Y�!��Y_���˩-��F��`�uu�?;���A�#��IH΁�&�oN䲭��.�f�7��вַ�߼{h_k��J|�r�0�}t�ެ�%�O�Bѐ��brde��2��.�s�������I�T�V���������O�Lޡk���#i�L<|��"_I�u!q� Zgk���B� E�?��V��1�?s�~\�_([xk�"�<z�2��=��z�jW�&����~�<_.�,~��V�
x���.B�����|�?"f��4X�uy�����G p�QMґ���;R�q��#��â�\բ3Mx'��Pl-��Ɏ3��ʝ;��� �9�&��T'��.�ȋp��t�X{�������Ri3���I��O����.���ߺm��R�^�R��&���s������Rc��y��k�ķh�:�����N$ڹ���ʋ��b��"z2GX�'�E
�$Cl'U��$��=qe�gv�BV����x	�a�>~-([�J��
���~�G`�-�j�?]H��]��ش[J��������n�D�2
�5=$�Z�|��7�� I���㯶���J������C�
m`���[�c�\�2�<8�O�X����������Au����#*�*4���%"�7b"<=�.��@�$�ѝ��)��n��G&n����Á���W{���P��6qQ_��߿=���V�D�d����Q_��ß���d$���Q9m�g���f���Ў��g9�#l����O�U;ؓ�Iut9�b�.1.�Cۏг{��}S;�$��#�e� �b'�g���.�̓&IN�{���wQ���My��U�yv^�&�9� `�"�/fb��&<�K��rپ{lP�ͤ�gҒ*��1j��Ք����	Bs|���M1�$1��Bi1>�{M�����#�G�W&lf�1�{<��G�%�1W�7&Ied���JiN�a�n�Q� ���÷ͱ����U[��5ku�{U���w��JP�ʙ�z�4�S�BKl�K���Hx��ư%?��-6�eq����M B_vb5���p�W�����i�w��i�^����������I��Q��u���Le�AG�N��oYx��_�QH*��Zw�(�PMdC�j"�L�-��c�乪�$�CMiŨ����m�Ǥ=gdT���	Ry<ݎ����<r�X9wδc�x�ţ/9ŏm)�KT�|������@`�lS�����1NV�P�H�e,��y$��A�dP��U~�7�����Y"4��U�-�î��U�&� �L����d��v8�c�l�_m.����3�R�ƣ@R��p��P���ᔥd�Τ��� !�2[�@g��ـ�#G���+,�^rI��+Y����[����Q#i��@����ߛ��Ӣ'XK�v����h��$v���ѵ����&g} !��D��{�([B�3�{�oL�CY���雳�;6x�NX�n�z8�l����P��bH�J���7�}[S��������J�ꒀ1c�cK�U��D���B��֐αXԫ��SE�s=��@�ns���<%��.�j�{�#;R��\��������{��$��@������B�iё5BA2��В�
�����=3l�G���%v#P��~m�� }�`�h��8�^C�Y�(�JJt��3h� �/Cw��šO��V����v�K�h������v�w˥�L�q�f�_�)	׷��� �_��^�1i�~D(���� �^����?Jd��'qt��H�Ɩ����MѧG�{:���Z�/Yϐq��^?C����l[iAk4��P ����2�Ԃ�h�c��#JEG�����ҕ�5�+h�C|T~ԇ��q�Qě�����S.��E���n)᷋�6>�'�N�j�H����BA�20zK>toiWvk�[�Y���1������yL�*��������&�R�]x`�WvO
��al樃0z���wq��[,�L]�K�������k,���> ��F>�O�����UC"��h�Ǵ�	?���o��!�[)��m�N&e.������+0e�����V����wo���߿@�ӓM=�����'U�b�(WaĮ�V�4K�ա0��\j��g��r���M��7do{$^ats�9�S������F�{׼��tG��>���٣��#�keGX��/RB.�%݂��j"~F��3�0F3�&�vضDD�=����j@B���V	��..oM£B��[���nNJ��x��f{�S��	Oh^�wu+հ�|_��Q���}�X�T�j�߃9���!��>3e�9k��W�(g��{�hH��u�|�&�F`E��?�j�1�,捉V��yo���)��wn�U	RPө�c��/�P�yDTr���5��9C��r����"r�O�>�3�!��t�l%���xr+�_*-���r��:��A�O2�i�A�S���YVռt�ēI��5U<C	�qs�0�)�^����z�%�Y(l�q��X�!��*ͺˇ��{
�d�$X^�J�9mP�*�h�Nr�$Z&`[\�v�m��Ap��X��̀�,I��k'���A=�:��ir� o-H�����\���<(���N{z�:��~���s�d*"��DJ��#����4��]�(��TP*zt'B��H�m[���f�R�s_.G0��=��S`ⶑ|���f^o�Ԧ���>&�nk}��jPH5�|=��c�~)�i@���$Il���g��X� Jc�d�}<�@M����Ȟ�p��Zp"n:W"E	�g>=�]�r�%�!˦���e���������4��9�D��o*�I�k���&ܮ����t�\��.V�}����ގR�L}R�)핱�*��9�)�"I ��p/ԣ��3ĥ��9�dv ������L�T�n��#؀r����.HG�*r���^���cb���<���C�D��d3M��K8k��P����j+�y�w�Y���9a��N�׍�d)��׈��}�U�b�%��xj<7���;;ݎ讀��%�әf�
�����cL���2˰����n
�,_�똟7;2�KF��ҿ�ܤ̲�%��O�!n��sϬ4o=s~7Ӌ���el`�Ѩ�
cһt��t�^5��Dڅ��))���E�6_	;x.�z��->D�=��`&�c#a9��M!̺�����Zj;���z,���r���Ѿ�h��p	���Z�r�w0�	`p �Y�.�n:�������5%3��O��ܑ�Nȱ_n�����N�]Ȫ)5�p��=�i�?�c���0�����+��bZ>N%ٍ�"��Vl�Z��L�pS�j��Pv���'��MPP��2����#V�4H����xL�j��aRV�w[���M1�~�R��o�&��;��f���3э�#*�K�C<�˪1���J�X����>!-������ٝ�w�	k�t�j 7>{!(�Ÿ[g%k���g���[v	<q�=��؞����7�?�k�D5.�e�~g}7: ��'B�<43� \-
G��4��+p���:C`�gl~��eaHC�wYbC�j�=
�)0�iF�`3c�o]��3*��M�L�B�=�f?��k�Q���nJ�Qi�@�F���SF�ܴh9��u$׃HCt�ר|�ۀE7���u�^�@
y�f��Ƅ�ջd�gxŋ��G��O�3��8���������g6ȲP�x��=%������4�&��ɪ��/a_,���4����!��Rz�}����b�T'�������e~c�%��?�ٵ5�Z��2>�ZZ�'�զ�)D{�Ŝ˟.G���'�H��J��t�����h�\:4���$g�:�g�8?��?Έjw���vl2�#WbF:��-��^�%_5�G+���W������*����)U��5��w=���j�����E@��أ1i��[N�=��vw�����r�Hb�J��G��kmE ��J��eV#E������� I7���b_�M�����Y��k�dM.��{�N�j�B�}��]?iIؑ�@�YӾ�d�cF�(ëp�ݵ�|�߭�6�e�H�$�,��!�ǣ�?�A�`��V#V7�Aa����/��q���)����L�!ƹ!�����-���U��q�Z
%9��)�$L�R�]�K���3,D�0&/>�a�2}��𼓆F��]w�?Թ)j�A{�+'�vj�՛7c���Xg���oly������h{6/5�10� ���#i��L�Qpd�w�.*� �*N�Ӄ��P��V.{�%��S���]��~a�:�������Rk�^F�bD��5=��:W�٧0��
P"8�H��N�a[���_?5�_����?�C�lWƢ�#אYj�~��ԓ�3�b�����ư����SP[��_�p�m,5Rź(o	z�m�=���}�k���b�r����ߴ�5�}�v:�كǊC����8�=N�H�˄�*�<�!$6X�Z� d2|��EF��<޷z��,���q���� .�9�^�ob�^xG�^f���L�yWח$ehM��ʹ�'#�+����:�7��5��gE�d����G���~Z�D�����`��*�2���Z�#�������@��Vʭ�l'~?W�b���{�{!��[M�Π�R�g�öaL��#�~<�����|`��[΅gmPz20���&��Ή��N/�m�e�0橒��D荧3�<�e�@��C}a\?��cG�4�|�9�Y]�����O��&]��@����Ƒ�=�)��<�D���x�2�����Dr2F���0�F��µ�&���d�;��p�'b��ϻ�*�*-��ݳ�.AxLOｹ�=;����M�XQiv5��C:Qy�|�γ�o�M��u7`͢�b-��3�K�t^�{�DHӼ -�d�2��V��>x
9�킙�T�����
"}sG����Ѓ �L�U >C�4ͤ�����:�~ƭz���zku(�;�胷�*��@�s־p��Viƞ�S|�3�X~�^��O�"��I�2G�oH0҃��9z�:���!'��=�V)�赪��5�V��8�rڶ������E}o�fd:J�J�S��LW�0�)�c�L,+5�m��"1w|Tg�h��x�)�
)�v�`8Vq t�7�zZH�K�4̪,j�z�5�2|���ɭ��Pu�)ذTn��F��e�(_�2��T��i��o[�(�����E��B����Q�Σdt���(l`<S r����Ģ�D�C�#-��e�G.>ɿd!<.DyM
�e1���9ק�@Ux�l����H^�b/�T%��w1�Q�Lu�Q���ٟ�o�E:�	��鈇؟�E7ް��$�$�;~��p.��28���9h�5 K6�Y<TV'D�L��F�^(kw˸�����lS����xۡ}�[sh��������䕟���ڝ����ۘX���C��r/��n}��5�um���$c�q��qbS���g�b�ٞ��Y�r<���G2\�l8q/� �'�.���8�aG���RTP��㱋�Ss��$��o���ߺ9�>�6T�li��ܻ|ZL
��e&�,�j��2����`\"�0�8�{�T~����>�E(:�
U�Y��i��	�)���� �S;ߠ���y�"g%�PϷ$fY����۳NI�0�83^�ݴ�����Ghɂh�ɧ�/O���Ʊy{��&�S�ً��N����2	*�l�w��j#l����˶��$�����b�?����4��y�< +�R
l�f�_;��G����?"���%�+��@}�4Qo���̘	�� ���zi�P?�xk&q�}IG���@�^I����m���ِ�����-�Wa�㞁���)uv�.�۞h,��a2�}��Y&��a��/_�SE��9�T�
W2�|ϲwF�W._Ĵ��=:kf��6NAB����u�����;��Ȃf4M�P��/�'s��N���Q\�⩬��GdC)
T�FS��>g��s
���W�/;$!�i�u�u�7؆���F<�q�_6K��;�����RȌ���$��C�T4_�d�E4}h�+q��ʘ�#�!��ŋC"��4u�#��]������i�y�����΅�����Z�1�t����}ֶ��T�
>S���5�&kIk����
�#�c��`��%ˢ�K�(ܹ�%GJS�p���fMa�(7%���!b��0� 7���a	E�k���?�(�qr���1�\(�	�BF�j�\�dͽ�~]Z�$W@�/�Б���h/��HԆ�+L^� D��Zf�s�L(���S�>�%�v���1�*^"�vNM����?3�ƥ�r��>�ؔLK�#S�wF��$��&��4˻���+C�]0�T^���>���^z��⃌ܣnc<r��Z��6�Z��ǽ{�u���w�D`�ɗ�8�ˉ29��%FP�&�Qp65fK,VE����L�n��M��uR%��3a��S���ɻ�r���C]�������k�h7��"@�E[U�c�Y=,Ł�W�^M��|��[�WQ6�rEeU+Ť�{q_Z�����jI~����BC�"���բ�t�x���0ؓ�L��;�L���n갃����k�V���?���U�n��܃D�7��sS����њ4Ra�:nJ�D�Љ�8f/���������43*>�+������)ݓ��11Ď�w\݄`�'�4M�=}U��}� A��:ȭJ&|rN�Y��ِVn�
i%)'Ph�`�k3��u���L�J0����^јH�~B���Џ���Qu�2�d�G�i=H*YI��swD�!4}��6�5w�1rӎg�^o�U��ZB��ۖ%Y��!��ٹ��>UY_2��B��OH����O�G�_M�p*��#j��;�E~/y��hoD�C3y�x��EW�lHY��� =_%�=C׳-oUxÂ�i�0+A�R�ױh<j�FG�Ӕ�vZ�-m�IC�~DTj���D:1���ْpR�x&�X�1�GO�jG��&A@9U,�B�G���]�nB���sqS��C]6�^�M~>�r�@ƌK6w?	D�)g>.����x��T���/��Ǯ��|T�7�Yi����(J�[kHr:�f`�)'�Ym(8�x��&�X�π����u��{�%w��,	gK'�����D��}��%�v�ʗ�q�Ѽ";A��ή:G_F�[��g��{�u�S��(��DZ
��������2b���؁/���5��?9�Z2������oԱ�f�����ϴ�_l�,͈6��|Ӌ��'��n�E�q���;�|{���P� )�� f6�i�F���5�� ��v1�;;�^˾�*��,h�`�#T"|[�ٰ)�w�m���3R�-c�چ�ET��������>�����[�쪞Ǳ�-���:*	�h&�+Q�˚%bvq����������R �Q���|Z��IU��6�8�;��Mb�������A����ɜ�ň;-Z�%mEJQGB�������O�� �*o��U�Z�+�ב�[D��!�Ύ���IP8��v�|�I"��M먼���f�iJ?�=�j���D�a�6|�@�n���h��/�3p	�M=����[#�g��W�b�ni.�){YP�"�DV'�_yY������n����ny�c �O�Wq��˄h�7g�i�r�O�<�	5X9��ݭ�?��Hh�hs���G#��F��*�r+V�jN.9-ʭ��k�����0�?�so�)�y���>n��At�Ro44�=��2�m��CN�p�̃ͳѯiY5���2a~���\�M6�Qsk�Z���@�<Ⴤc�һ�R�{ �v�1ShP�CHۮ�#D;kI��E@@����5ɝ�Y�t���1ضo��\-�4���SPR���,]1I�5��
����l`i������D��j`��!��6^gyu�<u����Fe	��"���0�&/ʙ�ڃt�#�
�o���3
�h,?���N�R"������A�8��x*�8��L�X��}6��\G��r�@�y"�-eX8�j2oM�1�z@�\_�Af��?}@?x����f$kV0��u0��s2��ܚ=L�ߛ|�8�ʲ��tU�z�bC_$�a-)��KJl�f��l֖f>��F��uk��.���Z�B��m�#���P�Of꒻T�t�y�a`�H��U�X�r-�]�	��h(N;��fW�MuM;��b�Ls4�~@Șp�����,���׉�?nV�i�Ui��3�`~I��\)�mt���4�m�{גL�*0�	bR�"0h窱Z�|r0��E0����7dF��E��y��7r84Ncr�m��Ax�->?%��.�<k��(B!u�7��Z�TE��\l�������jA��de�$�8����2����8�Y�����5u&��<���_�J��>:��#3~�#��ä���q	�.��pxM�W�'?ڑLb�4A��б/���]�:1���՞���q�����/�k�0�0̈�y�]�|�Ȗ���V�s��=��e���vh2}�[iƏ��kl`r��Ϡ-a�I�m(��0�
����hX��GU�յV���r�7 ���\���r�j�L���9�n)�ͰҐ�phMt3 DY�pȾq�
k3sۀza-w_�=�w��љ�3e�ͮL�cO#� �����@��A,�x!�B��H�5(��Gv���k����s�}��.�#Ro���3=��/hi�P���2�W��˩�m��bY��H<�&�Vް��
r�Efm�g�B����@Ʃ�T^ɯ ��f<��D��W1�j#n��c}Z����3�R�*���o��W	�
��׭��Eұ՟��Bq��ċD(����>ŅK/�:�p�	~�_^����l�7&Xe���AA�hB`�T�N�ƚR���G3�����mb���G�|(�T
�\V��lO�6�3��fEO�oP�V�m��4#��oӞkI�l5��c�@�?@_�^;c�V��MBD��:0q�L6kV:��&�k׆�%b7^��~�F��l	3f�����F�K�G2��������t��<��l������gA[�p��_����AN0�����mEt!�_!Y��x��Ծ}�tO&�m#5ɫ�TZ�ɬ�\��[&6�im���mEj�j�r���J���{��#گ���q�Y��p!��1%�f)�A�(����&��&S�>X����6t(�\��.BθT'��ohy��8�Vxr0��%/ɬ+*LC�X~rXӶ�g�n�.W_������>*���~f>�$	�E� w
9vL�2�����Y�VT��Ҹ���Ōp��g��K�x�2�� ^9pQ%�l�����zKg�Fq����CH%����i����y��4Z�z�N���`�s%�>[�7������׋�Y�c�/j�'�"��9�%5RP��H�'&>�!����T���7�&y����7n���W��|�s
vCs���՝`
�W���A����"i
��4t�_LQ�����G�^��oM?�7�"��^C�a�;�N�|�tzG��ƌ���;Ԍ�������z�9�d�بE�T&��`�u	�ń����e)���� cF����EH�]^��* �RZbMot��I=�'q4�A/� =%�V4��;h�6�r�l�O�Jg���E���px P`W=�Kщ׷"�	51fjU$5X�W��@.��No;�u�]����?���=_�1�fz��R�`���-5��a� ��p5ALP����u�.���I����X�V�4�Z�W�7,�R������A��@��v��S�5v�v�%U-�B��/�B�56׸ ��R����p;��*
� ��~o�G�9r�C��1��R�x����m�ц0�L/wA��/�lF�?X���U���&	�
���I-��l$��n0F3�^�o��/ �g���P7��K}V��7D��+Ԥ���#mv�]E4.Շ$u���D�:�=�	�h4�V/Cv RO�mvl���f欯8�
N}�{��b/��V5���N(��-����v}nP�o�b�w
�U�chc@�ț�DY�#�Tҙ嗠Z��kXrb�G�x\RϾ9,#������$�S�(#�."Һ��y�&����Et����p(�05ծgF��3��Ӥ��PP��/<x��6O��z���CQ��ox�Z�ơ*'�K�d�AH�Vt�:��#�i�}�P�O4�Ki?����}4����� ch�6\�Z��fx(�*��o�i����?��"�q7�����r��_������&
��.7�����&�L�y��:I�r�n���4-��N(���F�Ɠ�d�����9.g�j'�|���W�I�QG�:mi��J��E޷j8MD�� __��n�QZ���T1���Dwj���SC��Å���+wK��3�ԟ4��Q4tUXvf�P ���R*&qve��<,
��3�>5CF]�_�g��t�����^��|�}�{Nv�����yg�N[p=8|AQ&�}�(�?�>��Û�M��]��%��p�8R����E����X��ۯ(���kx�i$�go�M�)t%:�|�K����O���gC�	qh:�
$��M�������7�AY�SlD3�b狵���ƏV�~��a�&+����2��uձ(���A��g]{m��f�Nr�]Iw�\gc�o�m���M[q5aM.�Z�	k!]yѩ�ł瞾��m{��S�0!��2r��=�JZ�)������~� ��yuq�#Z$�ȶ�aܺM*=ۢ[��q�Q�L�����Oza̝�]��H7J
��Q��4p��X5�!���R�tŹqwA����>��t��S�/fA:��B2��T�~���_tؔ�,���S�9ʂ�Gو�._:�ne:��l@�Q/��m|�|-F�bmk�F��-�0��1h�Q�c-� �
q��ְqH���Q����[�0o���l}�G�d�e��E�
Z����Mb�D�ʿ�:��b��m�\0���I�S����ߠ��s(�b�n�D�rF[�:�~�'�a�fb���[K���Գ��)��S76=z��i^K��u��X����_1 BO �W�"��։B�������0�d�3��2�!���n[$����"�I�Ww�'JS��7H�e�z!wj,ʦ�JKn�6����;S�[xǧ�z"��� ����ڷ�	����-��8��Hki$k���rw���V��7J
�o����_�d�*��+t�|M}�)�tFG<8�)� ��Dwkf%=�<�QŌA�/+f�+�d�m���
���ZM���l�9�ڀ� ĐԳ���qx[i � :���޸{5�ʅ�}ނ��O��)ͳbW���g���5�tG����>���R�鷓���7������=������u�.����	��Ũh@E�֎�G��F^�g�[,�p�h�4Oo�#��ߙ�=H��ib����倒
.u��g�pq��S��)lN/A<�w�����؃B;���jPȶ�^���w�Ggf�(��Q5y�7�O�Y�m_��M*�]NM�:�}s�Pb�P\�J%�)i����"��q5}r�3�/1�3��-�f��q>��zac~N��%��,%c�2EOH!K?��q	�67Q'G�0K����D����ʁ��Mh۟�,�H�xQ���OBt%��Q������gT��4-���������7�2����̗>�yξ>�cve�I��ny��^�ߐY��R���9Y��_Gִ(�?P�5��X�GR:*��_E���լ��8���9bG-�b�|䧇jk�q�#k��尤���g1NT"�8b;�s.��B~������tNx�r�,(�d�c���ƕ��%� ����Xl����?�qg�Z�=�𾊌��W�Lp��^�FH"�( �(EJ>{閖k����ﬕ�R��j�a4Ψ�\{��Ӣ�aA������m����~ev��m<w��zx�j�uN�*��c���Z�Gk�Z�H"`_�1(�&����T��9eF���H:K��?�Ӟ�k<QL����~P^� /!HBx|�l �?J�����Bp�X�O��S�;Aj��Ä�p��GZ,Ă:�i6ϫ��r~f����Y���ia�	��C��	O�,;�o��X�=n��|�q���&7wW`��d�>Hp%esA�����p�L�|;xWY�J�ś��O\܄|�9�6z���l�91s������f��%f)\ "���2���9���'7:ȳM[�as%�4e z3R�J�Xy���KCb ��	����D��B�L"����ǚ���&V�au|�7-��AX�j�M�KzmԳ����N#,���%��*��Vx�Z�'�D��_�����@�"�Ƶ@L�8��jD���=#ձQ]��yy�$V{�^���o���/;O���5TVqdk�l뿺O��Ԭ-R�Y� ���3_�%D�LP�Q+T�0���)�!$�Ƞ��`����Z��pd|v1@xy�O��b별�$��O�K�dC�uö��ۦZi��
��J��s�ԈK�ֻ$*ћT� ���5�3�T�E�S�CV����4�XT�5@��(�dڜx+�n���)1�kI!gJg��I����Ng �>!*(�_C㤭����а-�i,�1�DӞs�J%�Y�(�3)B�@{]\���|`�U���2�;��>[z���p@���T��"W�������.��O��X��+����s���F�	�q&���%�Yk%���ч*wX�u�ױ�Ry��4�G7���L�[��j��FA�?�#q�k8'�:�t��pЩ4�̈́�_XK���/��5���,����d��ӄk0��>F?���� m"[K4I�1����C�rQ;�41rp�F�e(����;�T6�X��꿢����zY�V��Ek��cޔ�����04���\]WX��6�k�.pc+�0��F��e���'�;�~���rK��HGh&��#��t'���}�ӄ���8QX�N�O�k���ie�~�����zۥpM�Y���"(H�,��:L���W=�*BT�m�IG��T�\����'�^��1M*e�hn�[��Lh���\��}��>�0X_s�'͘ӏ�����/}���?�Vs�
�?i�Z�\j�@k�E2����(N�3�İ�]�jB�- �1+����S^Īqew�vy���	�G�5�D�_	f�9Q���VJkAg���Ϳ�{��(��Ϝ��L<e��2_QQ{@���"��s���_a�N�1��&�S<z#�יtg��G�C��+�x7�,���9�8�V8.��7*\Z�İ'ڻ�/�rX-FT�os�s�朻4,$���S?/���[S�)D�_6 ���~�Ck��46����Aj�/�.(���k b��:��T��b��yD�d�]ĳ��0�'�e>{�;8��ѕ�S����$�:,9��rHIK�n/ ��Ս���rp����8xۯ"Z"���h_�Lu@C�BIR��Z�vN(�<�(O턲�PB�iߥ�`��[@� /��dԙ���˷G���W*�XM�q���7���/�+в���Cn�_�#E�1�֓��:@hDqv"x;��ZA���D`+�ނ)�a�%��+�#Ĥ�8�[y~k�� s)�]�Vm�-��4��f�a��Lgw{���l��st.��-���uE�<mzm�6��oU�,��D�ȷK4Gq��@��vg���UCU�fgx/994�]��VH5.sY;A���S�#Y�B��S���|akٵŮ\#�Gq�Q'�O׭� )�+��*bl��*]��%s���e�7=��h��鉪/�[ț����5��G��/=+�����@�frm�@���0����}̪�c������l�5"�kɱj^���Rw}S|����.��k���YW�(�FL�4�Ű,^����:�L�~��7�R?�O�'T8�"(e���9��`�ҕ�$f�=iGm����/�U3�Qi��� ;���Y�aB�QkY?�x��n�+����Oͩ�`�Тjp,EP��(ř<q�B��No���6��ּ�|aP$�kJ����f��NBLa �I��!���?�2v`I$�Y�Djǳv�']��Qګ./�!��&5z_���<��z����*�g�#_'��R5����aJ���Ch5��x<j������1Kn�ìq�k��(NRͣ�}���{���
��KU���z��G!ޥ��W�*ўLۏ�g$��7��W��L�ݦf+�;����F$7�-��PT�:�擂���8v�J��	��E�g�� u�sܥ������L��J)+�M���X#�y�=�.뤽�G͸��?�mÄ��f�@q�y�<_g��2a*���dv�U�нc�r*Li:�}ɧ���[0*��@�Ve��e�YP� �MѥN�ː.J�4H	p�Tj>Ƞ�����Y�K������Clͥ��1��n3���eGN��1��ʞ�C��RlP}~�3�+�Z�LAON�؎Vh��9���9K8� �Ѫ^ɍ��<�Y���ݾW~��k���?�,����F��Ac��gt:_�1������� ���Q�(WMKu�4�V*!�'���G�{ +N��8=��owB�p����p�%��#U�_4i�LnT������~zH&�8�T>�u�6;(�,��e���#C/�P�_�{��+��؝��c�(�o<���6�As���{�3����al,Ƶ���>G4�yR-�������^+L��N�<�nt�@�c쒄xŅ��2ò;��L��fj�-�$n����L���zG�c,a��)u���F�M�:x+�N�L��GS�.�]�6�g�v>L���p���0�����ŎN��{d����!!t�=X������E"Aߺ=�!cB�x�r
���w;|=u����wI%�����1F8-;!�G�;�I
�f\��y�Y
�?�x:=�:��