��/  !5ц��Fc=���F�jgg�.!l=l%!�uN��S^�6�)�Kgn���H8�`�BH��RXMTl#�4N�3����;p�)o���;�Xu^�V"΍I%���V���G��!��g� ����A=������4��Ó;
����6F{į��0Ѵu�;o���E�r�:�!����$�3�4���!��T0����諈H�-���J��9�TsEلY�"ð��x�(�/�&�!\�W ���$���[��Ა\7=�[��.T7�pā��:��4 ���O	�G���nQ����/�u�l0˂u�t���ZjO�4_1]���t؉��_Ё�[���e� �}+rz�-!SKw*XL�H������Pk/W:��1����w�R�{�].�M�T#�ެx2�@�f�b@]�qA.+`'Y�+R�)} vի���2_��e
�r���e�2�R���Ǩ W�l�v~�Ī&��k�L�aC���'�x� J)�8�՚�]��|��N9qwV�\)�Eށ yTǚ�l];��u��hUx|���_�/T�V�q����Ea��d�WyM	i6�}��,A�/�+���*�y5�=�����q/k��|Ka���e�TU>�������D���Ҥ2$75I�����������z�PϿ$�mX�<��B�}7�Bފ�Z��2���j^��������;eN�SC%���r�w��=r���xnpٔ�A�n#��6xĩ"��r\bR�1~ѷ�3U�孶ϸgR�Z�E6�/ێإ��ņ.�h�i^� ����b�QԒ��"%N�,)���m�d�	�����i^Ϳ9K�GfV!�&%��`�V��q�[ù��W^��-��<�k���[+���3z�/U8����P=�V��N�$Y�[��91��ϡ|��w��9R��x�_�[&24�v;(�zi�~n��h q�&4��,� ޫw�u���#��rb��^�m����v��7s��_4u�+4�^��gl�ٕ�
>���3�.��D��ou<�9�W�3�󥴈�-;r�{'��D�v�\�==/�U�nI+��+�Ie����׸��Y:>��|cp>Ce�o}O&e�����W-�lrυ悤�3T�
X����s��Cvr��E-�?+���Q�SgrZ�mz�4�<�Ǩ�ӿ<��Łt���V3����p͝%3�	��ӵm����-�#KP�j��ş7�I��y�gd�ka
�0U��:�!ljd��_ӎI�VpQD
I9]�D�,�"��Ao���� J�Ɲ��CkW���O@�
e�-���SfM�
<1��i�_�KZ�K.�*��s����\x4�� ����3p�/���c�u�.5wt��ȷ��1�|-}�j�����19�ԁ���+���f�=�R�ܜ�zTM���-�}-O��W�zH��K(Ƨ%�S;�0�B��H�$�L?ÚG2�����rE��&�N<lc� 0���a�����{��j�ɼ�_�"��L��i���%|#�Hg�����џ1zkK�]���t�bYMA��8����/<ϑD��U��G�s�,G;��p�\e�$��?o?�LV���Q���0��Ԍ��T����׷���@�,-�M�'8��K@�yx��/�5:���~ih�.sJN�K�O�B{?��Ts���ˮ�_�Bމ��$Y⇩���� ��f˄� �����_4'�8�8��_�Җ����#"���~W��|�ęTΰTR4݅��>Jŗ��*2+�3ҨH�X�K-U�3�,2�6	���n��� "2(�'>�eN#{O���d�l�sA�,.Aiw;� dvS5l(������ޕ��g{~�h�ǯN��i� �k�c�*��ۯp�+֕?�P��:���P��=U��5|�:���z>:.��X���<��L��8����Gv�@9!�8��R����_c��_�)&�e���cHp��4ddE��3��2�ƣH��7��U/_w?� �H���vr9+�ţ�{��7����T$<�N�P��|�L=q�4��GOFPK��,Y� �*N�m�p���:R��E].*T�5!8 a�����%P�*�_��M�ᄊ!��gZ�rǡ��Q�,���+6l������R�^�ӿ	x�Ӏ�=��6|�ɏ%)9���4[�{�d��C���S�c�vQƜE@��5�z���m�Ӧ�8]tWr_(���z�/*|�A ��By`2M�-	������>2��R�Zu>���*!�+�P-�8T(��3n��$�T!>�\bV�����z� ��09����J0t`}#mpӦ�5������}��]��ϼ�i)ԍ	�i�SY.���[I�"�F���*�j��E���h�C��+Y���T+�7V�e���O��]�qj�V��}��I�,AU6*[�&�OB�pz�䧱��*�N�w͹3t�_�sV��I�6xA��%`��R����^8x6���v�S�e���^ ��)�ɣ���%:��pF܉�Ae��u���� 6��)M�*_xǘ�nS~w���Z,�]����LG��8	��+F�~��l�Q�=s0NM�^[��jK�ptX6(8�V�B�Wh<��A2���Q�sKml�`B���kbu���$XBl�thU�|Uq'A���Օϫ��>�F��N�6##�?Q3\�v�y}�g��2�kN,J��>��%��*���%���Q����[E����ٶh��8������XNPg?V�S�nS��ʯF_͐�������+�S��I~�MK;�)�����k@�tU���c�yȓc�ƺ��8���;��ވ'�,��H�z?ޢ+J�eҡ�rJ͆��@�q)����|C3)�ލ*�7#!qz;�����"�I�8W��g����8x�+?����9�Ư�� �il�����I�&g�u�i`2 �@c��(?f���d�i _2$���o�I��>��6n&{��ի�� ��5>�In���lr�]�4m�WQ�3�qֹ6@M���9r^�U�og�y?0ُ��6�5�l�Ѣ:��쿥	e���a��퍅N�6����j�8l啗���xչ��Y�s졆�~��}�  %�	w! ��LA{ӝ���m�U�}�sO����e�5R��,9?i-A���W(�9��qS��dEA�ֹ�L;�G=�&j�fBRL*U�uY�Y�ĵ��gK�8����u�e� P�N����U�� Ҭ;�TW���D�aXөc$WW�ł��^݊�BSF��q9s���K� �[ڍ�iu���=K'�������F3�`����j��g�n��`�^�f�����S�����I�!��)B��������I��#n�y��/��˅��Pܪ<�=U�����SL|��|���f��U�{�Jo0/�6�X��~�5�BC�[��a/�M�C1�y���.�ǩ0ȥ0��$�a�[L��QnP�yq�>�6ι�L-�f��4���*Y%Mz���4�F7������2�!݅����B�;(�������X�}�D;2������_��8�f�N�6u:	�����-#���1K��C�z^SE���f�{S�X��m7'f�bU4MW�9�P��̡;����'��ή$����߀����Ga�a�5;���?|L:l��h�!��;�s�m�>�)��䊏j��bR������529�*c@�2��K��@!�C��F8�T|X3
�f�HZ �/A���H�+'�8��ӶKC%��4�o(j�Tc^)Q_h�Q��ň]^��Ug�gw5�Or�qX�Y�buV6�ń�5;�|8StM̙���N,��Eʸ��#0�؇?��X����4�N��s�-`i2����C�v����<󊔡���4����Kk1��W_ȶN�l����2ި�o�oe�?U��z%iO�;l�,�Ҏ��Ε�U5.R/�
�U���7B�:��<ٵT�ʎ��]����P�\�G:�e�W��_�&b�W{Պ벪|��$/݅��V��P�k^�)��LRG��ȊY�a��.��ɍ@�/��C�4����l޷���C	ِ��6�
nU�As0 ����4=����qڼE��x��+�r�n�ۇ�D22�hq���P9�]�e���Ľ��ϥ���Aߓp,�9��*��l͌|K�hI�OE=l���OV���bK�,�?�{?&b���yt��ߝ��{������ Yg���1g	���,_�	�s0��,Vw�F��j�%� [% ڽ�#�N�cչA�'�r�E�g�Ş/VJԴ�֯���_*݁5�1f�C���wr
���י�#�.��$�2g��Z�`�v`������-Cp��a�o�-�T'�ow���Y�LA2�w�ظ�?|v4��`bC��"D�ȷV��L3Q�s��h"���sO�����%�;���˛&���uV~;�,���E��pc)��]8�(�4��~�m���\.�����4��Hl�����Q�q�˂��>��/�[sn�eҦf!@�~D���k�g[1��3�5�R�`̸�o�A
��L��A� �1y���e|�[۶����Z�? 7(�섄��hN��y�*��j�� ����SR|SX�e���?�m��ԒȚ��:`J�a5�K��6p�6��SMƞ�.��Y�$Ե�_,E7��#J`;�t$�TH�X΋�/gO(����ø�ф�""�;c�Q��ȑ�։�S����W�p4z�3��븛�G���awI��̫���o�t���`�"�Հ���H?#p��:����H@��\�+p�k%rJ��|Y�i�U���c��䓞��M��������Ց<g�E����n/5r�j�]3�.-�U{��oz L�,yP�LD�gSY��0-jYk��Ǭ��n	��W�6��9�?ǈ�w���I���g1��k1;h&f���Z�*�!H�r�B����r�s�=e�g1|{�u��7���`者HV��K�z�Bח�By}����3�����'�Aᗝ*��"0���-��^,�O�`��]qޜ���Y�3�4���=:e �f�s�}�}��x��&K���obD�&��H�lH��*Z��ZF9��;S����Ş�L�£��f�iՉ���$�i�Iڴ<�l���x-p�W#ξ�o�3�S�ń�2bu���;�}s�� |I:�O���?�� �I傟���#�Zh#��$ݺrT1[y�(ݐ�?eǉ<������Ko�Xt�
��(���X�Y��^�jݱ���}��k$\~��_�A{�却���o\j\�X��w��gn㤉�?�!��(�J-ے1�F�a,�p�۪�#w�{U��f�j�z��iH�nЀ���=�����V�L��t�雰�Ѐ���8N���0��5�1��"o"9d���er�xb��}�7"���2.H�1{%�;I��j�$�q���������8�c�o��=� �qHi���g�}c�LA�Y��ą���QOv��tR}�9����V0�عI��=>Q%�=]�h<Q[zZ>�^z�6�jCR2.�<r�׆��eJ���qg�iݴrK]���Y���ܳ���1͟������$����A��U���%����	���KeR�2Is�g�Y^��#�-�\���ps4,�lCy��Ø�����t���zZAx`�r�Ì��z��Z��)ʶ*�`�{<Qq�3�����d~E��)MC���Xk(�U��tK��jIދq�#��>�g,�P\V�8nÛsC�*%.��ໞ<Q�c=���?zނ��?<`"�c����;5��~�����ƼI��Zr�>�C��R��bKE1��9�����Ծ05s��f��3��H�(P�K'�oO�BQ�sq$4-�wq
A�{w2W����Ňjg�*��Z�#�[����E5��ړ���y��ݮT�OZo�v��)WQA�Ok=�����o VYcaV��ܟR|�Q����'7�o��O�_����w&��ȭ�=b�h���V��"lZ?G��t����"��&!�X����B�@�U��j,�?�YI3Ch~OY����y��#��������u��o��(�M<h+n"F�Rhr}z�j9��%a����¢����>ʿK���q��;U���{߮���=����"+��KQ��`/���w��\y'��$q�-�A+E��Jb�ٟ���TDal�}�a�`'�A_Q1�*o���
Gw4��������B%�dW9iZ"֦k֖�i�D.�]�Yt�{��&�"Dd.,]�L�8m�&�
苦*n��I#Yj�}��H���,�C��.{��'�՘�w��9���-�R��D��DjyI�-��=L�fA��`�9H��-�Cx�=� �U��9�K@T"^B��=�r\y1��ʶҨ<�d��(�U�{{��9�r�6�L�}#�+��m
������F ��zH�@�;�@_X���(;��_'�;,g�k�O��% ��&NP�::���5���0e�"���e���k�+
�
�є|�.�;(��:��b��c���y	SDl�k�.z��J��[�� ��+E�;���\ڐ\��'u�@�t���O�ugN��c�\���	?G�W5@u�|����fߗ�2$�ŧH}jF̓�d��F�%�/��ɒ�V��ᒡo 
�=l�M_&�LFb!��D����ѐ�f=�P<�$��_w�pj�J�q�C��>:��'s�m\�k���\ߔ�hVo?�#�!�D�L~e*R�ϡi�W��ԑ�̞�[1�	,&��"���Rǅ�ߢC0�ZѵXc7E��4��KS�Z��R5�a�ڥiхU�����[D�>�!G֞�O�O^��4�g���y������[`�z�Y*�U����O%|+����'.;LK�N��U�sa��iF��޾$vn9�X�+�'&�?�Й����=i�,�4���>O�ba@�}c1S�G�*R]�O�����>�sL�t��XS���u�C|���!�BOè�<\0�ǁx#o=�L�gP��-	[FO��@w��J��s�q����GX��.���$ ��T5�Xdu��s׿���tE�w}ֹ��AM�3�����#���h�G�⁽3vutG����:'<d�c�!��3q��� � $��R�c�Q����N����-?fyq��$��Ho;¢Tb��>�y:�6ҙ�w[6���E����U�!�3+�x�h�"�tC�H=�ڦ)Z�3��!S���������H{\?�I���p�'N�6R��*MY���V0�Ш��k^d9͊�?f�X��*���q�4 ����4�����:��`��w�>U�-ؘh���P���e�/�d �fm��uu��V�Ň6\��*N�����켬��U3}x�c:c�\�S��U�"�Z��͞g�/�w���'�A�9t˹��Z��*�8���0h������>U��Xu>U�d���Q�C��4S��&`N��Oi����n��YC��b�������u� �$�y�}UUJ�/["8 ���k/|0v�A���+�lF����C@u^	K��0f%�5OB�ho;>���q�Y��������]���f�J^l����A9���g{���������9���ڣQt���=�HD����?��k�/V��.��#���[l�l~x䔍~Z*���7I�<`���R��E�,�#O���e�q�V�[Üh�4�%��wX��{%]��?������JC�٘��@R<_oG\$�ʉ]m��y 6r�J���!��&�0��N'�{�>G�|��e��`	8�v���0�o�`7J��� �_g]��I�J9*h2J����S����ID�T�)�G�vB�e���{Q�F�)�\�sk��M�4�^x��y��Ⱦc5K�L2N"� ���y=H5M�8�i ��*|����l�\A���S�)*�E!��'-v�j?~�ƥC���g�ҷ�@���ىU��6̈́	��L]�v�Qx���]��B'��PQiv^Q�H�p<���4g/��X:������;=���T�δD�}�&m��^��o�̑Y�?;�q������+�ћ^�ml��Lc�P��太�-8�`}[���T.�@�Z����8O3X���#Z���nH���.�Y	l����i��D�1�&��
[V)��ذ�jXN�eѷ��ut��ښ]�	@�����h�����z]�\�@�����@���q�"&4�&s���0`��9	��O>�����5�����ݓO���߿f��D���\@�µ��˻6"�7�X׸h�ʔ�8T=5�<�jn���-�ۍ9��N4б�"f�wۄ9�%;V�p�`�@�,�����3ކ|���c�I��߆rZ�s����R)�ܩ�3S�R	�O!�5�I.���ǋ���@���U��ڲ�NtԆ)�*%�x���3OuTH3��nj��/+妣���٫7����B�s !���/ڜj+��W��s	B~�)����f�NO��>#A�-A
ȫ:0QW�:{ 3��É���<[	�<��Lt�	#7��V���'^��BZƳb!����í^���ܱB�87q�F��US�V���	�&/"�%�KV�A�e&�c,K;�fQ(?��l@M����"X.U�XO}YN�p������ ��`Ci�� v�D����9�g����D���gC�N~g��>K�#b�<���XS(9�b,q_94[#�vN�w���6����T��)S�c�7��r�d��k�#���of�������^�WD�埔���7�!d���W�.Z�k}*	��%��9���n�9B�ޱ_���0�&�^rt�M^$�\uC%{�����-1E�;{cm��x�Q��?��C�����m�h`,n����ء��BaE-8-0���=r:l�|HhWf��~���w(��>=��Xm0I1�ަ�6&�N�y�pm"N@�\|�HMw++�2@����o�i�K�,�/z��s�\a�3�|� ����t��^�����w��ר���z�ϋ"	O �q��M�B	�]��ܜ/IN\=1�G�\���	������ r-].%�|���cUK}M�R�U�XU�
��B�$��*�!f���^P�@ew�K'e7�%L؀L���R���jJB�ѝ���o�6���Ja5�1k}8��)�q�>O�w�'���jnt�`�R�J��:��{z 9ur�X��!�j����4VwR	ft^���[���T}�Oy-N�&��?��m��F-S`A3�_�T>QU�/�	'L�:cM�v0�u���}˩pp����u�?w�����HT��{��>A�Z~���Q^�`.lK� �#$I
����x��`̏q�M|Շu�'���%�V��\0���o�#B�`����=ڑ�t��8v+��V�������2Q�S��W��Ձ���3��#>���rvV��.�I~��ӊŘf'3�H���~�Ŀڊ�� m�����aÃ6>�A)'᧬��ψf��(M� �M��+�m����*w�Q6u(O"��˵������@N��-[��ޞ���"����H���U�?L�؂mu����{���x��^���F�\4��{�&۹��78��甡�����G�YVǰ�ªMj�N����օ	������@��ڢ��5��ފL�L�*��!乆ORӌ�������n��`.0��Y��锄�K��pj{"��F���t:��8-��-m��r/�'И)CH��w��:�i5�c��r��"�Es:�a�׊�!�^�,�h�/]�,��� �9§��릋k^"*6S*������=ˋ	���@-d�Iw.OGJ!���r�>�.6�S���%!�������^�w^���t"Q*ps%b�h{�9�Q�{*�zDzB��I�)m��T���:s�7
����N������>��>�H��O�3�i�u7�� ���i ��n�E�sA9p��Zn[Y���%Y=���h�T�|A���2��=��1�^��,�3�8QWts7<*[�
��c:�@�'��'f������RR���u��v������x�( �U]�VK�o���S�6ٮ<HNܝ:�t(�����'�	J�+�nθϚ�&�=�@)��;�`�V�v��3�Ip=R� O���η	����~���.މ�N����d�����)�ce����V>��1��{��q7����^�<��Q�*�H�Veȸ�ј�bd3�l%�}Dgx+Z���K(��1�I����HQEo�����JX�aOjg��I�fJ:��]�������x�����m��.����g}��+Rhi[p�xLᛝy�I�p!)�<�c�P��}|�J���m����ڱ���F���>���LfC�0e,�V���W>���]�����&a9Β�m�$\/4��G����֌=���m�C&����d�hP�ie��]Y)��s+J�!��d/�h�ORl�ʢ�=�c��ۂc�
��c�o�^R�^�Fk�j��\�C;T��J�š�
L&!�-��6�����ݾ8\�l���2�Z}�%��2Z�{���y]�"_��y�(�AF�Z�Qn3xe�j����ώ�4(�r�x�k��3�]}�y�kw$?G��������ő��f ��ȡ���t�8u&M���'��������m�|,T�g�ld���}��4�,�'��m�K�<E��RUX7���(^�P��z�#�Kl������%fm��-\gҿP��Iާ�����`����߶��G�_�`Y]��V�W�_�[_(�5���#�F<��9��8zl��6�i^�L��b|�:�k �{��J
�(N^�>�H}2ܪc�h�b�?�X���60>;g�	o���.��P=z�^j�H��L��'U�HS��(��e�"�/u��� �����eCZ ʌGX�K�2vv5m&r�k�]�%>�^y�T��|�d�+��s	)d��˱.c����wZ�V't��`�lA�i_���J�9]��
�̆�?��JhF�*Զ=ț~����ƩN��&U�/��X���w���x Z�����+-��jB�v<�H�v���&&���I�_I�2���꿑�I�8������/!��kW4��ac\8x��l��(q:��%'Re�����X^&!D�-Q��V�a�"�m�a<U�'	�ް��Q/Ts:��N���9ϰG\�*�$U>%a5?�u|�e���lۛ�E8�Cƌ0�Pj��5��[9�y4���5B��x�&�~�/oXb�◓ຊf����	���3�5��Y���
�Kh�N�Ԣ��  幼��]~!}Yg���6i&6�
�y�i�GI"���	sn�)N�Y/���}ɢ$�?G�Ew8��a��ymj3����0��[x�[<�WW�_8��CmC����2�s��0�U4�s?Nn[@q[��V&Q2���,+1��7���i�,1��hM붅����ԍ|�kyS�B�K�^���g��N�nw�)�%UZR2�j��^罻M(Y�wku�,�o��>&��y�CSo��!+����4cD�瘜�e�#���?b'23q���ݎ�(��ض�;�K*y�R>u��f��Hԥ;�4��:�M��x0y�����"sF ���U�D�B[p��c��x�SA���V�e�%M���˲����ةd���&m2�ig±�]^�z��Iv(Q��D�̃���.,y�/�ia�F�eJ	�#+i��������RJ�}x|>G���P�ưw�W1��r\_�Q���!��'H�$L��}7��)�l=�v�����_vѠ]ֆ>��^8%���d-�k}���t������Ҵ�N�u0��j��q��7��"�V�F?6�\��C��%0���梀���k,!~��'S����u�Z2Z*���f�Y$���47Q�!�:u��h���}�_�J?Kp���sL������ �Y ��)J�,���%w���Py<��z���;O������`�����N�
�|��֗�1�[�;n�t������7��]���hM�Z����EH�O��`��z�B����l���.N���5��Җӥ2��1c�)��"�^8{�W������-�8?~�d}���6gl��(�]�^�T��ǎ�g�V�rj��2!�$Ƕ���Ru�M'7���#B#b$�)ن T��}�?��БL)����r���V�z�'	m�*�k=s�Ko(+�[��i����1�6�b�����O�ՙ�vLEy���|�y��aRl�c��q^��+:C`�K���.���l���M��8T�gl�����˟N�e���vL,���
ɨo�8�w��afF��m?�,�E�aQ�cL��1:"{m��?�[[�RU���c�^R�~��b(M+3n��ਟ�`�<Ǿ�S�E'A��;&7��1����=>?)��G(����L�뜣Y2�9::�t��$&�C�/�cr�oD<�&Or&m�i��
v7xtص���ֱ@��k�����L�E=�#6�˞��}[s-|\m��5��t� � ��	gEzF	4�3�m����4:�`���9}�P���&i�K�>�)=���h���.�*�}�MdR~���V�W�[;��p#8�A	xE���z�}t<��)�Kd}��2��T�kо��=��nڊ�QoA;eR<�]�E�����2��X񍗑?xU��"{S�+��݉ԅ��t����H�s���2�_�L��MLl/|͵Z�UE��>P�=�7�x�<�LTt$��r�z7��$���6�o����"n]�dcg�E���Xϻt!U �j*%3:S���c�	ȭ3k�jE�#]���;Y|�XXI�|<�`�f����z�24��U�>�P��er򎷅������n1:��/T��j���Hŵk��
��k��AY�n�i`7Q��ܒ�
�]�ɞ�U�(LU�HN{�!��֗�;��OC�M�?��c.�R�e�t��}��X�3��Wք��F���ÿG�˴����	�n�:��0X��j��*t(!���J��`�M�ij[g�����������Z��L�-Ѱ��O�4��:+��a�r�5nÛ~\aS!{�; �цz�^��<-�)�L�}�x�n���r��eD9%�W�8���N�^9��X�������5<��5F��7��nr#�����D gDa8o'�z.��љE��ԧi��Z<��i�z/DwF�"e���9#���Ϭz(G.I��`���^�s6�{ⳣC��RG�񃚉�����ۯXsg�S�(�[�����D�fM�w.�r�)�Ge�w��"}�\�$�n�)R�5I��|��-��M����}X(=h[}��g~6�E�W��s��[:��/��Gb�i�X������)\\iqQ�V%��JV��H�݁�n).h%L�;�F�{��3�睑���P�-��͆�;��eܰ6�=i4������e�/� ��$��׷v���gw�<��ا�NБ�9k��?y��X�K�`�l$�lV��N�:'����~���N�[`)|~' �\��+u�GͲ<}������!�:N	�?��WX�q;���,Ϳ�P׌�x��Z�;c�*v6/;�v̮��J����S/�:�X�=Ɩ����S��� &���R�Ճ��"�˂m`g|�@"ɦ[/b	����r���Vk�-��f�MT�
�/_`�Z"c����2!��Gl � O)�O>���L�p�;P�����9��.��3�a������q��&��f���&V�[�
�c�����D�EU_\�y�FP�w�%R
JH6p�)��J�f}�e�T�P���K�oI�������`x���;<"��	�&@��I }u ��ϞT\]��,��8�(��o�~���;2��Ӵ�)Acee|i^_`���R�&]�T ki���a*�k	D�2a�4#t�Xܵ�j��X�3��ԛV$ָǅ`]��؄
NL��P��F���GTt�t!T`�d @��n\P"ʒ�uCq�].Z
7c�]�77��eGu�z�t�?r�����3�3� ���RY�R `�&Lz�����D+m��7�Ko7 �<ج�罏0�A�YĄq�+]?����˻A��� ��ݬݕ��Sh�A~`U��X���
�X<2B��џ�1�ݹ���0��":�w@�[;�06Hg}Ur�I�*ao��!�p�j�W����D$�H&4B��i{�|��#$�e�|&t��L�G����x��ˮ�����6�Clj��+&��2�64=���H�au�X�!�[<*i���-�zL�v�0n�7��>|��S�E@�u\~�'��!F�4?���C|�P�� y~,�eZW�U]y��w�9�e���v;����'���De�ҡn��z�Ad�ܐ��,�H�esMi�/�G�� ہN3��+&�g	!������o�q@B��*P���낌q�n�+��N��:/b��u�f�N�,��'=��N�/�Q����{�p3����z�%f�<M����G��]�I`u��ˉn�XN�i2�|7��=��w��w3�a��a��c�=�F��D&}[JMq\�й���qo+Gm���r j�X��S�	��	�sâ%��&m��f����nxR*=��)�f�_&����;Ѻ���,V�u2�M�_��H,�5�(]Vќ�C�n�vZ�Ï4�t|V(�`Bױ_�n's��ۡJR��� �|�-r�c/3{-��C�-n�A���y�.;VY��eQLǤ�yT	P� }��1�X1�}�g���ZӔ�r�R6�z3�LZ��j`=��fö��.��+��$�ec��yvI���X�\��o��6��.ϛ������/Ho:�O돢��m��B�8�f2m
	�-7+��I��pb��4�b�2��Y{�ʪ	����,9@'��T�h��'�\�w�Ńd��cK �� �03t$�A����9V{D�����0'-��y ��,�R�恁��xd2���o�}Q�>`����6����C��y+zף#�Nѱ�탢t���n��<G��������j����^��4���f������Sgh�WS�����f�9xo0P��칓�1gi ���t����Hc�YY
�9
 �J��ч�
	��.j�cti+eq91�a)��=���dBw-	���rL"D�	��5}�䖪�ؓ�h
�ȸ��sb�wp�s���ժd I+X�ӎ�����W"y2���7��KA��ӥ�����P�W�)�:v�8���t��D�L�L�OH�AѤ��*�pMμ�O�k��J&��'���?�Msj�t�A�szKd	D/�l;� "bQBN�TdM\4e�S}�^�1O�yC���UKV���gg����=k����O!���O7�l�:�}�����z��^A!��Ru�+���!�(�j+�x5Z�B�Nn�� &$AǿG�ـa8�I� �8��@Da�up���B!�3o۰�',2 O-�Vv��DE�[�M�A�à�2��1�R݆ҡ�j�0��O�*���:-��.L�$�>e�&,��S�y>��]"E�뮗���3b��X	�M`X�X���hz���P�\�>i�1T�*/������1?��J��gs3_GT��Ǯ�Գ�=y�������J�W^�AuRS�7��*l���(�v��{�XӲ����%�4]|:�M5�S���D��G�o+�5�Id�5���1+���We���CVo����[i�0�'�zT�l.��f7	*g�i�2��!zF �ȹ��nn����or����q��(OS1㠼��'0�[�2
+S����y`�w��3��_ �#/sjO�lr��'S�V�{��+��uyd77� ���Zce��_)zw�
`����!����?t7f�����#8��{�5��z�)t�㩒�N��d��F�Cf��1�i*Y�w�s��;*�2 �mx�:19if
^?DI?@��O�\}]���H<�m�ߣ�$��f>���.r��կN�~TI�nBK����D�����~�x:�O��`�0=��~�}ؼ�(J@�^�I��kV��ֻR���� 8F�Շ�J#��£.�*��������֗�0��G�$��jc'l�76k��;��=��Z7:6渪kN!3+��@u�{�̜�B�o���-F�[>vס��R�ܘ��m�E�س��������Q��
U�;�`��ҳ�F|zU����VL�z�?'s燡�/Z=B���l��e��gIdo�F)�~����,|�zw��a`��vl"v7p�����8Fs�$,�'��o����@�:��4���k���;��#��9i��r�!*����x+I^��,KPf�u}J�(>����3���/	kN�r���Jg��j���������i�ޏ�lw1���yҁ��E��k��AO8�Z��|���!}���F�p��(���H[�%x�2�'�W�mn�P���;8��XLق��c�����@ph�ׁf���9��M;�H]��Y�~T>t]rPA�J��A��;���}Q�;H��fP����W��<_q=gs���5�D&�R�V���AN�9A7���X ��"�����Z��޶B؊8��{	P5<��������=V@%x48�JA�X.Jay	_ k������{ǬV���!�)�����](�F��R�����_��XT�NWv�G���XS�+C��c�kP���J(�	�r�"��n^��#���cmP���	�e�	��\���i���]�X<MqJ��&a�����B����M����e�mS�1�p��L��[*,����,杛-��è�ٲ�Tfy6��{ć�z�v/��c�]���Hv�_N��v
[��?��z2����UA7��>҆N��������ґ�ڍj�w8�ȚPaa� >�He�ߌ+=����p}�ˍTi�>�lV���4�����ot��*04r�r
�z'?e>����(�Oz�r8�3�)�3���8A���PH}�T=?`k���IpHwpĳ2��6�42+�!A�B�����.7>2����Y��OcD	�݅�]q{Z|e��ŝS����LԂi��11�N�%��$�O@�>����,>�+�aI	T�(�`�S�4��E�ަ����$a�:t��)F�s�Y�U 5x��q�:�84����a��S k������W�AC�!j������o>AR�й�M^�{�I�i����=�5v��,Ӿ��=�w؏��_��k�T��烊%V�?+�Fi�&����K=Q+�Y�|�O�{M�=a� ��?� ;��ຕ8��� t �=����D)%�7�p���iH��1�x�����oI�>j���V4 :�"�c\�n�9���	�i�54�~�2��3J����(J��k`/Q�xP�-��1>J����/�7��HZ���l���"��n���;��	�x�6�h���v��p� ��\w݀����~u1��xt�~W��QB�x
胆Q����N[�K�YQ�����a��fKe��t%�Y!ۓ�k�>*1�4�]\V�.�8:[Vj���p�?jgk~[�뿬�Q�ϳ�aY���	�UJ��灈�[�&[��
Æ�W@%���H�Л�??���1���� ��sWׂ��,M��I���K$~c�)���y�G5�΅��f��fF
niA`�����q��.Iَ�i�3��ơs�'lH5���}�΀5��,^����mHp����v��Z3<����s6��T������#tg�%ǮJ����'�����h�2�_�F�`�1r�Q]�%�D�Nr*E�D+�D`�)��14��u�c�B�ʤ��E��?PhX�o0){%��G�����z�0�^bFaoE��y
��rt�s����i|^3݌>�'�;(�D^ǫ$`gG��'�j�
i���T;Ί�p�>NΑ���A�FD&���y�_��v��p�w�?� �~���DB�:-' ?o0�]�̄��n�~O����.�b!t����K,3��]�>�k�#}����w�w0�OhT�c�P"8Dm��C���'�(֮Rp��g�'�UDa�������+!���H��0���i�ep��\��瑕�
�]�������PU@4P`ku���Q��pJJ�%��K�!�k��[N̑�2 �!]�k���ӝ�Ey�=�t�h���������Y�sε�󄭭���9�p�-�x��5����,�6b�a �%�(����T�+t)���xa3��B_��J	_�������|��I ��% �9TI���V�c�Z;�_e�-�E�A����BQ�/jc$����~?hE2����T��%�LTfq�Y��$Ϣ��1򥍽?&�f
���a�-�ҡ��f���js
 {�;cqTKv%�lh�JU3����H�`�;�S��ב%GFΰ�K�ûj�۬��@?��nK8���V��=b>UdWM�UH|+��8�[��3҄��$Y�Y�[ޔK���n�X��J�����Q��?�t)^��ņ۔������ڏ�r^���<�N;*�[��GK/Z*����!p�[eۦ�}:�*?����|2��2/���[�涤��Nr���T
�~Y���J����q'��G$Q�+������k�~c��qH�ؚYȊ嚲ģ����~$NH@Au"�Ϲ+�'��63�6����,��?ݍе$b;
sm�0��ҭ��/�x���q"�'N)s�֟�]��{���E߭m%}PO��7;q���~ ׃~�S_<�O�ׁh[1xqxi@�_庲��p���l �xօJ��!�\�a�)9�����B��RE&�@�~ܞ���cA-���?�`�/�Y���G1��&���xm�Yk"��j�+���xv'[l?R���H��hݚ��V����j� ��{���e�����ܿV�@Ǌ���t�A��@�	V��E@���4.{&�K�o_�d�4L����Yv�ո;�*���@�x����E���wS;q��c��� �O�Ѳ�l|�JmE>�! �^a�����G���ჭI0)hמ>)B+�N���@�Nn"+��4��vQ��-*o��4��V�]]�h N%,��XtE�i�j���v�{��:��ق��4G�#��C50�;M�����E �H����PY}���Ŵ�0z4dB'��F"sF�B���ǩ*�z����Ͽ�b���"���Qxζ8q�
5�E�ڀ6�ZL'b&���F��8�QN��TD����o����V�	P�e�qO�z[(�NP�q����u�:s��1��%�T�1N>r��s+��Q4���NQ�/��p�F�6�z3���z7Z�3��?
x��P��qou	���!���E����̉#4,�F���5���Ǵ��Y7�����Up{�+������o�S8nв�[�G,n�<\�� �“�\���L���p�y�<^^)�~�%n�r�0����)I[���6���fDW�T%�g0�*�>rB󤨮�O�'��ϐ*�R��@���bpjO��B��y7�#�������׫Z���2�gCΚޛ+����F�B�G���;�J�����8����+%�Z����Z�� ?�5\����r�}|G���݇�~.��I^b�̢c�%��__�^�Pm�� W8H��&c�g:�e�0̑�|��\�1ڄ\'Fm�U�#~��C�yo��΅����cƑLG0�q��"o.E��@i��i��=
4��]�҃�Xdp�*��z<�$۬�R�!��ޮ�Vɾ��V�[� ���p�̟��Ё�O�������y)�rʄ�9��}&���/�퍹r�l@���q�z��&�5�S	!��qb��L��Ry�cJ��l���:��(t�lδ��+1S����ƽ�n�����g�d4�k�F�\,�"w���Of��^�q#�ޒ>�)������Z�d��L� ���_���ʨ�<S�F�PB��E�h�u�ٿ�|�5�p):�*sc�:�03���C�T�$��<Ƒ��ʊ,1O|bc/��ȯ�F[�`��9%��&Y�'��b��nN�8��!�%ΝP�\X���t��5�|݆����_��! ���NPw��c2�ǩq�s2A�o;�2�*<{ϓ6Ӄu�mL�vQ���1�j��/k"�(@K���#%�un}�&~���zQ}oC,�T��8[�^L�
�Q�C�~I���w���M �;�z��̰��L=>�VI#`��)1�KR�2Q�$��,���9O��<�T3 ���̹�TV�LY�l�$�La�Mz6j��lQKҟ�L�����]ں�Jq�@��l�{J�x���VI���ڀH �65 p��/7�fU�a�A����ĺ��@8l&��J��
��z�.9{�S_�+�'���j�?��Qsr?������.03�����fk�Dd��X��36��P��5���yr�m�u�̙�����r�Sr�=Å��pP�P�VU��?��R[�E�(J*�����Z���kj�6S�qP,<q&�g�x(o �0_m\tc�,����"�[�c�+?4HY0F����T]��Gd���>=�ZFSV�;���1�Ǡr29���i�=�SG�o�:����X!w_�[��=^h�{��Y^���m �������r�qM򯳅*n���յ�Ue��Z��Ș8G�\xQ����v�v�S�9s���b�M�K{�����d^Ɋj/��H��9?�=d2���<����t����I�ۋ������lN�#冸�*�<�Ԩ�$�L �)�;A��M��I�R~uo��򦀠����g�폡�?S��=��P��.�ゆ�Gy��#U�>y>�G�� ��^�X��
�ϐ"��
�A"8�0�E�0��2i���	$�E
��]�qM�kv�����;�Uzc�H�je,��y '6N}*<WӔ���4[���@H���k���uv�����:ÜS$A��GO��;��K�9�Vʔ�N$�k64��(����A��4��SY�~k���0'ύI�r�T��S*�-	�e�9��WV�2q�E�n�e��tqJ���2�퉵��C��_c:��O]{KIq�0���P���/}�0�K����0��l!>��Z����ߛ	�(�n�����pi
�G ��C/�	" O;���=�~-*���{vEK#Qq�G��=@��8�UNM@��mۭ���@�~$\ꝱ��f��� ��~��J��ok��L]~?�x<���s6���hl}B�����\��m~a��Y����3#�]�E��\���~��&���/���Y��"�n$�^:�ɋt:X�+9D�_����@�\E����K�w_uzȂ���c���V���Y�;7*d�y؀��v���5�3�}~���+��j�VN}��FR1}BC�=7a9���7��z;G ͺ\�kt�}�\ܞB�@����BP&�O���o�Ϛ�K���[5U��}oJJk�U��؂i~���.�+z��vс���Xvv-3*�T���Ƽ������{ķ6�V�fVO&���#������[�=�������V6�k�٫�vlkr}�S�	���$�m�� >}�ٱ~g�T'%���n���	�{�޴���u�ڻ7SjrP����"�9���3�0.>RS,݆AŎQ��_Gk(���K3xxtdnw�m��ԯ�Zh��tb�鈴2��x�N^ �.��8���H�%Cp/�S5��Ӛ���ZV��,�ys`=#}����̹^"�O�JmX%f�49�B���M����q
w���Z��^P2ݮ��[��f]�v[��	R ;�2J�;]�c� J��?oQ����� ���$����<s�OxI]�X��̻e�j�v���;�<M�㊸Pm��z*W5
�u�?lcs���N������y;������C��b[�J��'Ur\-��tc��jv������hD��P�{��������v� ����yb�c�*�rYY�+��_�\�o����+�*�]l�GS������Kh�Q�20���S�����s4ȰF�f ���$Ė�G��]��YK��@F(P]v
k�j[[�Sp]�pZ.���ܴ�&����n. �i�_N �d�0z:%��h����W�(�J�C�Do�ә��YV"��ǔtNnPR4~���5~`��H��>@iP�t�M���s-��~�Ӈ4�V�?��e�|[!������(��)5�\L�Ӑf�HzMa�����n1qW�����D�'�I빰TgA���QC�+I��ɔ�'qp��:D8a��T�X����h�g���T�g0�U�ҋr@�-�sGR��0G���}�<I_]��eKx��\FM���5��{�o����lT5w��69����Q=�d���A�[K{�Y�~��W�(��+�Rٽ �M,PA�Y�_��y����PE�AƦ�-&���B�1.+�j��������_E���ɜE5J�T�u��e8O�m�o���D+U�RO�W���=�]����G'����.�~�%8�=G�T'rwQ^a��I��iW��?�B2�E����[�,|9���%���9"/٣^�7s��< N?�����H4�u^�(A´���0�oI��z4�+όBܑ0s� ���뽏�P8���bǋ{��ثx�EL�\T�0��-+����	(�o;<vA�tQ�.'V�@���*HmK����=AH�"�q��i�!4?ay���Dha5K�4�e��%�.Rwy,m�S�b|_���][�|��ѩ	z�c��<L�_�78��!Cc��⺺�q.O�7{���⏦(���e��tM����\���.�\����O��U���]H��<�Cq"���9�u>{�6��Q?��ѱ�D<q�}-ڣ�(�ܳ�?�v04�'7�ke��Zv�Ai/�W@��y�k۵�:b�t,�B�-�уүR��(h������Uɥ�k5$e�"R�I�<���P��%I:L�YDC���@��"^B 4(��
A�����y���-`�g���l<{��x)��8��w;��G�����O1A��r(oϏ���Ê[&,bd[�-h��:8�J���갑�I�ܕ�~R��1�&SI_I��Y�Q��\{%��I�7�O��B^L�	� Ť���[F��3<��P�Wc%\3�@����,u:V~�M�Rc�1���ԥm9����C93�򵄜d B�J� �V~�)0�z�i���k\$���`���Ef���ɢن?�#���3"h?Hx��iް%�Dy�$�O��;��s�0!OO�{Y�EmKWg��}t�k�K�,���ƞU8}<
�J)t���ނXK_<M��h��|���I��V����
g��#�1}IC��me
��%���o�����K�"�ΛeRo{�%J�ŏ�d6"'S�V��w��ȧ�MDਣ��Xk�+�+nU�Yb1�@֞){�9�P��]�2��	r�wpKX��:ؼ� fn���UG� ��-���	�4
� ��J��if��8�V�Y�(�\r�"[�k{e�%b%
d�&�C�5ֿfD���}Ga[=��.��'LW��b�YԠ���옕պ�I�8�����t-֢l���33�8&Y�!v�&D����X=,ɰ
��+�3�T��!.�-b/WO�ܷ�p5`�-��[���Q�?���������&PuɊ���J�qX&A�.ȱ(�oqT�i!��}�$[�9�J��O8�/E���fn�#K��N�E�����Uf5�)��`F.�s�I�gϝ��ɋ���'C;<S?H�oǑ��&&NnF ���Uz5�zm~��^�k߫���[o�/�^�(��������t�wF���;g_�䢒�pGu:���6U��c�5��L��c�+_@i���$O/VT��u?oq�g�HqҨ���ܬ���ѡ�Ѥn��[m($�0�
x�ٔsT��HSk[ԇ���?Y�!TȊP�Z�:P˟��r�KV�}��]�j�\�����#P:��QΪ����_}bF3���� {L%l�=��h�:�����$�;S����ʍH��u�f��I�-Ԣ�4�[�v�cD����jN4*$�$aIu#E�`�]ĉ!0\ʨ����Hj(/��V/ȹS�����6��5aH�q� �%��T0ֲ�Ȧ)U�r�ņtS<Ǧ�&Ƹ`-�k�;Q��{�CI��눖�|l�7� H#�� ��4�Akѷh��0�ciGqڗ�ê(�5G�刬��]��5�����_�_�9���z�UJFX,���vg��J�+�|\�� ~��e���HG~5|���~MY L�0��R)���P�>��^��s<�Q����j�1��BW�Z�ߣ3G�g ٘`���M������-2>?�?�����x��b�2'0����t��fbm)z�qk?�����Gb$�H`�[_��6n���O��_�'� w��4p�d���p�.�պ��g�\{-����1����y��%|<�p�I*�)�uq7���G���xC0���+��( ���;ҁ���og��I#�w>1��%���cG~&��0��ݭn=�`���F�L�pq� �W��d���A��r����Y��f(�A�*��������u�%2���(�k���B:�K&>_x^!���P����c�â:������ԥqy����	����t�
9�Mb�r�Wn3qqkF�RJ��3K{�(w_�]�w^��ٱ�j���õ�mb�tad:CU�ܚ��0��P4q�@�}��F[Ơ�B V���R���+��6���PP�}.�$�*ՎA�o��d�l^�Q���Y��ka�8�_,��p����lV_�Zԑ�/{yPj���`q\���%B�%�0A]L>�}�@�6�l��@�n��ߧ�j���h
s�էo'�Z�Y��η��.��z�A����м�r;��b�0g���q����<]Y�v&�h�{�"���Zh-��}c͡Ҋ�����Dg73���c��^���`+J꾲M��c�������>���Gf�w���j�a�&�-S�1Bj7���O1�]D����#��D����5�L��|��JDU,����#@z�i��AU1�l>����{�*�*��|�r������p
~��OЭ��f(���?9�}���k��Я� ����)ڏ�\�2�̩[�^g��:��aMS;��|�!T[&s�[SK���P����`��8Xl����:㩝zQV�d9y�����2��V��1���S0�Qk�39W��c�fy>^fC��l��b.�l�@����Q�����xe�	9��ظ`�TI
0�/�A��%��ya��N'D�����+���4�����p�.J�vI&H�\A��/-<���T���Py߀�9��4�T����>�2%��s��,��%�Čp���&�x�@�a|���K�Pr��U��:�����N@+Ͽ�0v���$�TlI��wP������킍6���Yϗe�Q��Pd�˚�F8�vq�YaV�}�H�����hQ퍫�����r����p��r�i��P��'Ay��e���Z2<�0�)��b�w�KwGl�Qe�!��3~w���̹\�-��/y5�@-�D�~�_UcE��h�|{]d�z����ۘ|��J1�H���%���`�7�x��d����c����u���S[��5�t�'L���E�'gN�p�q���G��{�jJ��F:�����˹�Ap��pP��j���h�;�Ɉ@ �aG:��[L�b�H�F�����#R�u� �^4�,�k�˼������JOD3|	�	]�A��3?���#
wɀ�>W&��ty�*츗(�g�hxDU�fj�z?E��|��<�*�`�+�#a�YP
�3hn�����qeR�frzj��&v��iI��'�;,BcB�b%���\G���C, �΁�:�юf��b�4ɥ��O��_^�T ����a�nFB��@�_$T����r��SޕI�e^������լ��&����Ã�c�"�3:zƼ��N).�)�����c�Ovh�>P4��*���^	�b�̿6}����F:�B��.�RXxVi?v7'�
��	����Ⱥ��i�W��ixpt���i��.� �q�lw�0<x�ձb�Z��3�8�(�5�f� ��f�~�E�!�3�"�S���lp�`�8�h�4X�A�U�q@�nST�ʹ�gU>���������J���^!Wڛ�9�A�����F�!�`����g�g�!A��}�(A"(=w��U�=��#Az�q\#mj�LH��V�3��%�=r��h��a/Ԡ8�E�X������[c��j *WCy�tO��^Q�p�X��I���¿U�{A��T��mL��<�|�1��M���yJ��:Z�Ǌ�J8.C�v'�(kz�˵����ǻM˅����Q"ݡ��_��ȐCm��U�}�F��
��0��@���v��H,���/�z��q%{�4��6`U���U�m�r��b���jY�Db�w�5�s����g0�@($�������~2�^�:�%}$U�#�^=�;Q��~b�;ْ/gҼ�V�\0}Q�хB+87D'�(����8��B��k��o��k+l�C����OZ݅�\�!���SH�Cg���G����^HR�y9R�[d8��2��e�DPB��0�y{�s�[E1ݔW�R���\A���2�Z���N��Z���ʮ��|Gf�M� s3qFV�8?�h�֮�~��\��02���A��H0�R�����BG��f/-_�&S^H���4o�&� �@*�g[�{��t� =[�|K<�y#�_ٮQg�E�\L@����=��H>��-+2I� q�`G����'j�Y�z�)�eX'Ձt�ξ�������>t���n��ȁc0�]��2d��Jt~�h�Hbx�{U�4�1�^�;\�xT��զi��' �
|�9\ډ�o�Oyxlz~v?�am��"�o^��^������=��ݦ��V+�B}VV���&�DRmy�i��&/�E�%���\%j}�\���3���� [spI��M;�(ꞐC��5�a&���/2�$�X�J' �	a�ǔ)o�"��u���;j��l1��&��� p��tr��|4��Z�����w|�ny*�_�D�ݹ@��{��t۸٤��c���fGL���W�;A�Iޙ �h�c���Ù\Ŕ�;p�v� "���M6�!ʁc=ƙ��μ���Gp��P��ƻoR�X�?�G��M�
����z��nIf�u���	�m��_;u5�;ܤ�0CA�a35Y�T���cZ�m�vdE#�r(F%ʗ�N4�t�n7j��s�9��bI�o���\T���̟���7a�ͳ�I�B��M��޽��^_��A1��v�܆JL#�
� �E�|�x2��!{b��WF����{����Vg�%����o3���SR�Ɛ�C?)hi�#��@t��yҖ�i� ���mY��*�6}�� ��,zd?�O�8�rI�K�ED�Y����!Z���xy��!�����j��[�2��wBD���*����0W 8�� ���Ԏ�rjtr�.䗩���A`����h����9�i�%*"�|��:��?�Փ������*���d_�7L1`�;�<C��0���$B
]�ߛ��q���m�\P��V7��8R1|'�i,�aܫZsG�� �Y�u�	R��� �DJ�	�4��|1p��#�:���.�"^�္��K9�p�U���Ip���\)g{�芛��Za�\Pz�@?�XT����1S�x �7z��Y&��T. ������W�6���s��g�܅�������cZ��^h�P?�j�G˞�X���3.p�y@\1��zz��۷�#�#�v1T�5%lh�t���0 �m@�d)C)�nC�cI>��B!�Ί�$Ȭ�1݈]��Хb�u���cP��?N֡�0@rpa����D��h|�2%��T(�#Dg�
h�X$A*r�Do�F�g����L�_����93�{7�>7A�Iq�$5'k�:Fu���H,�o�u
K�D���N�j�	���{m����8(L??96?���Qx�҈�=�b���ǈt��{���f̚���B[�w�A5b�����j؛EWVɴ���|up#�і�Y=�%��[FY���s��.�E�}<ML&�Y]�_�)�.2�GG}V�B��":%@�]����V��g_�jiS@�w
a9��Wt�_퉃����}E�H"d�����W�o����	Ҳ�(����Z��������]W�lUKC�d�a����4Ę鞇ΈL'��G�E�ʘYj�/�l3���=���M��XDNDW�������eh.�w�����1_�mE��ٌ�}�R�ԡAO�¿�4��-��sr�y�NW�x�sq�J
O��Mu�9]�)��k}w��U��M�X@�/�1BjW�Z��O�ڤ�A��U/3(UN�s}�!�@	�>�z������2k��^����44ޑ�٪�L��༷������t�5hq�Lq�b�Uo����_Դ��!�����%DY���>|���+���}?لM.����=/=iHc�:j���!�9  cr��b��e���u}i�s�d֍y�W�����p/Ȏc4|�%7��s��{�J��+���c쟛�	}���kh��5����[�/�+�u�
�����%�0\�ib �~��?cc�����	f\ @�5�T8����a`��Zͮ�^�Ø�h�U�y�}jI�(���n��HhM%��FQ�����j�dfnUV_[��be�MM�-��un�N���� v����F��QGi��Ku��[Vr�C�c0Uł���4�`A#>}���p4�t�(x���7�zQ������nz��>V{�"�� ;q�
���.�{��=F���3��sʃ��]��}A)eX�] ��[(�֧���]�QW,A�|@��|ۭ�qi�+e	�
�X�IˣT����ֽ�j�6�S$gm�2l��D@|"PG��2֡CT��l��Ζ�e�{�l�({	�(on��^�Vm� Xp�qҵ�v���!�g�F���Jq��^��d^�xS�/�i��m�D� ��̨/��K;�,���M��L�ӕ�T�� ��O�J~���V����g\1�R�pdZ��-��CPL�q�r�(�m|�r6&Zy��Y��&��vu����z��:�0�ov��#� ������j��y�����T���Q
F�X����y.�-ݶoTd�'�7O�ñ(6U\2j���C�Q��C#���Ze�V��N}�@��%L��`=���>���x�ſ<f��3����~�Tx���R\L4|y��<�+ǀ�����L���Jw,�x_f��+�f�0�E�*F��E�( ��qwdp$��#='w���{U�g�~���\��t9��	�9��!:7:�SokR9=�$�(j�i�y!Fsǃ�V*~B�G� �����zӞɦ!E��F�a�ΙF�!�jeN��|nUf��kJ�'p|p%!�s��C-����n^���ŬI�\r����a~�>�3(h|��緈YX̯ox�\�4�C{��G"�5>$�h5Y�ӝU�a�O)��8D����绠NS�dS� ��>�<J]�F}rk����0��uT~賙FMmz����U_��k���������R�,��>O鱴���215|,�9��y��J�"z����镸� X�q�h@ސ�I+fݻ,|���4���k%,���;s[,?oΔ[�+�B�[�\�#s�s#�I,���-��GV/���qu�֒�5E�5W��.bVF�}�8�?iui&�% t��E2���7Uso��;'�8Fb��ʋ�9Ҭ?�A�r�kڄ �TɍP��v�ۭ�y���UE�7���p8[)�WJ��د
mj��(��A'��ؾ�M�Z��WP�X�����7s���:d��^���F�zѣ��3��*^��k�5�� �S���e��3$�.�b��zB�d� �D��dH��	*L+-�ي/�!��Q� �	SV`�L��b,I<�OeS��o#�I��ے������'���H4,�'J��[�Ԭ�,�x��Pi�wAh*�MG�W��I���3�/���"�w_��	��Y��V��i�"�/KsW6�|z���H�,*;�Dd��:8}���DX�H�RN2�͆@E�e�2̓\j$��J
���E�����	�I��m���'�i��H�PZ�8�_�F���W�!l"��!m��d\�Mu�E7�}%���ߧ#�f��T����ݵI���]��qR?�����������H ܼ悷�<^u��I�h_��a�B(���3��{Q^���ԛ���T'�[�L$L\�
���mݬ�E��>����χ$흋O�|�x�<��G���v��gm��U�"�Ϲ��>���ېR�!a�*�w���ѓ������=/���Mm�a����b_��+Y	]����H��%^.:CػT7k� Xizy/3���` �H�d�b>5��8'"�(@�J�8�Z�u��&l�n���aO����Ȳ.'��&�r�		%�p�n_�Bd,�
6��(D">y&V����sG���X�"bh�'�V�6J��8�̕�
�a�c���<�1���G}�}t�RC}k��n��5�k��@˞����ZQ3���]�?��[� Α�Z7�F �:�'lG��N�{D���P��f�H�~˒���2��dX���?�&+h��6����b�JI/_�9l��,�G��c#�2�|�Zn�C�tEN4��5�N��7,�U+ˎ�F��f;zj�L���m��T���"�ܙR�b�Iq�}C�=�
�˘ϣ����iw��#�͟�-\���r��?�a +�d!�pH$�fN�����K�e3��I�7�u��o�8��[Ћy��D�/�K����^~�#Ci�
�`W��?�ZYl�nZ�$_vΏ�o*�΍Γf�n8th��6|��tʬQ>�'���(YL|c��s�+�'K+�td-cB����!����Ұ��6}��\Ծ��@�`�=�:���4�5�*�c�r[V�l%�Z���t��� �)��:6���Cs;�`�� ǚa,N��p�a�������J��$]�"��6ƍ��Q1ӯ9d)����-��_#�\d ����E��y���]���}ꋭ���Gv�XY��ԇ���?�rzV�7��%n�����C< ��7)��=1�$��Ծ#퉃�u��`�c�L�z�oK M̶��&�.�d%vP��7i�c�3��t$*Hu��%�d�	�$�6="�L���`����j�.���Z<Y�fl`3'c=�ڔ���D����P�4f�2�D�]��^�����m5�
�hR|����Оx����L���oh6K �l��,�����H�`
y[e�b\J�@qU���WS�E�\�hZM��/w�ta��r�S0�w���,�q~�p
��i�.�8� ��#��jF��,k��e��{O�B�5��С�^���5�J|�� R�`[2��h�5Z�fW��'�������$E��}��l頬fW�oB�>�:11���1�/~��]����sgrTt6r7 �PeB�.�	�+9����Q�M�ĦH�tiws�Ǯ��[rJd��~fki�_�ߛ�k�OՂEx�<���pEX&]:� /\t��#�AXj�����V@������g`�N��� <��'gT�v�y���� �~U�.V��o�g���?��ZI�n�ؒ��"��g�6އ�E���]v`ʙ�������x�~w��k{���u�a��uT	�M ��
�[�A8g��Sq�atUWŵ�	*o=��'s?Q�� ��8�p���*F�!F���J�����Bk"�oh���q;�z�ٞ���굙��t �ї������mGeuLW�9���=��〬�����^�9]L�a���6z{�!�M=��d*��-cTj�<��Wpg���h6��j�H��n/MڌR[���.�_>��s�ԑ�{;�b4����u^�c�ݠ��}�'������ՖKf��O����2���$���q{��)^!-$��WB��R"ﱈ�+[��� �����5�t�3��a	��H��5���EP�ۣ?)�!Q+_�s�]a1�X����k�W"11$�u?���m:��)� HK�*�˃ӻ��L�;+��#r1VG�\|����-#�R*����@�3d�����E��@���;���-�D�(�+x��*�J(?G���,�*W�`�F�ZH>�E7^�OZ{���H=Q���İ6p�?�q�H^`���!	�|��$�T�[�(˙�n�t(;�ZVC`A�j!8�@�K3%4Slt��W��
;�������sv�R�_|�g�Q��Z���s��h��[E�K.3.��O�'~N�f��ѱ�:{KqF�nm�(�]c��R��B>�M�����*��r�|�*�^������W����xΤ�[>�.�|:�	��l@|(êSC�>��я1�h��UJCf�����c_����'�[/�X
8d#�_d���=��֠9���P�w�S��7b�1y��S뀍-ƅ�]w���*��˽+P_*-Of�;DBC�=�˥۝�	������_���Z���t
�\V0U��85�Ŵ;Mz�Y|q8�1��Q� ;���]���KTs��4nf��8u|ř��N�>Sc~ڨyk�C����U��0 ,�`@ioҋ@��X�Y}�NL�����m���*5|Ғ�}�7�������2�ۇ�<�i蘯��� KeW���A�������w�as:�W��&-b� U`��g��%I����XW���{6
9�0R�L�QW����uZW�N�ڹ?��G�i��3�Suc���\�שH����?.�z�f;ۗ|o`��e!�cAOf�n^�*_�	�3K&�!���e����!�!Є������e Q���ADG1��ɥ:Kd��z5'6������S~�0Ԏp���b���$𭥌6��X����vjQ��r
��H�v:�rB}�]��u�����
'K����a�_U���4�dAkK�7��7��|UH�&�ڕ��
j�Pb5vqS�l��9r�2���C=��sh�sRr�$*�Ϋ�"{%m��0'�7�=LhiH�:{"tf���9Fu���BE:8�"��A�%�qA�@��K�;��D�LB�)���#�������׵�&�'��(%��l23pȫ�&���3�b?��a�����h}ͮiS?�=���;`�_���ٖ�]���������W�i��@�YmU΀���KT�Si�?�����qk���6En�O��D�pE0� (Z��¾F.��pE�G}���Ӥ���M<~��1x�ZCEj�Gϗ�n��og�1^���pF�<$�F�ؗ�/!vF��,�et��%D��������u�&��n���<OCtD,��W��.�Y&�����+0�99 O��b� s>����%��!V& %�O�I�,z�'5����_�L�I���:M#�ywŸ��	�F5e_��)��f��� �Wp����t*�d������,�t�`P^h�uk�%��˶i��0kU#&=�
v� ��9?Xn�7Ck�;#�o��Ѣ�r��ܧr��vO�.��Cq~'k�7?�n�4{���{�:�B��`�V��-!���Ȳ��o"�ְ'�6TA�c#Z��!�`�Vf�(k��gq��#3��٣������]��7$w��%䤼��P"H��ܰ,��Y��$�#j�x*ۏKfz��7x��g�:��ߵ�)����:����Ff˫��؛�e��(�/B��&Զ�k�j�8�ѪQ������֡_��r�IQ��8:�6U~<�P������m�5S��F����{�Pkl�>.a�0���-�����fb�Y��f-��5nh���B��3��]E��"ԟ��Sg��9t ���6i��&�q8��� (뻜m�}Uv2��_�:�d��G���",4q�ԩ���j_P�t�:��ǎ�)�ۿN(ޑ��9�8_L�I�
"yq�hב�9�H�d�3B���7����?A�Y�y��S�-�+���W#�d]ȓ�R�[3tڤrjgi���`pLq�~��nX_܀�Y}���ᰋ���&a�e-�{���)�S�N���F*��{��)9�?Lx� ��{�}P�23&a?`����<4(B{�}�72�7P�0�;�wz�D���~�q�p�A����cqks<!�����gL��ǌ7φa'ņ9[W=���e�'N��$��|�߀��aJ������j��L�Px-�|'������K��=$VsS^�;.�B#C��|��Iƭ!���,0������%�m� ø!�2w&����hF3�h�.��B]���"���OqfTTҞ��9fO���,a�� �B��{n#����P�l� �Z�c��s��Z3�z�&�YOx�jt�Y0�<�)J���e)d�6s;�����{>�<��x]� ���g���c��f��R3$X ����%�<6�rŽl���Z�I�ǰ�E�@������E�1��x�?!������.�sS�7L<�/mi{ֈ�x�C�١#i�Oc���+'�b�1���j�/0q�6&a$b=�]1����]����	oZ�?`,j��[A�ŪE��}�	����iX);w�x�j�>���Cbڗ���׋I���g����*	�Y4��n&vb5�fX�4�)g�J
u��r�)Pj���D��hZ~dTf����1T�mi�\��v�//O� ����多O��W��o��;	?n�C>�j}�LX�R@ل��rk����ǆ@&�Z/Z�5J���M�7�q4�I	zF�,nG��w^~U�Y�ơi���q|�?�|�
���<�)C�&y�[����_3NA����H� n�,�R�ޤ�� �<�Z���Պ<�B�c���>U��`������Q'=\NoZ<-+7�$��{(5�3L����2~�ۮ�E"=OuӹW��_����D� p�������>CL�ɷG>�z��\^tH�R�&)��~\���i--�����e$��P��	aa@7cO���q�U� ps����%Z�MUD�CS �Z������$���I��UJ��_��M輸H��$�[d�K*������U�\�����*ش1���R+��� ����0�m��P`�!�%<YX����[�����cw���P^	�]/T��Zc���|�2,:EX�J��ؤ<��޷��e�������#�f\{޻�o&�۶��Ck⋩���ԂEv����(N�"TK��F��9�g��]�^�I�=kvo���կ�Z��]�|���X��*BSJ�z�,�`�z'+�Ē�6�e	�[�RF����i����M�M�0j�u*�n�Z`��]����auB�M|ÖA�	u��a�������n����M�/(Hӛc�|����˫��V	RDR1�E��~
�ˣ�,�DJA���jC�A�� �{�k��X�j�߭�,%����,�����#v�1+��*�t먔�3�*��Z��euL��U�i3)�\X��>۴Z����%�ͽ�ll�Ï��K)R��d�$�a,,6N )��[aE@H8�f����b�a�DmC�Ў`|�'�S{~�D�E�wٮ�uA}\�� τ�8to�1ș��
�_4ᨌ7�����,��Ǡlb��iS���-v���OhC��Ѕ�3@��I�^�7_-nř]{�,a�q�X4�i$(�%�8df�J�~"`���Wl�9\Y��6G?t�*%���Ș���pI8���;�y�C�+�s+?�����?fh1����<��v�d�v#��Z
0T-fP�C��c�8���R:�%�#��k�$�2_h�\AJXG/m#��&?"�s|����R��b���+]>.�%8�emJ6i|v�����K	��Z��o����h׳���[�
xY|�b����{��_5�'k����i��TX8� `:������nN���X��ϱ�q�.��2(���}�>(|��I�m���!�r��'�@�I��^G\����q���]9]�B�V]���ƃ����	{(������k�VԤYj��-Es�7�u�Iզ|-H���[o�ڋ�����i�U�%��0�zB�;�k��&��>�N���r�:
L�ڼ䦝���h�R2���t}�s�'���3�����3�
����d-a������E'��!U1~.��גM84�8�Z}?�K� ��u:ֵ㭁ڼ���M0��7���3	~�(�'�نQSP˷�wyv\>G`�����W�ld[s#!{���=�����.T?w����5�'����2����X��=�!Y��:#Gt0�o�0��wo�H*2k��]��	&(�0(�)=b�__K��DnEu����ޙ��ޕ�m��t;�l����qki���k�Iw<7)� k$mS�NT�с�w�it��� ,�)�#�� n�'� �D0��9�TD��;h��|����NWK�DM0�F�1/Mk�ţhli��u'�ņ��>Q���8��	���S�|Y��U�-f����q����z��E�!���.�l
�*{l���b�����&��<P������lC��������K�nE���;�0Dy�-j�O�8�����(��'";�
�,M'�s������A(%P�;�]+��_��'��Z��ش���Gދ��%r��/���m+�������F�H�	u;{zdh}�Z���y���o���&2%����"{0��Qb����	����l∴K-��E ��7��)�^�HS�I~�J�_z5/cB�ٱ���wFbj@Ifx�5�6y�Q�'��v�"�>��4��@Hwz��N������<�T���a��b7����{��AG�n���{b�N�d�|㫸)�
U%����eK��Y3�4�m����H�b!(V�s)Ρ+�Y����<�2��������~u1*v�����RH��!��<�y>������p�[2$�Yw�/�a��3���!�5�i��P�`L��s&�$n����4�w�?f�\8#�[=�X�ƻ�bW��)[�:�}BƑێb��
��\�PY&��;�A�txw^�ggN�������_���hn��M,Z��C�7�x"�G��C�5��[chc��#]!H������Cr �0�5���6Ŵ���
y�V���[�Vgl���|c�총H�W<�2����JCr��c���[lJk,��=�����u�	�|�:���?��&S���0������l>���]��?n?�ک>)h8*�.���Uy��p�v#@-����L�+��F}�����G���S���l�K]��˄��#�U�f%˛�eê�01*��{y��O��q#�9�iQ�m����tJ�� ��:�35�!
y[������+�;����׎���)�qߵ���.O}��Ĝ>���N��&Kr?�8��a	T��&E�%�M6�̎u�NK��K�d/��O�Fm��;y�aIO@��R��%`T>�qG!b�ښ0c�o� 5��Ɏ��<�a�����mߟ�rU _:�Ɠ�.͎��]X��'�"Xi�y6
�{�r���׊��d[�c�g�%1b�p
*ͥj�k;)�d}�{�۷�L�|�m>�y�fk�o��f)Y�G�}��sO��K:� ��ʪ�D:�SK4�(��/�B'���v�Y�и�S�a�N?�-���9t�re��+�f�OP�8�8B�󼢼�g����k �;2 ܡ��VZ_ˇ:���U�� �:�5�^R�mr܁_�gU̔��骧U�����
w�yaɤ����G��2��+I�{ظ�h���,����}����l����� ��9��o�@��=��3 >��JfhV�z"�y�u2A4���mZ+��jv������n4a���S[s�Mc�����=�zR��}�+�K=42ȰT��ȶn�'�U�w��dB~9�X(�H�WPU�'��a� ��Q�3G�Y�� WC�;���l�-����0�\�����>�I�qp�v�%%aF.��6P#���Ϝ�Tb��$�R�׸���{ %�e���N�p�n�ܷ����mdF��ʭH��}��eg�6���p͛+��7Q
�Z����%@��l�9ЊK�����`�5���}	�ȃ����ލ&V��o������u�����+R0J���*�S}�U_�}
��k#�(�Y�禉}uR*����S li�w���\�߲��%`��z�rB!�%&��ږ����3���+79j$}��L��3]k�������,<r�עO�I���ϼ	�_����V�7�����Y������P$U���ǭ�� 1��x_>C��t(���,2_�[�u��'϶�麏:��T�&Y����ځ���>�*��+���v�7�`f�n�1�D�����SLa}1�m�o� ��/�d'O�xn�J؆	��s��;�B�a�Xy]�>.�~�/�Y��"���.k�xj��� �;�n@U��q�g��*!A��	;hm�؅�^�>��Pry�l�)M�{�IB�}��������:ƣ�Ԕ��h�)iJl��KF����t��3����4�8O�'���������I�||������K�.��,�E�ƷWr���Ūw��=���Z!���Φ��(8��{�=�\c�^�3S�	�8+�X��)�w�L޲��!��7��Ep}��!Co�<s� ˑT�?�+�H�����4:va2���G��]V�
��c5-�
f��]��ǎ�t�{	��}���[�0�x��? y5�:���	��-(,:]Vh2}�	�^�g�W5���Lv����T=(���=jYdr/�yN1����V�������ڿ��3�e+�"�z�{�jߐ�=j�>�I����Ȭ�K���%m�y�5�����G"o�S a�K./��k����٥GV:lc.gX.m-oT�%?�~��b��C�D�31�|	�s`R�&#�a��Z�Ⱥwx4�w{����e�
;���iZݥ;=�K��c�B�����A�G���Զ&׷Y�ڴ&W�� JJ,k����ꅥ�M���o4��42s��od{�ĉ?���koN"�c�HR1��u�C��V8�����+��k�=��r׹��.��6k�紞�X
����?oWs&>���q�=md�|ZC�ƾ��Q��mR�ѝ����R�N�O��Ҳ�T��e%�a�4[�3�� �ܫ�3���at������@��~�t��LP����-d���~S��F�+�u���4�7%���I��J�hd�]�B��8>[�Q��6Z�1����s�3��t��E�;��W�]S�.������4�d˧���]w\N��CH��_~Muߍ����@1��xS�OIak���T�m~�Gԍ.^$*�\� �2�0Kb_�V2a��N�rj���X�HDW ��f~T��fH�I{ J-N6R[x�˯��Q3�5��e>�`��I򋜲��x>�/�} �i:�^���g=���ԡ�{����~x~�E�T�ɏv�p$�{�;�1��[?����i����.Jv�h����&�S*��Jל4�#��?N ��m򺮗�?GR�k��>�.�L�����{���f����]���Uj�o:�����\��f�	��:�l�o�91!��������?.��H-��1p� �*�e[���R��T-� �F5���j(��7�/���񁫨6��J��X���+_��(aHm��_<����dl��Y�A�?�>a��͂�j��N ���O>��w�Cc���rM�@�2����ǃ��nt|�0=F�U��U��������rJ �}�_�tn"Y�"�	��1'Q�ÞI���/��t�0g�C?2��\�DJ�yɫ��Y{>P��"�����Ke�XG��=��ZI��j�h���GV��|��-�G������7��觡	���bдv�BH]��^��N�$p�f�ꐀ�z�VD��(��;Y^��H��&�O-��mU?*t���R�P")��==��0�a=gb&�$4�_��_/5�CU��#��ݠ�;��a2����y�ͥ�/�5=bk��g?:'�b̓/� ��t�|�뫫s`���/FU�|�A���nk��֕���lQ ��=>8 U�@�_o���{+"��J�C�8��OtӸ��4:��go!�D��g�>>c0\���j�}���l�[�����w�ľ���n��)��Vȏ�[@Y�n�[k���cD�����֝��=�����M��G����{������.���x�J��$t�,I��%���{V�4as��K�I{��,���񺊧�\P��;�1��|�FaU���|5�B�a��&H"f��d��]ڽ���W�2� B�h������Q�pk�<@~w�}��|ۦ\W=�7U"�Mi~���K ���❧V�8����G,c�p̝���b�b���ܬV}g���n.�{��G��Ph�}�w{���O�̐1���x����o��W�=<���<���v���0vCl�]�_�d<� �&�&�m�ܲi��Qik�z�2�"d�+`Ɩ"K�I6����$X@
��h��'��;q��٤�(|-^�>)Jy�^8��;x�;�F��鴯�XN�T��eȊ�Qߩ6�{97�k6�;.a��{,m-���Q�[��K���@/z��ӌ��k�f7=:���r�S�f��RJh��~�Y�ٝ�1�Ѓ�ə�^�����I�=�l�K�_�,@��Ȕ���S��L#iRk=��g{*]�5)�&�2u����ht�t=�Čɦ#�9��/W[�����嬽����loPB���yoxx�$�%���Q�Z�"��P3[�im�9����麧`�F X�Mmgk+��v�i�7ˋ�х4�vP��yd���T�Ɲ�ZL�&��2(D�Tp��3����^�v{���Է��t/������B��|0��A�*v:au��A�o�� 0��	cn���Q'�G�ۀ�zu�ǧ���ۢ@VF�L�v�����2�l+j��E���e�����Wi��^|:���B�hM� ����q��	�HS'ہ�$%��V��Csk���m�ґ��1�?�ӛ� ��o�D�\�����Ϯ��`zQ�h>�(BC0�2~UZQ�H�~ۈ�쟟Z ��kSu:�ܙ����Dg�� ��w�I���w����-������M�*�dSv2����hs�F�U�}��}=V�A.��6O?����`�W�dG�2������pY����.��/! �E���U��\Iĺ�K��5Bm���<6Y��=Dy[����S|^���|�!�C�PMr�e�W��&i1U=��ch><ڊ!Uz���6)�,oƁhc��b#�n������Jt�}9Q�`�]�CA�����|��m�e�UK����(Q�~�"�iW.|�Ӣ��8i��p�X��o�#�p�m��K05���\�U\	U.k�	%�Ͽn�ۯ���b^	�mם���DͶ��'�N���n��<���V�2M�|h�_���]NX����(7`roސ�V� S��1���2G5�K/9_>�s��TT�������~�:�������@yS&x���l�)C����bc��Sw���u8�pѮ���'	�H�oM3E�Q��8�=����}"�^�XըG���Ա�"9�GN��T����o��w��Puʺ�RuC)&���ֻ�ᥠ��$�����t��G sR/���19#��$�j7�a��z��%xp&%�D���Y���}��xquy�͇|�}�3'���
�J@��d6�SQ�~�Q�������A*>��#���rvŎt]Ż'fQ��D1�fDOڢB8�0\8qN��v�]Y��NX�Fَ$CA���0��8�լ��Mǳ��;�"L��4����U�'%� �:>:ߙ��b�l ��U��_��)����D��^�{�Sϖ���K#��>�[�.w?�ĺ�Bmp��"�S;��9��;7J2�o�\��"VÙ�������R�]���_w;f�d10�៎14�M��V���t�S�!(w4���1��^�ݽ�["�GQ�Gx'*�PAr��X�a&�����0�(/���q;��гS �O|���}����?�׉�)6)s\�i��;��]6�/:�7pTkBSB��,���2��,[)Aqⶇ�?)�If��֊Mʬ�{�{mu�гX'��w���w����h)�[Ή���hD���kuI8�S�8T�z0�p�e3����2fZ�x(��������~���>~�j��>1M��۫u��j�+A�$� �)�E t�Ң�S
�u[���ߣcd>MJX��:w�7�\t�XmC��3\�^n �D��Bۆ��A�"hk��NdYr�<���y��0��*x���x��R�vi$!�vLL�w���X�3��_�u��d�|q2��P��*����
������ȱ�&��M��/��E?U�~���+�������]�kK���J�^BZ�[;��Lb�*��Sm4�?n������� �@pn�%[�0��IRx��h�h��%�r{7�'�n��qd�T����}i��Lr���!�	N _V�
@E�W�`�� {��r��%Pg��D3����%�U[�N�{���T.;/_2ޑ-�Ȥ/GX˰�-hc�%#��NJ���V�*������}��1(�~���+����� bl�q(V�f�.H�
M�3o�6��,о���	��������T�?y��L���>�����T��Bm%+j0O.It0��Zs���xP;���ι��C|����"؂��G�+e�te?T����܅ ��F�PPp�H}�G���<�m{������L�U�Z�`e������ ��{��E�e�Nb`�s��<_w�3�C3�<��U(��)��i�Px�w_��~Ds�sn*;œ�!�A��8��Eg3�vt?\U�����RO�ۅ�����U�hZ�f[����X�N�*Z����{&<���S�v���>�9J�Ye9�HVD��mb�7�e�����SKv0�H�W�
��t��2ģ�Cb�%�[i���L�C�>8OV�+9��fێǛ|\��KB�G�<k������㩄k�Ƌs��PB3��%�ps����G�-�WuJ3���\\���̏E��3@���荩^	z�:�T���ٯ�eH��P�����.ǎ���[��"�QcA!p�9�sJŚ���x�~�?ɴZ`R5��j�����$&c�2���ρR7�C��sW���1E��-�@�9�;HLTv�f�2a_R{<*�u������{�����j���S�����B^J��LU+w7@T��۰3}(
u�8���m� "�O�h�@�����!>ɦ��4OY_��9������'c7W�"�Z(z��U��#~�R@R� ����5[���j�ҏDK�B���~�q߽)i�(�?Bs�oB�XL���Z�o���Pwj'��P�~w���;w�G� j�GJ�>����6�(�L�g\�Y ������ ?�ײ4#� �=+3��m�\��?�w
�#-��0��Ô�w�
(����w���M��켃�E��]��s+�#?�(q�0NYr�bx�:��P?Īɝ�vL���O&�0'���Όm7���~�и�D�l����O�>��W4
�������+�ʝ�+ybǠ�+�}�iI�KW@k|��O�\��؉���C;��#@Rf���.�Ć�]<��[tHh�$�:�+��/+WT\�R�	����1-�l���⎑-�d�˛�R���I5R�Kn������m���4A�X�G���\;�T@�\AT4�YS/���b���u�.��s&���x�H��5�y���ϭ�-:�jX�b�S�����T/�7A�
��t3�2!V��O�Ǣ�?׈o��k�3I^�PN����wM��DO�P��b�z���z���9S�Pcb����m�gQ"|��]��2����r'cJ��}�b��7��5޻��K�s(2wD���]�ݙ�o���7Kp�?M(�a�A6�O	�?C0�:d�*->[;�$�4NAJ]�{a�68"ё&��"�S	�J��
�՗a�/���N��%��z1o�s^̶ПR@��ӯ��a�KܓB���	/��1S�� ஶq�a���Niy��~������n���g�X0�qÙ��
9�ԇ��d�C�n<��H�0��DT'�M�����j�X��aJ�j�?O;C��nd��*�A����L�!�0_۴o���T��oa�����n�9��ͱ8��fT+L��E"�@G`(�2�b�砦ǎ�
g1_З�*�W�o�;������㨎ntW2���AB�TU$� �C��j�fC~v�}��R֚�M_p�����❶L�(��0�(o�EĽ� 0!��\�1��=�3(Q�O^����㘻��M=7��:�@	����AߜXW	K��
���5"�5ԑ�/��o�\�u�����ܑ K$�etW!��)���	qDb�!"|"(�I轉V�pC$K-&�_X���vm' �5��Ϯ�����c�w�զn"g�u:���H��=��M9a3�'(��L䋐��3�d@|P���
���5�\!z�JQY mi�s���;�P#!=����K���D�5�*z�@�8uသ<�Eѷ��d;�a����(ZA1n�9�\"�Ð��.��?���1/�f�tӭMd�*�~�C?��X��V~4��`��,�Hq��2�&����[6%Y�����K����;l�a�%I ѸS�^R��`ԗ��J:�[o��u)�q6������ƥ�R\[��/i���E�֑������]�94z,E�e�B;��}k|=E���cN���W	������Fl~cJ���O~��:���+�i��*��UHh���q�1C�q �}�U9i���oVO{�]��Od��<s#�zW�xG¹��g"B��$�i���S(*��A���Qm%��_^����V��vEcYT�:
Z�ywL~K<\p
����>Q�(�q��� ]���$21X���#�~�{�n��LѪ`e�B> ����vQ����J�d(��s�M�} ��	JoX�R2٨zѿ��fát۫v��x�£����#M�o�g��RUY��MD���ـG��W+�a��~{�ŅY�U�����:�=������1���e�uIR5J��&v��y��w	�ƛ���dO�8#Qy��U-����U��)��EܙU��L�����I��B8���N�����lʉ3��V1�Tm�jcU��m,�1y��YK ���g�\z��C'sD�ѧm8�'R�N�Y�\�qTf8n~��i�dmDv�0�f( �e�-g˃�������"_y ��|��> ��¸u����A�y�=��&}T���}�W%D�6�'���'@�����N�K-{�k��u�tq}]I�1�d�8�g��<��S����
,}8ض�u���"�]JX#ls���4������F�N:��m��c!wT�x+����Кr(]�6&�t�(� ����4	��̫l�xb1�����U���5��`��ei���o?{x�ܾC~�����1�m������n�}G�o�R��zX>�J�QgAJ�nTF�	R�Zݓ.�q��b��m-l�Ʈ�щų��)���
�9�x}*�Gj�%�E����E�,��yF����$�YHKN�kN��S�W��z�X�v�Z���N�I=�y
w���,�s\�me%2�����g$���!�:d+����!C6�܋�P��޺��5nq&�2�(b#p���n�8�u�@�'���ǉ��/ T `c�{�G�Ɓ(4���p -f�n��V�QanvT���H^�܄'vl���	:�h��(	MV`�/,	��2NI��5�r���[a������q�m�I���&�\u~�l�|'���5�B��{QҘ��ւ�{�6�V�&\>�U;����ɟ���CB'�,��Ą�M�k6�ov�|e� YE"��N�ܸƖ�����ja0�6��
)�Wł?��z�ġmYuP_I�7����s��t���JR��FH�=TE@��Ѓ[��
�ɉ{�^�T
�U�MFd^�@f��{�Kݱ1K���u�]�������}��"�>mQ~L���aU��_���p[r�=������yF�ݱmjH5�L	�yb$�(�dH�7ͼS�E��K�G�w:q́��蠃��L)J�2)�a�D�x$�v��I1�;���,1+�I!P��Am�[,�g�b �fM��ֽ�����,��4���D�-3����m��UMG*r�أ�1聵�$�m؞�;����y���bܬ��?M*%N_�w��Ke�Ë	àL���A>�����麪��
ܿ@xE��k_2�K`�		$�9�P��9$�	6�{�Z��^�Dвz7co�}��h�v_m����g<tL)t�3 ��}�L@Apv�z%@��{�I�k��-*�J��w�y�TxZ�׶+f�ɚq��a� �>�=VK!��4}�t�IM�ˈ�]�w}�p���nmel,᳦��9W�5�_W� O�z��n�*]X�/�]��8�{�1}��O���g���J8.c�a:�����vC�NH%��'�n_
R0�,M7q�a�y���
.S�p��9�w�`��L��҂ֻ��3ya�s�jp��_ c���yŘN�}n���]�<2%Зa�Jp���t[��	E�ю�fr��4��R�o�嵢�!QJ����	3��M�N���=�b*��+��lb"(~�^�}�Z��n���KӔg���g���O<���J�\K�3���.R�W�WȢH�u�{9x>|����8�!���������|!h/��c����=��T���1��<�͹*��z:�v����Į'hMO�� �ܡyΰ�}�.��k��*�P�:<$ڛ��2�� �Rt�p�~�Ϡ�'��f�qC��i0˥؂��z�S��!Q����fs���P��JG,XY	ߥ�~�$:e4O�lV����f(3y�FӇ:�_ك�tyk�o����h˸�������6��9����ۧ*}����_o�b���,<&r���Ǻ��
D��}�\����[�/"���k!�9՗��s�EdG��/�J�w��t�PI;������qA.o�d_J�����
��ކ2�P���.���N�O��ԚȺ�M�,Cd�ǢT(�h�w��]ɉ�r�
S#|tq@�&��\� �q��H/`�ɶol�Q��q.��A���o#fZб�r�$ ���D_�������h�^u�7��DC!���M�qlm�C} ���z��Gڶ�[Yŷ|(�S�yi��� "Ɏ�$��[]��jFf�V+a��a��E�ݥ˻��A�M|q(��#�š1BF���o ��|y}\J4��vQ�R=��o�'�1p,o�p���Ǉ̼�hZV����k�����|��.��8@��(��CRC�ּF���g�1Kd!�V-lNY�$s� :Y]PL�����r�ȧ(�,�Θߢ��-zQ���CCxRƀ8�V��]2���aि2l���Tãʰ\w7:�e$*d��%,u�{�O���$>t�%�4/����O3'R�m��B0iH� �p��G��ɼ?�eo�~tdM�]��/�fD�+�!��/�[�ʉR�{�`MM��ְ��4�J>|��p��,c_ˣ[����Y�1"��^�� �TH�m����n�G���?�;�KあB�H����)a�~�>�ѩP������X�3�JcP`B*���\�����!	�M�ԋB��/����B��K�ۖ�w1ѱ;�
�'���JJ3���{�7�
-�^E�	�M�&8�'}����[��[q�xTi�i��7<��vs�6G��p���B�d/|z���ر d��vN�����Юڦ40Q�� ��Ѫ�P�1���'7��v���������϶ko9{��ќì�z�̪&9�S;Pz�ȃ�.^p+	 �T?@2l��k�X;��5-E��C�tU;��)��%�o����/���3�M�G%�6��N2��=Jւ�ܙ��u�|���H��d�L�F���'�����X�K|ʶ��S�G�&��~�b]pv&�|����b'UjFN�E-;�/�0d��ٔ�����>d>�D¨��p7�
��	/�2y0&�EL�/����('��_]z��������o)�`����BO��'�ĥ�?n�}��{G_��LV��`�-Ο�a����$Ǔ2��a)����&\�;������t������/#6C��b��Fz�45ݗ����\��@^����ol�\�vvh�_GZ<9x��b1����� ��A,�x���ַ>f���eva�4&�Gv�צ�U<g��J���ʬ�C�Go�+c�Ym���gݼ"f��$�0F�2�Z���=�a�F������h�X�H=��d�K��1�C����o���MnZ����\���5
�
������
��۰��Z/C��+���G�I1,���j�p�f):�MJ�'>5/�M6�N��Q������b	�5'm(��?�n�2+�� _��"���C��y�58�c�Y�f��et�M1b��P�ݸ���Y�lޯJ���,�bWE�2���U_���si_�Z�s��ծ7#���̌*!~�
`/�ȱ�ր�,�
��o��g�� ��1!v��B��~��P��x�5��z1S��Xo��g��\=D������{��Lw�"�����"�Oy���N�A�e�����< �+{�F�h��q����;�Ŏ��lkG�2'm�
G����:_�{i�8�t�����k/�	U�WL6`G���-W/d�f�K{���P�Zge,�^R�]�`�g������Y�9��-�Zb�����_dz<�y�p��j��� �ze��(�Y
����B;��_e��s.�r8cA����*�HH�.�fN��j]���&E:A$�]��Dȟ�K7.��t5K�M�f��E���To���a��m�7.A=0����U⏆f���C �w�q���d�THB���E��]֋�}��H��R=�u�.�k�\6�����ך?������\2����>����~�u"�����Ā��o
zQ�T�7�:z��G�5.�|�fx��&�@"S��c���l��5�I�,O!-���%X���ӏ�).C:~#���F��5bC�_�$	 qNxDy�V�5Ý�v����	$+�J)UI�k��P�*Vy�S$�β%%�`HM�(�~�ށ���6�0��С��U�_��IRK�<.��&3$��Do�����H3����A:��'/G�Z��|պȚu���|��Y=E��b��x1�|! ��8YU@�b9rp(��ҁj*#w �~��B�� +cEÃ��P�'�/p�s��`\@��$�lB 3�5�.�c�RS7�[s��d�p�4��g�(�.�%����`%NFɚ�\��Α�+�d1W����@�;��>���G����J�㒖����Q#X&��!������f����Eh���� ���M�a�|x;�����'\�|�0�����,�S���7\��Y	�O���p~œ9Q�qq��+r�3aa�L�*�! �.��_+4g6����Q�����3p�7ȍ�9��.�q���.���(�ͻs���߄^~�s�_������G.�A�K.L��d��qق�YbBT����`D�o�W� S@�*�l�<z��ۄ]��I
�1�xmsɃi��>/8@�֎��C��S�U� 0���1�����5`>E��S���|�^"sTh���g��OR"�H��/��)G��41���_�2H�x���$7��_(�i���� E���*I�wH|2.SW�����M������A�s��]�f�Zԑ咾�F7Ƅ˶��>mYE����5\�����ި�*�7���<��]���2�Xʗ���B���E���Y�h�����T�����W.;?N��*=�"x�����=H�Ռ����P��"��ͨ�dqg��Y"�e�`36�}F<"��UEt�0�3���ƲJ�d"�n��i�xq�GV��t�%�7�<$���"��Ls�b�*O��JX�-aa��K�V�}�ߴǈ����BUس���S�HOR(�F7���}-h�j>��#|A&p���hC�TT��NE\e{��K������rq�Տ��H� c>0��>�g��s��H*��N�㋃�y7����>��Nk��� /��
���T�FË��5|rv�8�ѝ*�H�s�﯀�ӴC�O?V��X&���r�� K7�kR$�}-�J�����z��*[a�����kY� �>���ݿ��,Pk/X���'��s�!n�Ԗy,�F$�l9�]bE3�|6!ֲY��5�߾��d���zY7�m�@�k�z�z[�)ڜX��
���^[w�?I$lh�<2%QOm�+�qk+ɛ�q�#Mõ�����t&���D׿�8\u���7�	�LwVq�"��`�
�=�$��ݠ&�?D�y��B��pSUh��Z���p����-gF5�[���0.���8���V��"ݣ�3�*�b�,�a&6�ᮒD����|�;�j�ګ��)>{;\c���?�!,/��B�����yX�s�8N�;g�"	4�"�����2��E^1����ߝ��y�}�
;����z=R���9Ʉ���ဉ	(��A|�f��V�o��;!`߮j�o#�_S*�@�+s����5�-�� ��[m�F����O�$K:.{��`��@�{�D�-^�E�g��{���e�0�FE���h��G��8��9�/_�����jp.�7p��h��kCռ�km����23yqNcrqD����)W_���V������P5�.O���U��?�c��ݰ�E���V!f�J  ��&�;�A_���;pA��~OO/Z7�y��&<m�!��,�A�ß7O�WU���:�ގ�c��b�&Bܠ��Ė� q������$
��1�˒�T�#�d���R���v7�L�ԾmD��;ԩF@�#2*^�]HY1rH�S�edc������ǹ.�R�����>6X�y��3�|��0�����$�wmB��u�>������2�)"F��u?�l�]s9���=\�I&ܧ�u="�kjN����7KP�XH��n��l����<�>WF�v�p(�'��Z1�7���+�k��H���R�cNPr#]���g�lv3}ʘ�KLa+�i}��L`��yfL�%b�+�lp'��=��ر1oo�)�����m��� q���P�t���Mq��
g\ͫ�0��BMy����'V��3"G�͢��[���c:ȿ
��-T&*l�J)>M��`3�
�"7��
�ᐈ�J�9�9
<, FG�z��� n��#	!�"k9�R��.N�Ѝ[��Bb�)���TZNǔ�������;K 6�uX)�O�_1]�0VO.��e60vL���9'�m�ׂ��@|ǿ
}Jr�L���I��^�n�B\��[���S��A��qf���g&r4m�)?;@9�g������U���+C;�ϴ��V8_mhs4�r� U�y�&ɘR�u���9X�H/"�~ɸ�>szM�0�/��Q���a)���)���V^(�h���yv�$���/���H�i8j�����2G�H��:_�T�į@�/Y#�MZo�k���@;_a�`P4����4�)w�TP��zSXV�I��l_��
��,�i_b�&�+~�]���5�;���Iz�J�'�G�B"x[�~	C��eNM�B��֋,I�/�3|X�@"-���ʳ�5��������>Blł�@T8�sViYH��`�o��6]� �PUyy�U��0[�Az��N��:X�-u���#� ���vmQ���a�`ۛ}Y1�P�@Րϯ9E��¤eJ��������"�x���"�X8���t�BY�w%��ɤ��<P:=7@�Ǟ˚@w�T�k�U0�{�N�Y�"�������{.�����,�*r��ϷgT��^�os_'�:�g��g��WQ,(�%��1m�ƅ�k:��˭y;�Ռq;��5To�Fn �ũ�m���a.{�׀��{��=Z�7i ~=S{�t�\��A.Y�pX��j���F
Ĕ
����Q��"����% ���!(L�a6a�,Ёf֜Vg��{_@<;/Ɣ��4υ���D�]�t*�/ՊL�)�(���M�gWo�V�v,rBc7>�Uek��*qUL�Ҡ����l$�6�j�����qijV2N�kC<����h������; �c
�4CJ�wd7���X����}Y�Pi)��� ڒ��GS4=�.;�)�JV<��_�5ʯ|�WO��R�6z&Kl@��i�o�(��*�d�~g���`����[����tF��x��O6�G1+,�n�Z@Hn{�jQ�s�&�U%	�4�ų����c��x��S�5 �ti�����x�C"?���%�Q���u��xҷ��dj/�Y��[ڔ�Q�Ez�"}yO8F(�2��ފ� �
__��#���ƴ�6M�"q6�&x�܊�:r��lh�f�y�vun0pM�$Ʋ	7����Hv#F��z�L�C�1��C���l?[��r�u}��ZY�̀g�Q�k�v��	\�2p����
������j�ci1j�͈Yo}�����r��G+��0�f ��*�~�[=���B/}���]�����2g�ΡS�Οb������ٮ/ z0"�����`�z����J��\��4���S�&��c߆��q&��v�7Ϊ���* p~2� ���!Q����aQW��T�Y}#W���FD�]��=����f��E����9e֏�3�%���CM��aʘ;�c�Z�s�� \���@�^��
�wO`��麐+Q����°�Z�`㶢p#7x�&(�tQ4k"+�0�6+ޗ!�^���(#,	�m��nN[A�BUC/��y��	�-��F��y��\~*6��UC/|1<��WtF�������a�����^v: %Wz��X��c�~j]&������x|U���Q�L�F� � >~耦���J9��~|����Ke���p�X2\)l����
r�}߶��!E3f1a_~���<� K�HO�N%�d���n�왵8����7B��GK��|�qr���C �yf@%�����Tv��:�K��K7���aC�%�#��)x:x��/4�R�j��h��ڕ�t��YmKQfg��k�n�&�	��%9�J�"5W�R�O�J3h�/:%�
o���S�ǋ���o������/�blë��"̬!�&VUP�Ɛ	�&��O[����G��
�^]"�:�^�W�g �
4� �7	�5*&zg�#%H��{�W�ԷZ�d8|�K�odҼ�3ܳ{�-�s.%�C������(�ÚgY�X���B�8�V��P��rOT�5�_[�c�;�z0�iQ�Z��]���|0L��[ݞ���Y1���D��/��iO���(路5��P�{��\	�%�o�`97[����'�g��[8�`�&���t������	N� ��}c1gw���.�"�U���z9@�мy�7$�^{!s]��MK�M}8�\�QÁ*�L���(����?(��AK��d���@4���<ndi��7]�������Y�:@��)������X�/�rZ��r?g�s����VV�$�`���n�y�C�LS�>��J1��]�s�gܼ`�̀J�����^�hҮ�s����L��k���}a�Mu��>����|�3P#��:�$�}{u�]��4ISp��b�����y���0�5�(��I�kE�l�Ġop\␪��G��B?'�Ē� =ѧ��&�W� #%qM����m�����:e�.��M����L{cxG��V���? y�
y�d��`��Ͼ���V�p�J��$�i�[Qd=�����l�l��bj0�`�ut�KqaZG�(�?�|8&�KOؖ���r���X��6b����O��h�)��� ���^��E\�S4S��K��7�Ymwٚ�^Vخ��v	Q�(E�D��[)c),{P���P���b]m��u� �.^�Q~���r��+x���i>�Q�HW4#�}ؑ���;Y��rWu�c	��Jjn��ۣ���x�^��k��Z�{U�o��˪`���_ �Pw;����2/�Н!s�Z[(�qu�Z�d�2�T���������6���˫u��iX���ơ�o�*I��_a������^Ѐa�6#����!P�I華�Ѵ�ț�>q����s&Ty��	I�j7q����U�	�/k��vemHM��Q�>��5#F�d���4�#B����f�m��c�w�3k��\�dבP�t��k�P�?K�M��ͯݐ |u./J�$���CxՕ�{��&�fb+���
#�4��Qy�S|]=���X
�v��X�O�J|W�*Z��2q�;u���������疻���J���7���^�3B��`��42����T���2^Ú
��P,�<�[��5��MjW��&�Sڏ�R&�B�8��&�-�fpXÎ��[)�_N�eΡHC�"�6L���i��5�����tu����6��Y���]ƙ��a���?Uն��d��
���S�{�'����͝����q�|����
����	S�sw��ܴ�hx�����EJ����A6(> �2������9jc.g�������#o��*�{��' �9�6���k0T�����F�A��ECH��GZ/����qI��9z�˻��;��> )�۬,5"�9���ט~�ͺ�}�~+��^}��W:����K��HR�k����rorQ6�v}����8朗J�c~+�;��l���v�6�����Y�t��W���K�n/�%~>�9	�ѨX/ץ_�4h�a�~<���%��i���y�N�ӱm��VEy���*ţ�!��1!;+M���o����*=�A>�,�Q
y�� q�܅L��f}��:��h%�,ͭ��ͦJS�YM�xR��TӸ�[���tlh�=p*dH����9����[t.�/v���/�I�|�(T����$�$�K}��
h_�����zf��輇e�����\upf^;�(Vѱ˼1^���/����Dr�=a�hq����%΂����84�/�'�^9�����*��XA^�m���oT�1]KSqcY���cӹԱX��#k�ii�9c�k[�o5c�;���j�;�{5$��6��͵~�oi�K��:��CH����G��#lA�Jt�N.
X�)Ռ�V�M�EVԥ��QQfu~w4t�=:��RӷC&+}Ǟ)J*Y�hͻ6�w��m�{ުt����~�UC�أ?O���%����'q-��gJ���-]>/_8-�ao#�����ǚ�el���/D�	�Ԟ��[�=��M�6�ّ�G��6C�| 1)$��<"hm8��\�e�3�jcr��t�m�UP���p�H/0{�/S��� ������tŒ����x
�R�U�i?� 6����R�����u;�˙��<G��<k�`�d�'���d�WI��,=�45�'_e�R0	����,������y�C�-l(�[�\74�0Sb-�$5��'҉�`T�ܹ�֮���*����^�^�Ǿ����ia�s関o���WW�v$[��>f�N}��Xl�v���J2����4��"y��(�B��_�\N(����x}uI��u��0]f�x��l� �>	���B�߿�{<��ְh�FlS�Ѯ�1��S������d�"\���p_���c��nHg R*{#��gN�Q�UҐ���%� ����&��5Qj4]�;�EQJ�~pE����f͇Z��:p*���Gg 3�5�k�d���#��R~�Ρ~��\�@>�T;,|э,-Y��*��`����}��+�6���&�;ih�Qm��y�oNw�7���U#IO��MQzA��nuw-u�!E��<��V]R�}EJ3������iu{��+:�f�_JD�}�M�����s���{��������/��y�eV1�=ְ6�� *k���~�7o�wy��FE��(�ÿ��q+� ?��Wt��~�l�sGٴ+u��,���}�`.�
	�5�éI�]fi������0�
d���]y���`u�B����QJ�}����sը������x�M��`��V!Ũ��¯y�vv�+��_;�
R�1\�5=:Ë�� �i���÷��7��x��D��[�Gh�&�We֊b��?#C��Qך
��1V�ϊW�<���$�UH7z����敼C|������|{t1�k	�WsM�My2zp/�;Oc?B��[��b�r�OC/ͽ��\~��lQ����J˒Vw����G����S�/B9��TPt}W���0#����$s�.�Q2�h����>=����G��`������Ѓ����..r���a8���)��1���"
cD���d�L/��`[�cސ��Kl�Ο�`�Y���f����y�e��!��|le�^�>���!�n����� OVH���l��-�Q_��o����9�>��H�b�(`�ܥ�������)ݽ��jK$"���LE>�8#'��0���}�����\vP�	ޜ�8��]��
�ŧ-=�$�Ug憙A�J1�G"@,����9�N�1%!\��� m�"��})�
������ŵ��L�W9}X�W��� �>䡐-�c�E4��������qVI*K�+B�PP���`Z��-CW���q��H�X��9X(��6�U3����'&Q��uo\�x:�`F��W�xK�^i4�i��V��{��D�H����fL{�Lۈ4������İY��Co��H��~�I��(%b;�Ư���3$4�]����0Ɋ=�h֬�tG�t?C����~�%��Ș�,��J��~G�cZ�Z�Hd%�2�������0X}d )W��r��I�����!#E�>|^��;��,k�>UA�ݱl�{vY�{F
��f\Vi��"�0t�F=#�>u^CY�?r7щ���`}���6�+������I�ٜ@�C���2N�ŏ��J'.Q)W���v�s�(}����A�k6)!��x��޳�j���#h�qcq�r,�i�N���A�Eq���x�R�)k����������'r�pOe/X�i]�Z��c5�9Hr(�W�˗4yZ��˗���eE��_��wrv�K�?~�:�|D��X�T]L�]��1Ȧ�-��>��	�W��q���g_�,�I�Z�Y�.���nL�t�_(J:K�°dҜ���u� �E ���}��h�\c-�&���i��9b4�2o])<�w2ײ~����cR���f�����L\q�<�Bw��0FpA���4f�
��
���̝[�{�&�w�Q	Z�%�Sq¸�k]4�BN�Z4x;�ʀ?��`�M���4�O���q��w�u[0� �9��#��$��D@��Mo)��#��ca�]\���Qr������
��4/7������ ǰ�LN&�~4%��
�fsP5�JDB�,f�[Awf�0bݗl<-sns�>"��Ha�ꡔ�@SV,���2�����Ye_��5
�q]&dO��ګf<�^eTQ���.�=Lπt�G�Ӓ'��8Nނ@ޮ}7H3�1+�Z�NI�[�?�q����_w��a�&e]���`��	E�VNƠN���SaOvA���������I�3N���x?���S��T�u���|��W��(s%s�L���^O����� F���f��{��&/m�,ٯ���)��.�^����;.�	�4 ��D�H9���3�P:F|��,�K��:�mjbpop�cE�lT��ၦ���Zu��k�p��M� ��]���l��a-��~��jxX�S��N]"1��MI�~j'.�f���� 7ї|6�(��6�3E�Q>"�De��I��3g*cךK�|�h�}rYU��H���fW�D��QQ)	]2�#�#�ٝΐ|+����(g���F�v"Вss�&&�W�z75��M����Hw�eĳȼl(|���C��
Y�߇�����#����p�~��d�kio�����?����5�.�S����H9�.�K�\�����6pH�����U����9,�Mg}EY����ڪ�"+Һ�
�Y:t���F��mI�S=���j/ؔe�歩:��XN���}�~�g^�/����V�Ҭ�X �T��5�S_�k(�ħ��a�ߛ�׹����^�$���"�E�J�ٍ�-C�X�<��ÜZ����=�^h���ʡ�£)T�ֱ����ٺ@�\#Ԉ�ƈ�&��Su�Z�f�(=6�q- �*�k���� R���6��:�����頛�u�J[B���eȹ�&Fǽ���pky��`B�+��ǚF=[z��R�̽�9s V��5���mU��}���z�
y��%�I�1��@����C2�"#�?��3]`>`y�+٘$���0���+�l�ɜ�Cr�+!o���9�$�p��&���)���&���<��t�Z�}����i�*�����/)/[���*�%�V�&�B��&�n^��C���w&Ni0$hp��k�������Z�bU��:�8�l3%m����WO}I-�r��&�;2|��cp�<��g��.�����a���_i�X� u�S!)^:��A<��bE�*s{�GGZ�yC���zR��2Sw(�S̽NU�$�0ń~�%U?�S#z��m\���S����gN秩����G%_B��sY�J��X���v�Ji���e
�����c[J %I,�[��hG���^5�%������o��������O�������-w<�=���47��d�̖>�5��CΫY��;SA�d�f���\�P7S���u>]X��Dz�[�IY���g�_en��Wp�=�qkC�p3�j��N� �c8�S�@�L�4��xWܧ�*Ɖi��=�?�s�+�����1������FK1�D��x�; ������z!�ٶG����HK�3*��|4�WW��35�		Vi��R�V�M!���P�~u�K�DjH<��/ͻo��|q�ʏ���$��;�]}�qLȨ�� ���~Q�%Fy��G�ȏv�S~DX4���o�d��]�YQ	�-N��U��?"RLu�v9�Ȉ��	�E�T��]��Х���l�Nyr�?ɳ�/�K�?F˪�`��P;��[wp"�U &��	?���*��*1�%D+��.��ݬV���/-�R�i��f�nߦ��Ə�ܬAt6
��#��X_�lc���s

�.��R��W�峤�U�(���TNׄ�x�!'C߭��r�����h@Ցsv�'���\�=6�����e,BM5�Sq�O5W'�t��N�1������]�l��
�W�*�%���i�����<p�����`��Kz��,�/�[��"ˁ������3s͟F����d��l,�VzYz釡�|��)����Z����Ӯ&Z����V��c�'Syd�O�F�v;��=�((���T�g�"=���BثN+?v��J�xA	a��c]]ޟ��P���J�`�}��Z������3��7������Ҵ�ư;�K�#�߃i����h�}E���ti~�F�Z�D�������U99*����� �;4���)�rf9��(b��P.����U���J>{��|����ϸ7$�B��� �3��)t��M����U.<:�2���KB�N-:��Iң%	]E�t� co`�8}sʤW�4����@4��	���_ܹFJ-8l�Vy��_��S�Q�8R�/S.���_�{��Z2�/9�n�-��J�	wh2�
���U�:6���{:Q۪$�W��� ��T�؂i��ww��+�.p�zL�56a�सNI(��yV�W��B{zC}b��/�F��G���0�����Z�遹V��p�}ؙ�S��}e�V����k�/R��Y�lՄ���[�o��Y��n�Z+��Nl,��(��N�쟆8C>h`=�����h*γ�����A۩�O��+c���.�o�Ҩi�+8<�Mj��,+w�gS+I��GJ��y=ẖ�8J�js����ɾ$wyI���M/���4?����"u`���F�s�x^M�~yG%Yx$��.JQ���/�^���PQ�j��>�@̶���A��/27{@�M�.Wy�x1�O�h����;O�)��ty%b#�t�h��S��Y0U��?wA��{#:���o�����#�d��O��M�^qF��*<��j�di�?c�C�F�F�1�{``�	{�co~�s��-BB�+���]���MX	k�z'Sq�H�ӖD���˓�p�}i��F�Gj@��eQ$�qB��S��D�>qsEu`���@�������}�)�����rE�at� A6����c�4�'�������ƕ� ^o1�x��.W�p�v�=�s@�G7X�};~/.$�"#=�ؠ.��� [���9��	W��1��E�H�C��<XJ�i�9�l���H�a�X7;0��w��
������������:Q,H#֕UH]j�>�'0U��5��k2[\iR����%~ZW�D�3�������a�]*��~$����0����[)&��Q���sfX�%̄8����33!�o�����܆����$���W������d�t�D�xg��Z��O��� P
���_���+�������G��H��o�}lC+9��g�X�X;;���/(�=�Lel��,����<�z�>��֕��V�z� �W���z����@2�o�s,�;є{<C�Nz �δ�0���^`��	%�S�d�XZnC�0�u@�)�j	�$/�8�#7Yf�3��3ݩ���!��5�״�ېJ�(�"Q��)��;��~Ͳ�.y��N)Lobn{�^XzIad��î�������b��p��?(�x�w���<�=�Z��׸o��V�#,�<uS�=�~܂�~�%���ӊL�"�71�������I�0�}�-[�BΨ0��ah��#�C�����t�h��rI�J�b���� 2�~��&��<궞�����8&Q�Q�q�B>�;��G�q����jݸ��C���(zO���n�t-�#�Sմ�ݠ�NO�qm<KȖ������멤<ǜ�@��h!F��[�1F�!�i7��$+M�R6V��\��	�rќ4�j�N�
�	�)�Q��eН��O?[j��he��u��	��a�E
���a�9�����ř�0��~��	�J�1`0�R�9�5j�]�*��5D#��/����n�`�mPxUY/F��P�.�X�'���D���x�O�V���Ol�£���;��a��{��G��n����W'>�L�F�6�p�x�
X������!�R��NJ�>p��RcNh�B$vn�#�L9��}��	i��	$�5�����y�$�U}�P8gpxi�f~{Q�5R��?Z��bBG^�mȲ�Ja�~����U��VQ5�C�������z�C��n�(hP���V�������f�Թ�SqoJ[�����@J�~�P�eƖG�¹$���M�D�����ls�y�zBޠ�t�1�9³R�[F����`7�a cx���XR�,�<�W�N��.?
yê�̾�l���ZM|�&r"u�J�_N쨅��N��P������Ɉ���qH�I_C��m ��[�h�ʷSܢd� m<a�3�\H2h�n��a��JKۿ�BKD��ڃ�8e��]Y�x-���j����T+@>n��E(�F�@��!+R_g5�Z�N���LR�Qz�Cb�2z
F�\�F�ʜ5�qӶ8�p�#%k�K�0:\�A����t������ۿ���
8i�;7�ϾG�Ծئ��`�V��СD6m�El���_0��
���n5q��s�4�1�B#E��M��Fm����hul���d�������.��m��Z.v����ρ�|����e�	yN�������_[Z"�.�:l��/&v���y&v_���b���g�SM�qa��ޚO�r{����!e�0{�$���e���ߥ��yuL���]��B�M��y�eǃ�rΖS]���gX��&�Ue�	a���
�2��i�(�p�Tq����+)�IBd�a�k�nEW�?C�n/��Y9V����h���a�;f�R�L�Q�
.�� ͖��p��Lr������J����2�>H���.����v4���`�d�T���X�By�����z�
1�Ŏm=a�h��G� \Ee�㛲�AG_�͞t�j���[�3����m�hI�7���ymG���ܐG18G�6�nc�����A�dP���^C�5���_]ǒ�y�g)�.ڬa�,Hd*�10��,{	>!�1�sh���5¸�Mȹ�����Eֈ\���m ��j��i2�d������ �)�Rl_,�/�B"���{b����nu{�r��h�qU�����[�t�x��b��e// R��=9Sтv��"T��c%6>�R(l��z:|5�k������NZ�$�oS �}�W�R��;++S�`TV�o��j=� !|��G�d�ܟ�~眺8�P[�OI�CD}�x'���֨��8c�*86��8�G�A��Ǆ�zoG;h���s�����/�A�2�KB� �xN�� ��	�pP��bl$� ~ơӺv��7�SPh�] ض�u�3�t.^�%���L��K{6B3���*�lЕ�G��DBj�7���n���xu���n{M�i�r��0�D�U���E�#0���y�{'��d�\�@/)�Ԩ���!0���Ѐ,�i�^�~�s�Pu��l���Jan��b鰟V5-;g�_{`����N?��8�d<�k��?��������fL���R�@� qd[,�u4)�!� ?a\�}�h�%��}a�=���{�h���7������Ӆ#PF��ۃ�Fp@��΀�;SaiE��A�����BCm�
)<��օ���`M��y��p[��s��L��gKtu��S�u9������[���l޳˂�Sߥ���_�rËΪ̏�VQY�6k0w
ގ� ��
2!�h��r�Bs*h�(�|$T��m�:z	Z�Z��^���=��L#���s�S�ɲ�K�3[͂T�����7��5�nX��Hy�QN>��j�M`p���2K:TQ~�E���*K�&�<p�_��ΖȘ�yH#��CŚL����%6�3��X�J�����K�L`����.���FM�.�I�����܏�%CyD3pSe~Z*�#���������_�F]��c��	L%\j�Dd̧͙���pV7�ၵ���\_������9.¶�ϝ�?�㋸�t
7X���D1q�F�zhc[�ͱOuލ<+r�����/K�PUq�E?���Ov1�|$8E�5�wW���~�"r��)E[�&�����ߡj��G+Pv.k�o��O��C&@kmVc�.�>]389��_S(��(�=���b��Ӥ[W�̤.\��7ے`F�p��w{���ݷ�4�2�y�9k���>�u|k��Ww>������S�
x{�}*��X�Ln�ڬY7t�>A�N�,�����4�X��/'p
.�	����T3L̀2��<ȹ�N>�;!��d���K��'� j8�AtaN���9~5Y<���&�gG��"3�4K�0�no�VK�=���XJ���Z���]9� }8��l��H?L����
#�g ѫ�'��_{|��G���ɚ{��s�� e/{��`$>� Fi��8��?g�F�1:�/\C|)��2�V�W��	8�[<Ӎ�G]��B�G1����.lz�T�@�A��3�&�v6�6�s��� �e��%� �W����q��b.m��vJ/���Ǉt����ޠ��H�����t�&:��EpF��׭AV����5L���)g�����mz�0+|~8�J��t�a��>�i�������GH�N��"�9ѝO4T���VB�2{��u:YlB��7���N���| w<�~}D��ٚ���`�K;~ޞ	�h�/{��Z���j���O�aU�#�0��z�Pכv�f���WOg
����c�9���_�.*��$F�������l�-�dt���F�����?k�ǫ��*]�u�����O�äv�vx�B�Z�T��������
�r�X�\����0���M���`�xE�&u��,������K�	3i8+:7"�"�IG�Z����D;P�r�֘V
Jۙ=ۇ���(��F,b):���@x���=4�1n�YN0y5-�
r��N��1;]��~[�{�Ԍ�j�;�����n��>��gvz��!���c<.;i�^K��Ė���G���$�s�t�Z6�˔i��o��d�͝���Y��	b�=ur/��,�52z��υ�y�0�6����
�(�E(�A��~�`��BX�'��P=�ۊk���wy ����i&.�` u��i����(5x���&32���+���'�h���LH�tSuץK6VN�������ko�g}g�ϊ>0n�DVTW���^����U�d�;�nA'��]�a���(׏��*�$Lߌ������h�o�9B4ʹ�H��v�'���I M��fMSFt�N+z�jRE��u���3��$s��~7M���8�x��1,����KNT�����5풀��}8�8��TU4G�/7��z�W�%U��S���ڿ_�lPe�f�"�<���G�\��8��u���a�3:Y�F���Q�-��$�֞;R-�>�=��h)�;�9�}�$�<P�� XZ?2�bM���Q��9�^�^;�`�9�O=���(l�F~#�Q�	��80�;�%.��ऽl�].��2�1�Cn�����KAzIyQ��n��Ͽ������}��V�_����R�X��.\]o�׸=Ǫ�/@�7�����TBS�:l��$8�1S�~Eq��~���H#]�~)"����9֙gF˨���p�5���Z��U�yס�Ф��j�yDVx��@YU�z������u�NB��.��N;B�9��ۘ�  1�� ����{a���%{��D�
���.�?Y+,Yw�������#��YB���)�:Z�	|��8�
��e�r��9JlK�V��g!�j�{�9�9����@�j��?��l�=\
���$zKF��w��~�!�au�eۻ`�u����W�����>��}.p�u���%�Ҽ�V���4>m)F�%ބ"�2y�O/�Y@�c�,"1�ȵI����e���x�?������xT�^%�i�r�����?���8��/G��,&Ȅr���WFM� Ƀb�i�y�r����J�Uu�͚�@��qtE0*�+����3�f1�����L��`_�rJ�N��=�b"�t�%���ɱ�_�Y�W�Z�~��_���ˮa� �]b��_��}��ň�|+�.�&����a���9�և��K�lU����&��5����]�4��`NA��O�<�¿�E���lQ�l�C�:kcm�6�[���;s.0r~�)��ڲ��o����;��I꿿��o�`�CX�oT�&�1�nqژ�V��x�>邋��U�KIV���E����i���~�6����عQ���
��Y��d�c�b�W�@�ċՍ��5�I8�C�����y^��*h�Y�}N��\ɨТ� .8�����t�S��a�7����Y������U�=��\b�܋�;?��x���M�$���r]�p�Њ�}�D�\St�;���	�nzm��< �c�u:��՟����mL��k�%����Iȃ�j�|]dLD����O�ٔ�-ӯ+B��h�����D��#	.n��<�f[�7��E���{h���Tx��`�1#ܬf	�>;�ڳ�KR���S<��"�ktۃsŷ��?�G:���9=h�C5o�����x�qu�U�=m�\'�Z�׃�י��Eʹ��������7M��?-�/R>����~�zt�����Ă������`��/�|ė��q��)�'	�dFiDɉ^,���������s$�C"F��U}������������5���a^� ��K�qsL�� ��v��\^`��f}�=P�B���p	Kܜ���0��*:���d�O��Ҳ/&���x-�bÝhalsts� ��w>@!:H��-m����ʚE�;b�G��RnoL�Hxd�#�����;�M;-q����N��#u�j�e��?#�`�6�P�3"y~���o{�P�� ��(�(l�B�{�oB��<���{S��$�`g�`��AMt���C~_	�:��|�u?dn�|�}8��e�{�M�V��m�g�~d��]��w5i��`}�]N�8�O�nC�»L��+��1��$l�XDW�@�g=xX��-��\k�.�6��/����ǰ�M3̓M� ���YG~و�%`;g��&�z��0�#�T4Q�`]Q6(�b�1"�"��#���R�'关�۬��ue���M��5/�%~p���i�i�%	B�i��W��0�As�)q�K��x+�Nj��ZZ�/�AQ�kN������u���-^o,Մ��Nj���]0��5�^�F�J�ؾ��b��_��vm�H��o�i9�8���H�
Ok�#���"��@�^-�	��b0�\I�|�J2����3���`��൯iԏ�|*Td�À�č��'��,�4�L����� ��v����D5&Վ�I��P��ole�5�7���tYD[�b�j(��K-2��;��i�'��<"�QD��=��`�+M���2�f>�I���X��l^V��u�a6�s5�s翤����K@ٽ����AqFZ(�K��݅8X��Zw0�6�j��WH�x��O��@��9�n��a{�Hv4�bo�3-�e���b�,�|�Xe���}��ٔsk��(��S���ڄ�/�XD����� �C��5�2��!��=�B+zfr��/���BOk8 ��#j���'ٖ!j�_�%�w�zz� �$-o�!�r����Yl�!(��ū���Bh�, ݂[95�â�[y�u��A�X�-��hщ4ǻ��T]��fP3�_ϯѯ�Z:Ebɚ!���K�ªnm�m���������<���]`�u
:��nJ�IG`8��6b��(s���3�p�Ua;�P�9#�d6&�K��t�m�!�O�"a�)o�+w���Kt�#�!4}PV9>�G�2Oc��g�c}T"%���{�6��66'���T��^F���8m�d��6��[�.�,΀m�(1�I�,�湈������KJI���;��U#�}���c�IJ�s�����m\U)nrk�5Pf>�Zm��=ꝻEU��8��gN�0���4q�&�=$�X�p��c����d��_�*�\�Sy�o�d�#��x�}쵾W�-��<�,��\�0���G��H�P&u�Óo�ľm�5�B`#d@b�Q|���I��Rv�[ͯ�<�����t<��K�Bm4��Uxq����N���󟦷�P��N�������PT�e|M�y3�7�!�����D�����w�B��v3>�TՊ�x�z�zv���PM3���^Z���b`\����\xu��Y�]�j(x۸p��t�4�zX��)[BU1��C��):��hx9��������%,[>� �$�e�b��"��4R��$
���"�j��Q��6�������Sѻ�z��i���0y��8AˁU�&���L
�-���Š�պ��l��d���n�g���/�x��)NO�t.h��h��S����/�耞pl��ؒ%��a�g�B�0��X��+2& _���l4�*��:d韽��#xCZp��vyS��������zaTlj]|��h/���Jǥ/�F�=�3�N�^�������U��Ղ���a���VWKXwK�7 ֡�h��H*�o���V��o*B�4��F %U�� p�p�V�&�@�#�2�$� ���.��ύ	ݨĜ�~䋍;�$f�/�|�{��6�U������_Y��Ւ{[徙&Xj�2�T�twD�K�:&�-�_Q@�1S�lU<�x.�T
����jdYR�J�$XH@M��w��n�49���yo��%��h�9�S#��Op����������ĠD$L�3x	��J�)ۣ��c�ﻳjj�����c܇Z��L�pq}r6�I�tq��q�_���ÎCד�F��"�nK��:��"���*�����;�M����56�}��V$��:N�\l�f&���	��?�Vd��ʻh���w��fWٓZ��sIHM{~���@㢪;�����C��&_����()^eh�h%Zh�VCq)-[Y�c`��ۃ$e��r�Bg�g��ϙ�;�Sb3�2Cd����Zu�M��x�G�}�J�%���>6@x�C1���鱂Z� �ӏ}����h��:�S�̹B����'�Tl,�/��@0�˥��sXCq����(a��]䨒4{K��W�f�7�_��n�{�d4��җ_n%�g�]���
2��V���2�GU���`p�kc�Նf�
,jaD�3{��a�d�k��}��K,����ӯ#�����4�E*'1G	�U��}�l�S"��[�k�����EJ	b "��#�ʮRq� �2��Pž�չ���*�I�w�j�b���!�S&�����ݎ�3e�d[R��A��I(x0�]�h���do@@��� 2ܱ�ߘ��I�oɂlۜhc�zҐ���;�z]�U]�A.�%���ED��䑹I����cj�+f��K+_#|Ӓ �$���qV	v�+0Mv9�O?S�����RY����y�3[l����,���?X�x����e%�ۉ�:���%�E��.O����u�_�5�� /Y�ZY�%Y�ͼ�-ti��a^�)�qnQ$�z���o��YcY�Y����f߳l��z�3�6��<&�y�=Q��ڍķ\ڧ�B0͋/
c(�k6��<H����|���B%l�C���d��Ӕ8�z)bg�-�[%���'32u����~��M@��Isk?�1��� 4�mۡ�N�Ԕ�+�K,�w�j�M�Q)�
�(�F���̲,!����)�ޣ������"9]�üϣ������f��Dվ`z�`�72��{α��|i�zؙ�9�Y�ҺFS�>��j쵀L�oF!�,�$�T��\^D؀��_�������yU�'��;0�a�����C��-�`p|���3�/n��Kg�g���� G1��
 �Ai�� uC�0kX�Տ��#����Q$�_�4�M;F�f�]cl!Ua����^<���Ju1$��L܊2�#��ٚ�p�F�3�=�N#2�߿<�VU~\v����=a�������ha�z����#�n�4[_8wu�. Z�1=)�8�"�g�U���'P&����L�l�*��Ǝ�Vj�UVZKYj�qP�6z�S�=?�>�����G���;�^�}ʚ)��Ȭ��sy�B��v��ѽR����~� $z[�/�ɸ��,Z���!�ŕ �tK�����̣i��}�b6H���>k���?��m�8x�*Y�X��=D�Ϸ�,���^�d�4G���(�E��"jn��Y�g�S'�S.h��ϡ��,��T����X�����oK����;>Ӂ� �
��H-Z�s��p�{:R���O��@^�^{��d�L��)1�����Gƒ���%�^����m�;��UF�������Q$M�>gד��s��S8��v8E�fS	��t��6kQ(_%a=`�J/��JS��ܥӊ����\Y%�$�L)�`�]�3�i�49meLf߁ ���j���@`R�m?\���g�u+7��TU��!�ݼ/��VY�v^�.�yٮ|�B��%	��`H�U�]Ve�?N)@~���!籑"��G�.�ON|c�@�c1�G-��1��h���0MJu�h�:r���b�tn�z��q�zuf�'��W���Zܷ�Ű���k���Q�p����V�inqB�c��H�� v u�%,����>�N��`:ɑP��O9;��|!X�e�Y��h��C`#��� g�"U�)�Sɗ_l��E�_�5{k��d�T�~)@/�2!^�b��z!�� ��:�=4�}��9�b�p��A��a�n���O�_�5H�B����zL�9�K��m����Y*�O������ԇ
���ǎ F1�R��8��_�'�3e&�˝��+F��K�t�l�檏�U˚���-�� �ݓ�����Jw�,S���Ӕ)_pC��`��^>�ij�}r�å�vy���eI�5�R� �v�KK#���J��Py�ϥ�̸�b(�I/�UD����F8)��:Tj���8�g��45����mni�#(_i=Z��Ydr��~z9E&�Ta�O.���8��k*���8n~��Kj;�w���YTt5����6���J\az�>����d��~V�S׬,�o�I)��Z���W��=�O����W��1|k[�2���JQeY�HW�]D����	�E�&������R�&V�}���k�ו�&��_��4q����?j/�52�*
���M��p�r5빝�5J��>IjuD�&��&�G��G���m5��yE[���U��j50X�	�5H��<�҃0��4�v��pR
�n��^�����{s��W�L�/1-s�����pfs2�*\t/�PI�HMz=�ު( |�:<��s�b����u���
�H"��{�KH��`��T%�����R�N��_H�NRs���� ����h7�.dt=�5� ��Pr��?ށ:!8 �raLx��	^!�a:W7�_#�A�;��T���Z�v-�����hVG&m;Okj�|���܍F��3ٛ����n$���h�����/S�Z�f��Sy�S�o�#F�e�yN�<��l65�%��Wr����gk��6�zWwk嶈}��}��L���~A�� �_j�eZ���7t�Պڭ��Oȵ�Dy,)ު�0-J�������s3���A����%36���\��-�d���B��+?��x��E�+	���BBF�a٪�(�W�k)FQ��4�U=��Z*B6n}l>=���$8K�X����ȿ�Ss�B���
Z�Gƛd��n9������]� +]��m�XZ6:�$i�Q�sۅ�^���X�F�QnUW���6�)�0�/8��9
����|e6>ٜ���[(4y�S��˴) ��^�kR�N� w��[�u�ы���fN���+i���T)1�ZY����93/ϩ��=��2c7�9N�k��������VH��7��PZu]��֐�j�� �d	�*7�B�%��~'�X�%SMͺ�ygN���鱼,����/�Z�k��"��tĂM1ZA-�ڻ�`�2RD�%����b+��4 ԝ�G���p=�U`�c�L�B���0E��@k A�9��葬Ey��2�%m��Ig8|- K+�5�A����9w��Q�rW�8�eM6]�ʩh�h�^{�qw����?������2��wiMW�=�A��Tan�|�W+�IW�n`B��*����$z�k0<<n��P2���w���ǎ��LX��r8��e�7b�AN���������YrG��j�M\>}�	{�P0U�Sn�a+�c�����ſ@=A��u+���7�|�[���<{�ɢ>-@�9ŕ͉y1i����:��c�\{������W�n�اOϠ�A�:6!����u �>�`���F��S��K�n-�3������ �H �����U-��h0z�U�����G�i�ѝ@���3��'���E����HA�4��01f�2.�	�Q�7�q6����խ_����2|�L4!�5Jl��a᰹�xm��rf��z�K�k���%��^"sE2 �%�r���v��f��B�U�dv��0*!B��?Ӹ�Ѷ�=���#�ݙ"�4���ㅋW����Ry�,-F@\�Uf��C;pÞlyh��-��X ��*�Z�'��1=�%;�iT�ke'�?)�\�[���
g��(�Pk��D*���r�Gs$d��cK���ػ�b/��g�'�&N��RV��t���2e���>���Q���$Wm��kz�C�+���u�����k�Gv��Wd�ϱ!�id��j��k��Z�ݕ�����S*_X|E�H���P>�I��6��,(�DX���XƐ:��h	�^1¦|^#}/w�L�%$�6}_h����N���h9A��~��)ϐ�c���Z4��T%}2"���:������H��6�U���0�-���w5��)+�&��	3�a5G߹�!�M�U��~������!t��|��W����]�N�b̙U0C{�5��f���iE�C��`����`���[� ��9���S�[����RJK�u��w��㯪�{ c��\�LM�8<���*O��В�ES'I/���xc8mՁ�r���F���eh%L���=��>���N� :�L�J�)�zјO=�J�=#f��Z��xǾ��ZwL�K��P5���,:G4�J���1�����l~��U@iQ~[`�=/�y��~b�
��E���U��f��캄�^���p��O��/����&"]�.1�l�0�G}Pg�t��H��T���n��D���4�|���9�<?�'ډ洅p���_d����u57gut8��W$$����o_���t����)������ZX�]]Vp��aÑ9�a�)����_F,�v���`�����`�7�m
�#F��<C"�$$���8����{�@�u|��
��}r�$A��4�l��8HD'�&]��a��dV͡I��ߥbclg��|5�l��D#�b(m��2�S%������iJ���a�Q�K�˗���'���ǉ�x_�Q�2?8:�iz�&`�o�/Q�g%��	����x�b*-�t���5#uᲰ����E�Yqp��1x5�)��ەJ�v��<'�|��"LѢ����v��y�@ҥ8թ���c���;G�m`�|�gʶ.uhH*��E��uH��TΛ!���Ͷ=\0~+���׺���(7�>yІ|5��=a7����8��u��qz�%,;�ǸD�~�݈��`�$.��8� �F֎5�\���a)7A���@�0+g 
�c���ȫ;�������2ݶ*4*�]�ˇ�7�	!�[eɰ�/,A^�uYP�m2�UtӤ�F���8�e�Yb�,99�NNa`p"�z�x6�U�� ��0��O�ޱP��V�4(�Q��<�#,����Y��2+
?��3��	�@amgVW�V"�.����U<� �@���xHґu\
��Ry��R�%kv�k<b�? U�Gu`�N�{g�h��&�xw���O[Qխ"Xhl�6�N[�[���KGr�<��,�����&��x\L��`�m�J3.ށ��/��\0#�șa�*��D�����
-t��c��'�a��@S3]��%T�G/�G������r�E�v�"���
Cܾ����<�MH4vl��\b1��!�g��J �!Q��8F
�r"��o��\�s��~�rٗ&�i&�5;7ir�Tr!��hz[�G�ǞL���S�%��#�yS�_�>�xan��o5��>7���⡾y����C�����t�Q$�����NhE�]�f؉�������)K}�sr��?��;�k� E	��p�|j�7.�Ȑ��7U䟮��+�`P�k��Eй�Pڔ@:��ŕɞ�x7`]��1J�����ER�HƦ:�I��eX��bUb�,��s~��I#�6��K�O�����"9��X~Ө�0��lra�i�bΨ�׭$ ��]�ԧ��`T��~��~'�� X����v��F���y��`@ҿê5���͔B�$�E��-�����G����U�=�(;���p7 r3��ƪ#Y2c�gjy�Wx]��>-늧�0->��`�Uղ[2�\^��3]���,�S�,�݆�~��]�H�>f������`$E.°�7Dg�m�mv�Y]UV`
�۲�����B;�� T�����WsM��
d�8V5h�Q.]H�
�fI�+�[��d��ךQƤ�_�[%����#Rv����OQ�>�N���:̓�}[��ϙZ��h5������y�=�Ԭ�qvH�Bٚ#���mx��3�Nw���H ����a����D���O#�j3���t(n~V��P�y�
\"�eZ�=� �@GQ��_6\�Wa?̟��aPK:�Q4����U@�=u{a��'��i�7�����mV��i�(�V��IbT2��xZ�`������h��%.�%`���'z	N3���Qu�ژ�ie��*O�s�S�McMvK�*����5�/cz
�Z�����-��m�b��< K�qu�'b���������o��Hy�܄ko��[�Z$?I�q������m�Um��&B֘1�I?Ү?OXp��L���G�jG�0���+/f��9ZY ;��O��}'~���G2�/��d��ao%4bST�������~�k:<������v���R�J�Dr��-R�-4Uj=�>9; �6����j/Z���y�ڪV�5l�'t:~'��Tbr5D=�7kݯ|8X�E���'~�rǇ~�,�S�!XD����]�S��ƣ�9�cF<�5J~���@�f����t�kONui��R�7u	�V��H^�Bb�w2\Rn������
�A}������"g���΃����Q%S�3|!�}�"F؎r�>��?��t��:��'��A�R�[�����Z��
蓙cTMm�|��$���ӝV���F!漞�����E�OX����y3��!�*r����N�Sz�v�I��IrY����Z�����	���E|���UW.y1U>��L��Y��SU�TD����sʤ�Ɯ-�ƃ�㚘w����@r�*��[��!�<���<��Q
��K�Z���m�<5:�Fm#���ں7��rs�������b�����)�n����G�M�=�ˑ� ��0�@��Ϩ��Y�%�K���:�dB��l����[fؖ��qJ�&{mjY2���0�%_
g
���W�$Ji�VҎ�p���٘;��9��euI�Ɉ�ܚ��כ|H26(-��`E
X����sx�ZN���R@f��,�u�&�R����C��$z��d��P�1���l6d4�!�F�/��bd1	Y5���h����K�0|&?4������Y�m�N�Tg�:�s"�}��.?Ҭi��
 ã%J8Te*�z�1Ӻ^�%��#j/��fQT�m7�;�G�B(NGIz-|�:ІIH�Dz���J�o"�'P[t�'IQ�X.�p�A��I����� ��,�{9�6�P�z���!k	��Pm��!�:	j#�W:��M��+�3=/�+_��	gq��(�X��)�}�l�����.���oI���Ÿג���:��j�%.�)?��Y�_F�wNw�s$��(/�-+A�&v�1����8%c0R0�V�$O���"�3�@q���
���|b��mؙ��7��)�Z�cpzBd�T�(�u����W��e�FcJӬN���VMM��2��}P�j�绣�_��z�-0���0�)鞖�����!Ђ�e/&���n=���0G/O���o#�ŃaJzp; '��h��9G0ॾ���L�XU���u�L�Z��4D!7%]!kt�%��� ���Q鈳�����ziȪb��F� �ت����%���o��6�� h��V��>�z��LT�t��Oa~ұvM��#�W������&�1��M�k�!�ׂx�E�DU�]��4� �B��&����� ��ptW��/F�)�BwU&��$q�IqYmi��k)PS1s��T� 6�m�j>���<f�'z��iA�g5iu�b�;B��K.�cDs7����m����SgK&#@x����9)�h^'���������~��u]��n^��Z�}�p�����va�8�o0����ˮD<��o����#�1E!Y9��,ߊt/�������1�A�0[�$�̪=
Q�@/4��Ũp~!Ğq3O�-�	S�1ރ3f��%y�3{I�����{-ѧ�ߐd�ZH�m*\�)DpH�!���A�����Z�	\��A�?����[f��J���]_����Yvk��Hp%Yc7�( M�����r�@ut��s����e����[�,���Z�H,Z��X�X�%G�úo�I��qP�*0~'�Ó}�}C�;�ձ��|��}r�	4yXEh�}��7���g�{�ⳕv�3&S�B*#�
�w��N�)��DC��G���F��Z�{���r�z�Y����Fae*���psHH�.s�!p�L��[�'������mM�4�9�sӸ��	�wͧ��^6[�dX�
���X٬'��t�5��y:���(�2঳9�̿�����T��0�X��}�	[r�c�5���&Db�,�)tT	�i�3'����zdVrv��Tb��d-A0y�9j�Zi���Ppt�~��4��;���gu��s�i�: �"��y�D��3h3�䢒(Y�����h�u�X�Y��pk-��vL��쮰�W�99/�	�	���hIث��y��r�|(�����F���V#6g������a��Y� wP_w�(�i�nӜ�"l^��;���+铚8�J��}���޼$�J0�~�'���rS>�bF5b�E*kz���N'~�w`�$�C~�l��ו"��$���1�&���h~���r��k�ܣ	g�Ǳ�o��������?�!����ԓK�h�2έ6�d|-i��;r�L���wƳ��m���sn\!| �5$"_��b�n�;ǁ��+��se>uy���gP[��)F/\�C��?$LZ��̍6yۑǖ��`;�Far�!�w�J$�h�z�J$����r�}}B.S{�*�,ۥuU?k�_���N���0�O��A�	R�@"ڈ)fJm�m=n-��*@�C>ׅUj�T���:$.>P̃!���:��`G�YPXX'��'���z ���]�YDt��ʝ�C���6�/���v�I���@��7�Qh��HW�_%6�BK�Ʋ������#���#���m������L��?��ۇPSPm����)��w@����V��$��{�����Vdm�}d��b��T��B-s7�ہ`�4�1�����W��z �n�%���i��+i��xu/��v��ѕ\U���ݛy;�ߛ��G!�q�b��
�0�ے���j&�%���v@��C[��'
�=��TS��î��ww�7�u��H�s&�D��6��˯��UB��gSUrIx�E�\����g/gj:�'�n��j�S^$?
HB����S���貮�Y�1Gr�i��[n
(qh�1���̓�����>oFL�a���3h�ușI���y��_��8��!�[�u@��>�����A�h� ��š��wC�[=�dنRԓ�/�[�J��'?R�~�B�71�!��F�<�ƹł:|Zk���x�i����0��A��#M���đ�����[�_� �ಕ1�(���L�K%D����s"?�on��J�[}�<��jK�o?���G^ߏ�v���y�ᑢy�3m?�!U , ��U"GX�Ү�`sECK�M��(3��ͣD9('&q����N ������c�k���z��j�K5�*QG��9$����Z�*!� W��ٳ��"�G�U ��E`��7��Y�� �"��%�������|J���О&j�$+V5,��?n��6��4��T��>y	=�:�chFyH��m��t�������X��9x�����bJ����~�M�i�ړE�bj��5��ݫЃ~���(��>݈%W�u�ku� y{���B �5�� ���=���̃$P���F9ީ\�e�>|��!G��Z�����7��{U�gK]��¦* ,���Ȥ�e�T�OY�2��'�ݓ�;?��7(>�T�*!Ö��Ng꿶�p+�X��"�~���r�#ۭ� ����̤3 ����oI��<�"E���*�y�����:����>��m@p����5�m*��ʣP�şדC������B�z]���ۙ�����jK�T���`���_���zЧȤ��������|�!�J��bJLM�"G�V���y	ܕ���^.�H��r�)'*��y�g���jj��r������򔥔 ��� �o஽�Hm/�!B�R��.�/�=��0�ψ��s@1��t}���	�ư�2l^v*X�Ij���'"�����('�ݧ��@F���U�E^����+b��^]SM�zW�4P1Д"���}8h�D􇦔���Q͐gB��OW1�+�'[���,��7t=���M|�9�s�^s��Z"���TH��eW�Ew� MlΪ�W�Q����yk=�-C��
�V�0��r�0�>�Yv�<os��7�E�B�5���Yi,��Vo���7-��@)��_�[��AL��忖b 2e:���A�F;�%���|X2J�;vz+���W�Ѿ	S�!8��9ش���amb����!��� �TV�� T���X�y�T��O�s����Ҏ YV�Ob�lI����y����k����n���;��{'��Ɵ�����:/��8�?�w׹Q"z(�Nf������CJ����*.Ɍ�@~j��*��6���yv��Է��5}�?�(���v���7J'(�Z'�����@����`�oWѬ���eZ?**�Ƒ�V�����c�l�`b
��\\��!�q��ۋu���>(eu[rV�@��{D��&�X�ժ
��:+0j��1�ly��?�ꑜm'�o���*C�eC�����.��;��ֆ�<��,�l/-�
t��D����d=�D�ڝxsO�^�����U�o��+}F�=��ƊLn ;̧�����&zh��ԑ�C���h��a?㚸+b���lo���S�π܅Q�K�_��� _�2�7scXƅ+;�Pk+���S0�~���qw[��[�))Y�e$�K��0�b�B
�)a0���)�J�W�G)G+�;��M"z���X�j�ŀ�v:^R%4n�W{�V�Z�������6��M�^�T]QӗRH�����@اW�
�SK���߇	��$�ܹ�	�ے"v�<�o��߃bҗl̈́��%�I%�F<�:=��eX��ݲ]r���Y2'��En��tEZD�=���6U_Pf��L�w}@ʾ',�z�!�X��__�4�o$`��=̆�r��0r��v�K�]��C�]�1��eܯ���U�]~�E��a�=�D���w�U��,h���	��01�2��}���Y]2���^4�g�g<d�Qz��wg�5ٮW`�2*�����ǀ6��bt�-�&*8=�Y-a��Uc���T;�:h�������/����[���|�w�1]$8��,O�A���S�j�U5��>.���8��Y�(�z횙�{D%��+f�M�v9lJkM�T��?<~(�r#�x�mm���h�3s#�Womt�u3�@�-����7GyS�9-���>���d}����2zW�;����2a���Q�X���D��y>9����CfE�.B�i ��g�k#e�/�N�TE��*�*٨{�ߢ�>R�	���9!78X��=X�������.B'�t�]���< t�@�rd�.��s�u+�١���>�$��}��@�XLl�g�ݲ0�56l�9��B9Zu�	�bq�RȄ~�통T�%�_ѿ{.�B1�U<a���4���B0���WRf��**�P>�p&�G�G��T#m�0Ǔ]Z�P!���.p��{�@(N}�;�|"�@qil�^h�c�~WԒK��~w������ׇ'�9��2��w(��:``��m�ȾL���������</X���т�ˮ��;SN�/Q�����E�j�1��!�x��Чp��̧[�����ģL�@`�r��q�.�*xH�����!�^z>����[8����}
�l�6a�>�B�Ws�ϓ�W�w�7�)��
��<�@��G�.BW��h]Ŀ�V�Ŋ3��FHY��D�k�H�-L�F����ѯc_��kqb.O��H%&ʖ�d���Ƈ���N�(F�N���g���@�rI�?-���6���I���<C������ɋ�-�t,-q�87:�`ύ�{oG��|5r[�a�;y�d��I�?:��V	�f>P�8��?=4�c´<�z����V�}1���� �[�xeX��S,H�ypN60�]�O�	t��[.q�|��Ah�Pw����ج`�U�҈@+i(t�C����{��J �H8�x@�d�V��a���p�WgnU��u��6o�(4�>���~ʕNd�L?\��k�R��t��9�S`�H��\�g�^ o��"��$�*��;h_c��A�[O+��c_ D>������E��#����i�<d�p���F�J/;��Td�:�$=��P���g$(.�;~��	`����G�IX�\�ג�&w�N�~�KAX_k&8�N��Z��O|���,��Q�T
'N���Jc�IR�%r�c��R��1P�#��k�i��գ,E����`�{���}`�c�R~��(D��8n�i�6����N�|�Xl��d���y;�A�A�a��4��`��X�� �7~7*���E�c7�twc�S���@X�@�抰x��&�(��.���q�����F��c��\�ʝ"�O�y�)^f���*7��[H�9�~�=oۘ.r���Ǔ�bo�>�,\�~�o<��s��C�HA܆WKc��q�8�clGJR^enՈ���<��aP!�S���Y(�9�5���m��;ּ;��9&]'eD���Y|AY�ٻv�1�||&`��s�舒�?���W���-���
�zGe#2�Z+��ɈK�?��������ˡ����	3�x��vY�H��^�'�����B;�ͪس�O�>��+�Y����.�G���R;Н��P͠��)���Z��D_y�̿�`���S6h�ņ���E�T��t#.��z�K8X�i��,� �5c�B��[y���FTa���h0�l�>��c������yS@�;R�z2R�AS�犛����A��5+����6�����oW=~D�Z�ݔ7�H�_&bڴ
�tꤚ	���ϩ���ӂo�|�'�j>.�k�j�d��@kO��0�����vOǪ�td�dg�D�A9��N��V����dK^�?�.��]Rr ��%�>#��윰�n��H�94a��[�N����KE�>� Kr�>�̡������0|/�O��wd���@=����.����<.mj�j�\	�����[�:Um�����k�h�Ф+�J�������l�g���P���`�;`3���`.G�,�s�C���L�*�T�Oi[-"o����v�Bd�f>���F"�	�����F �oX����3��a�����v�=��o���1����K�#��{yd���;�P�ҽ�'7����?���"L�wpl�z���@�������aHaal���e#�L��W����ἐ@��I�/��S�-nY���@�`N9�Β
:#o��`J��<��[�觱�FzCcUwv,�����ˊԱ;$��(��� ������c7��5��Lr(���bz!}��VN��~�a@�4��QMGZ���k����&v�Z��%n�T�m�ĩ��H��*]���
�F��l��!��.	6V]�Q��o4q��D�֕���a�r�� �� ��ws�n��EF���E~�{u4C�L�_���~8*����j�'9 s&��8F\���ϗ��^�R��djU�Ep��	L��l�[�f�/�BzT�d݂��; ,�T��@Tb�G���a�S>��H�ez*_�uྟ�J�����T�dAN���jE��87�+N�8վe$��K7�A��,6�$�v(d�zֈ<��J�qg[�8��h�3$��pP6 ����Ȑ���SVCt�B����q�n[��g_�y�C�z���	�U?��<8dw�����o��
)�"�uG���?&g��ˀ�ӧ�kh�Sx��[j�;ň�,��v�� PI�L�Od����bmŀ�1�=�6�^Eͮ���L���n�;` 	ݕ�L�}����?l��$�d<���M��D�S��}*�t-���L��K��Ƴ�	�33������d'�5�d�S�k�A�̨j���������k���Y�|t��6#U���Ad��f����6I�?L��f�т��y�G��� ��i��ΰ��^�,Wi��q�C���t��@,���L�}	�v��k������@����h��k�߽P�jL%����`���x�Z�
	����I44$����z�Aze��P5ַ��{	���M�?�.���>d����!��\#�o��N##)�u��1r��n?��H~x\�q'�� A�@�P7V��V\R[�@����nm�l����6�>��K��a`��W�8��5a�{��e�Zrs��N��_7��'��bR����"�8���� {�@ĳ�	��ݝ�{�Dn7{����;ȅ��	�S��+4ҽ�+�1[-�$ՈO������%Zud�k���h�E���/�ZE�~��V���0^��N����YJ�얜'*/���/��;�J%�pU�����9��bY���BR9װ&4]�@�Jˠ����������12!��;C��XN��A�h��O.v��1}i�z��yј4��`	I1���Wi����)>�zt���A���p�K%�����͚_���2}K]r�P���\֋�>�����@����٧�|��`��������'���)�UZ���$���/ZqҒ.pb�>.�>�'�ҁ礛w�E�%�-�6D=:CV�!Vե���D���Ą�T��oI�Yh[�:�����|/$>���%�<����D۪��~c}εX���	����U	IB��K���%�g�Iە��N~���p��C��I���E�Lk����7+,�eۧx0�D��̞p�iYp���Q�S觝r?��T�m1)35\��H?�*��ڴ���>4��ܰ�c�R�f����iS=h�'�c5&;9��#N��G���|��X$�pw)�2g�)3Pë�rI ;�����8c�G3��ĳ8`1j�st04���BS0�	J�lg�O%�F4O����w�&M �o@]�`P�P+�O�L%���FE�	��\���?|W�7&3pNǷ���R7�F�Q�/�� g�"�鑧�eiz��,�c�x��&���0�jT�⪮��z���GRƎ�7�H��w2����}�p�P��r�)��%Z�3��v(���FO�j���-a�(�/�M�fv��ـ��`f@	��d_��~͍�3� ��!85XO)��u_6�׍���
�{�;kB�Ԯy�٭!D�����-I*���e۵�Đ��s�F3�K-C�CFtk�zG�����!e1�6=�u�j�׋GSpg��wd6)5�@\���  �r�����˨������e!f���+�Jq�[�{������F~��Ip�0�H���}����[�w���Q$�����՛����O��=Sj��s|VYQ~�D,��k�`��?훷���UCr㬳�(=a?�� t/�;�'"f��u�`��;���eܠH�-���lͺ���P|1�m��N�R�w1�e��t��]q۶Egg�-�}$'�[�~�L�l<��q�M�Ke]X��Zxx��D�{��݇0N��
lu�J��D�(I2F��p��5�jF��S[�	�\?��~,�,������㷅�k���ŗd�;W��aB#3�꓇}��f�ݪ�fT��� 	ʋyb�E����3w�T�6�@��&2>�Q��$� A`������gWr�crY*����ص�eȇ�_�h�M:K_�������e)�R�H.�Pd����ȉ?���"f �s�P�:Գ�.�+1_SK�F�"��s�����c:dǦL�¯����"
(�_�/=�t�M"
��܎����>TI"�4�H�$ф׀"C�?�R �sy�6rq1�^�5�Y�����u��R�=ƉC�
�V{��	��_��u�}ú�Y7�O�`x�۷ma���	[F��b|0������n�q����֗�;�ӡ:~+�q�P��6k���=6��`W��D�Ʀ������"J�\�w	���7�����m-Tvq63ٍ)�
P߻c�[÷W�d�&�����n~`�Gq��?M���u�q��2{���J��]��/�ֶ*e�U��7b�F����S��Y�Kd�z=q'�K�Ft<\����i#%�6L�ܾ�� ����f�-AI��8]E��a�l�+Gt��ǝ�9��(c�p��I���F�F���0��r6`�	_���-�0�l�goOvbvׯTj�c@����wBB�ޤ�β<V!����7�e��ʟV�qGf�P���,:Zf��:3�뉁�j��?�atT"נ�7��`=ե��H5k��vt��2標�j_�4H�*���RQ�T> ��u\<ft(�M�jh���Ͱúr�lj�.��X�L71�߯j���0�h��x}}V/ޙ���"����T��,]bxS�|�g��SH�r~�I9��;6��l�?e��z(L�⒒��k�����ݛG �{0�KM�%V��$!JL��ʠy�q�4�����"Wv�����;��^�6��z����
��z�L�x.O����D����>Lj�%wp�
�Lߠ��0ɿ#]O�YN���P���s�A����8"Rl*G��w;��z(�޶hC�s���e���t�J�Oؗ�pH�ݫA�\�|�۷t�h0�Q�{O�pW��G�W�b��G�ES��d��/�G�6qS��p��ٌټ��{�#m�(���@*�$���}7�7�J�Z�EZ����ƞ6�?�u��4)�l�fȚ(��?\��U���by��ο�&#˞��j�_��Q�)�ȇ��7� ��#�k�%��Wμ����nD(�T�����������4�1v݉�GՙeB��i����=�P��"!>E����W3�!-Z}{#���C��&�U���wV6��2�xOޤwsh��\q�������{�|��'<f~v���U`4���I�ݼ_�Z�T�~�����O?OvT��2WH��Z�*�D�攃u�@V^c���H��sp��K3�O:S!xzi��d�g怂��_>��u��$�.���,�L�y	�X礼���8��4&�@K�MG}<>�Z-�^�����_+b������eS��7�6��0{�Vb1~V:�}�&I{&�������քO ��=D٦���h���yJ�=�tw���Y�PiM�L�Իk��7T���k���̭�)�?�T��^OG��_�EU�z�&�'?"^�^*�r��σ��xc)yL��xT)���)9�8�YwG|d@
�uX[i���R��i�<7�G���ֱZP�43�����2��y��q����Ơ�|��T����z�9S�
q��	~%Z6�2I��ڱ;�~���xD���� ����l�}k�{}׀��r�^�V����'��B櫽���R�(&͞��汴8G��`S�p����r��A�WA��x8�ݟ/�{��{�d�k�� �|K~��s�NM3ӕ�pW�*��ؾz��-�(�H��^b�{���+�oi�h1��kD��3Ş޷�L��l��/En{�̳5TL�k$U������6�Ԩ��6���n[ԩCm"k�͚.e�CR�u��<��;��I]��p���ߌ|-L׭�8��
�z%��5{��,�V<pf�v�ᮍ�k0C��C5En>[P���� �!@5������"��_�����/6v{!��Q;P�|dv�������:YXв%kJ?����o8�º>&�~jH���Tr�VL/�i��dAĬ�?�F�M�Ȝ"���L&j��5E��W�����b�q2��B�J�Ƈ�?d�n< �^�1�V�*��e޸%B�ltl�SJh11J;�P5�򚡩r*�-�G�"��)�e�ę��Xɳ�\ɹ����jc�Y�)5.ӓ]0�Ϲ>�(O^��.-~�Q���h�SJq�5�
��[d�'O��u��d��z��I�S�2N;T0O�EE����c��(}���6-j��GK-�T����7+{TJ��O�a)��9�p���w�~�7Z:�|j������iVQD�_zQ�1=��22^���E���}�e�ɇt��@�ϰ�T "��5���Yt��6�4
�SBy��v�K'퓾B�i?!�&�a���3����38"��e���΅N<��������#ז��x��=,��<Dv�{v�J�Hl*a0	��68��qUR� 6')�*��T�v{j��Iu�}�+��o^��er��C��D:6R�]GG0���:8,hxD������ݨ��ԺA�W�7:����*q�P�R+�dpRS�R6H��3��|/���{����������5��� &�՘�p��9�~������� $r<�Q��F"٫�UȮU]�N����Ba
C<��ؕ��up�.H~����鳹��t��k�`ԥ��!�� �W����X+N���r����\�xW��n�ZNWT�e��X>:��-�rW��U�#�����`���.Jo�%�y�ۖ4���U�Z��wk+A�>kZ��q�	2p^
�_���V�L��]�f����,��J�V���r�[�z���.�໥���3� D���2tDn�|{��Q��|������H-�Q����'��gN��5�Cm�fZɽ�����+�V$��E:l�pY�Ӳ��OM���/��D�݌��{8��%�7H�/��[m��wN�Ag~w����#����E|�^r��*�d:���X4��w�B�]�K.C3�=������4��҅I�U;Bl{��L�G����C|g�p1s6��`Ēx�����OQj�];Z�� s:�S a�O@J�ʷx_����,r����� �x �Z��ߧ��&Ρ&t�*�H�Q�%�?2�ޚx�fY��i�ʸ���`��_��:���\7M�'	@��V�X�C�D
�F}�k��9�S��Yb��e��L�z�X��+��&I��vP&��B�X�E��Ğ��P~�oX��Ǵ�(�/�)o�u\Mp������i%33*�W���nn���Ezf��������u��ԁ6�	@� &�n�]5��I8��q��t�"C6oۣ}j��!����1��W��%�Lr�'(��젃�Q�pvtPd��m�<��t�V!���\��o�T�R1B�_��۹g�;����(WhC1�lh�b�IX"�����?	Q�Y�1p�S*)����K��#��8h���gN����� ���	B�@x�A�D��h����MEܓ~MN|N��F}땔�c�1*���Z���7��,Ks�Q���lH��1��a�s��;�(��N������u^���_�V�����C��l;p.m�}��n%h��qu���81�/?��
�Oz�g����A�@i��L)T����:��7P\
�RO��U�!d�@�h�?a�=L��d����A�s
�zcE��:Mz͸��s�"�Dql�
���=��,O�l��b>��k�.rY�M�C�1U�)���W�9�ħ�+�\#7�=�b9�G6�%FG_��f[�{���ώ�\�?#֧L��ݳ�T�۳����t���� Btb4ԑS���څ�}C=斏hf}����}�+ϪW9���������N'��U�����3ӫOJ)A^�EW�U�A�p'��wb
?b{�7�,o5j�pJ�� "dL>��t\ބ�[��T �q-��|ڌ�|��kC\��(S���MR��¼��iZ�hrd�	�3������S����^���k�[�X˛ٮ�s�j%�{C�D�;=E��R`\b	eS�5bS�����J��FB����p���.7���M]� 29�A�̾W��
Ǻ-�5l�WQ�!��&�q��3���V��CՆC�D��o#�>��kZ����.�h�~=Z�5��	��k��}��ĥi����Uu�UӨO�
h����~0뾩�Hv�Y�i~^�9N#�؅�)d8ol���6�\,hl��ɥ!#�kipo��g�Qʷ����p.GS�&�h��:�#)S���㨕�W98�7���5��i�4=��75O�;����(�K9�z�k���m{=*���?���S���"��+i'�'|�'�o����|m��pJKn�'���:S@֕��_T��X?�����Xl�p���Q��.��4b0}�O��o���`�nh�\KX9�8D������{/@6��''w�Jog��n0�څ{.5�g�{���-0���ġ�^��0�R����<���Q�U��_ƌҲ%���	|g�b��I^�6G"(�!�r�YR�4��(o2�j��˃���jƽ�-���-��db��?�|���񆰩_V�]������T#���֎ZA�#f�� �%���CR*��ڛ��7U����F�S�M�q��B�H�#Lm' pnH����v�x�l���C3&;�H>�lYPMe�,d�Q�p�G�q�`m�(��^j �i۰/MH7:��#D�|�)�׽4����mC�z �\�*�܏iy³�)�M�������l(��ߞ�)��h&/���Gt�؃@_��xLՇT������[���r4O����9Y��	gE��d����+�VPva^�귋	��JF��د��l�f�:������**�tɜ��FEg(F	�X������!�nŃu����� [.�5�j8멐Q�)r��� �L.-�|���0�̱�X@w38�����I���p	Aa�)������00�h#�6�^S�^NHMft�ڠ�d�����Ypǽ>�o��U����"��9��s!����s״1���ϼe
Of��:�6ĵ��c�]�����1�.]��m�uU����ci�4 �����H��t�o&A�}8L��7�V�D#��8_BQ��e*M��=���� �;	�?ϯD�����f�┾]�	�V�NdFW6� ���-�)$�̮�ϥ$�e�~��M�S�]��,�]����:��OvH�<�m���M�G[|7�*�OP���n�#���ִa׍�M�����~��'/��c������^���\�j	�a����/��U@�4~�'l�kvw��r�^�^y;�B9�*�(w����UP��G/$���|��H�T�7~"
ߺ �*���'൐0�ؼ����q�]�'q�=K��\����ߵ�W�9�6�,]@���ܼ�M��o�B6��X�a���~J�O�}G���SL��(�
���k�0�ς����{E*����&���b������ll�Z�"�;7 ��ӈ1��k4l��~�/GZ�K��Is�u������۠_~��p����c'�����������sP����~V�|ٔ1]��:�z�[Pƾ (�zɅˇ���U�É�L�)�I��:�k�$�Z�X�|ql��%^u���锹O��dԣ_���?�99�Nm�q���ѐ�����B���+!��Ed�[�`�h���sSl*�꽄m�?��s����R�t�U�u̙�Ɛ�?fh�<�����>�
��7�mj�s���t�����C4�Ȩ`���<��<XzŖ��s�Q����ue[^&W�����.�_߰6�� `��!��V��?b�H6��'�b�_BA�;���E��z �Ŝ���C1q�6���@� 7��>����c4��A]�A�x�
������mC&;|w�u>̻�6i��jE;�7��%�ˋ7'������_#��ε_�21�Uz���q��h����2W���	��Э�"52U�r�#�oZ�g����[G튽YAZl��`PJՊ��@NdUQ`�c%�������a��D�$1�.�|�y����̯��7^�P"i�F���.`��%Mg�ݓ�Eڈ�U��ꙠB2�e��Xc�9���}Zt��Mg��F/�s�h��?�m*�����.~������Y�rv���0(o���aN3!�B͙�՟E�j�5İ���v���|��TSB��{�Yϋ�-�UAo;a���bqW08N�����J���5EM�rj�:.$�|wm�	M��f��[�:��=�i�&�����Ka3��C�r��܀�£֖u��HV����j5��ӕum_6}P�5��尲ڠ�����(��Mrd�x�R���{䷓CՈ�&�0���歓�t�I�&�8�3���SD����.)�:'	���&�OV���m&^�f�mbm#���p����u��HD8�d���g�Z�"A��:4 7:��un�c�_	ڔ8Q6��0��,����&8�Kd���k�,��R\����J������E��x|���������XBdF��2�ek�=p��C�5��L�皿E:�J��^�����n��0t$��+^���G}���Y���k�!75.Ԅ_t`������^���	���i�=�ȈѠ;��Eؿ�<�[;�wl���H"��E����O2	Y���Ǚ&�a�(;Tj}�h#=!��g�V/\fS��?ر�]��
LU�z�����9�@pl�;�;xy�Kw���t/��wr�o������k�A��L�>U�f,Ptt+��c 7F��}Q1��M���K�lѐU}�Ðd��6�:�N��)��Ղ�r���>�jU���+2�����b�Jl� �vlV�Xv�ԱF���꓇1�'I���u�7��W�g�0�܃�m\�6�e�L:+`+k{2Z&�|&�&#n�r������k-��@��7�L�Z��8[(���kb}��d�R�C�t�Xw�t�	��k4����@�>���������S��T���5DW�x��6��^4���ȷ����}c�y4��7C[��=i��x��ئ<jQj6����x3�:e��uA�|��\I����a1J��7� �'��QA�\Ə��ªYC����������WW���'�R5�)"m`�g7�L�Z��� ���뷺$�� >׃�Ĕ��,�/ 1�0UA��b<��p��p �ȇ�DJC�����(�SZT�ʘ����=�Q��+A
B���|�1��P!��|�?�҅��r�'�B������x3_y���/�#Q�$�ۈ�L_S����AMn��;&��X�������kF꒢�/��M߿Q2~�7�*�N h��͟���*�5?�,d�G��fIͪ��:G�%'��'��%ܰ�fo�@��u����Y<�'3��x�X.�-J�z�i��0y�u'W��p�k��>�~�����Is7���/}���X:���#Qg|�h�q�?;��4�ky6���M�FwPq��Ec�E ����l��hJ$���f�&n ,�k���6^�Г��<w�]c��:�=M�*Ǉ$:2th̿�1�����Zm?��6l��#����#}[��|�n�n�S�F�΍�����l�&�	h���]��Z2��Gqky	����|:��cKZ�^�&�3�M#o2{n��A�n3��e/�+Ug���ȹ������v3a�}���¾y�t�9�w? ��%��(�5P�<��I��l���
��Ǡ�v��4��NDڰ�yȟX�rlq�릤U0l�-�o�C�p���b��8�/��T_�'�"�N#�7�oP����6 <l�h��,�Q�'�a+����YG�\x�߳9>�C�����J	�9
e��
����M8�!�n��M�*P�>��Me��3��uZ�%|ՖR�oԜܼ�4�$�/mN��P��������A&΋c�hi4@²Jp��m��x2��ϰ���'���c
�ɷ�1C��Z$�ћ}�Po���Ev�C���?G�In��3���Sr]w�נ+��D�]�Ӥ����2���r���8�"�����R�|ęؤw�B(۷�CwT� �3����V�c�[cҌ�ə�Ma~�=�|<��2���u{ğ�k�P���d �9� ��ɱ㔐I6�uD�1G!7!�U=	��C��<9��T��%	�KU��$��Ǚ-��N���`� rR��.<JX&���}�YG�}Xw���]f���ԣ���H���mNI~��ͭט甒�ѩ�!� ��fK󖊲P|.ʚ/v��V�9@����d��l�Ạ
M�y��qZ�C���������3�!eh&�?,�
��Q���K�ʷ�Q�*1�TvN�����|Z�]g4=�<\]�
R@�B;���Y�s|Q����s%����΀��Y��]����};��wk\y�n�4�/���I���%�yh�x�
/�.P�F�FH���zCč���-�������AtL-=��)�tB�I㴪A�ƽx���=�rJ����'���ŀ��0C{�+u�A�I�H}Ǳ�Ԁ�,O%��E���Y�(����z�S$������
}�Gv��7T
���빈�Ž��2Ү���,'��=@�;��<�
x�������{ϴ�]B�s����|���ֱN��c��\��I4w���6�#o>���M,�_!*l8S� {v�=��fv�_���?�X�×h�0o�	ȯ�8:n��8ɚ�0������,�N�4GdM~J#�]��y��C���5D��I�x��JA	 �ɺ�r6=��@/Hο�������$#k)���ۛ�O'��D,ņ����oI6 ����M�'��@)#�ك��z���w��3�	B�ki>tN��T{u���Ӿ��Dr�$��ӥ���I��QG#�݂E����ަ9��w=T��Ƣ�E�V(�F����fI����'0���3��bz��@�\� �����n2�6x1L��MnZ�O%.�B�=��^u���y��I��3��[�P�4<��M�wֆ��v�E�F�R��Y�ń���?
{��2fxEWg����В��ir���:P:P#��G� �ir����S��c(W>��O>|�1�8>z�2�u�-r�_�㯫�"=�����b: ��G��f"�t�qf���xwI��Py�ex�T��zl��u!�7qEfV��،�y����}�N��*�qyM,p���k%e^쨲���f�-�&v	�VN9P������AY!	�������naVG��!D�ǫ@���Y�0g�b�Vo�/�[��5�C	p�'��@���euK���k�J��t5��#t&A2�FB������|CpE���0C��^8>����ĺG>Eh>��72$N�c��HD�p�ɔgb��`���iTpvs���i^��8�� �iQ�M+8_aZl�������J�~BO��~�A\��>e^�bb�U�1���=���9� ɷ}�0�U~�0�Hp��"#��׿<��o*�=�f���I�y&�ҁ����+�����KI�Y��8����1.�-�>��:�Q=�r�T������>��o<�zU���5dH�}������T>`,r��3�.L��*��"H9+Q(z7�r:�K��lܵ���;X2��*2�:d�Ɓ䩷~r��c�m�g��^�����1��-8S��YxS��݊daU�Fό�(����J��y]�V<>$	�H�';@��v�{�-"�< 冓p>�y<�6�r�܁�h���r�f��D����4���Ғ֡Cz
}@BκR�|n9��Y�-��W�@Irv�S�u1��>~q������0������vIrg�&0ud��G������Ǧ���!@~k"��	�8����0[D�J�PK�[�j�E������-�I�K:m��@�HH�U���&LrԎ�3�E���s�0��&�K�m餃��pU��qXӂt��T#��E ��q�Y@���ޔq�%��3ǈYek�3M��@%�T-�0���q�W�0�W�(���(�>�MD��~6�����5�Xͼ�����`���J���=�)`��#Pf�:����|�!a�_ΪWW�[HT��nQ���*�%	�"v;d7��]$�ܩ��]Q-�<���[r��N�X:���n�-���b�"��S�~���,N�7���9L�>n�CEO���du}ޱ /�~��7����w���W2M]�s4�)X�9H���/��`�va��\
i�'WfJW�>M���
��5l@Xԁ�J��.���ܞ)���8��{w>�����T�ET=��P2k-�y�BB��������N*�  M9�546[}�
ߚ[���o՜�3&�}�>�X����ö��GK�g���7h��e�x�=wwq]���f:�Ӱ��
������9�HAdu�o�	N6�
{h��WX'��#E	�j =�`�BsV���<p��՟��
�7�����!��^R�"QkG�P���J��>��MlM�}D5�T�%g&���Y���%���)5��JjZ�r���(_�H`�ښ��z��HkV]껥2o& �R�|QW��?��gi�F�S���mx�vO���������A�[��J�:=���4�qX��+���ƃ��<�{k7ⱍ[E�K��\V�BX��E��P�>N�inF�Z}�VۛZ)���Å�3��zD�|B�NX0N����ͣ�l�T��67�2M��D)(D�{x�+P)ɤfU�c�9�i1hn� \2Q#��y�L��R��d�nbB*�*�d���ф^8�%W�D��*�Igy1*M�@
�+I׈��_�_���ڶ}��Tv���� �OUf���)02J�����N�XT"���S�ޓF~�j�:�lCL�w���#D"�1j���l������g��F,Z5���shM��,��: ���,����A(9\����o}����P����8�Y��c���� iU3��2d����C27�::���������`Y[ѷ_w#��tI��KQ3~��Z�.L)��C�Vg��{;ی����o��V�d�`���B֐ ܫv,�Y<�x��]'�GF��>ogq�!��T�M��Z��m{V7��^%Tq�l6�@E4�do�v)`�B�HY�X�9��xy	OT�+*ґ�!�9�o��n5,����\r��,��.J#�ф�Y����{\��N6�NQ��?
�_��b'S˨[=G[E
͉x1��ž:���g29����:��ә67 uB�9Ba�=և�Ćf�P����{AL�=��AQm2��H�w@d�AӘ�Y����F�[���`l�d�ǉq�G�p���d�sPR���Չ���ҥ\c�F����Ϲ���P�1�i"{���c����74,�	�S�]����V����fXh�|�(.dR,���[P��L3��l[�#h{S$��Ű�E��M�4��g1��_N�� ��š��nt�����zKAM�x:ݶ=Ϻ/�?x��X�f3��ю�k9q�2l������ŲX=�k��|h�4�����$q�����ꭃMҳ�ܢ��h����qKN\�4Y�	�9͋.��;�>��:��dP	4&|\��QR>��s�z���	��CkK;⦑0%#Ij{���-����!�*�zݳs.���3�'ah^��FA��W�9㾩qE�Y�W�-����a�Ka����Ž16�v��!��I�)�m��NPu#QuL.^o�i׀��z��V?�r#J�6r�c�*t��{��X�T�ʬ���∜w�Twx�B�Q��dmW�5ɝ]yW��Yr!�p��r�b��A�Z���ծ�j�ht�Jպ,&����3��́'��S�M7�H��6`��G���p�b͆� ��ܗ�G,�0`w�u�F�_��h�1�"�"՝&y�J���
����>.�O��k"5��q���v��"כ�Rȇ�拌ÇdV���&�)[����1nPVӹ�i)g���f�2V) }.,1������t�U�	Q�!S΄C��=X�(�N?��=**`1ōb�8R��%rW�O���H�w�@�8��w"S�z��f`�:�a����������y�wpv��i�����T)�L�5������sn�@f��/� ���g�������~D�(#���׾��o��#�.х�����k2�8k��E��cퟭ\�܃�#���Ɯ*��cC�X�g�� [�|6G*�9?�/�h]'V �����}�uh����ŝk�"KX��(��jmo霜|;�rBV'����^m�[�b����9��+Aa6�>�����b���eNH��\�N�.#�TB�@�D�	,f���+������>������A�a���!E����r
��M�{�[e9��h^Sԓ�	G�4�.�3-V�C����ieE��"��m��_ܤOi�ԯ��tѶɭPcA��)�88�:uЅ�t��%x�]�U;�Q���Qմ�8�0��=�2'M+n�����������aA�8��jP]����,bR��#ޑ'\�xTN�z�G�	(������P�p�i��i���[n��J���F�ڇ�P%#�ˎ/7��7Y����H%��rh�w�6[C�*��Ry|aմ��b�Ӿa����ˤ���l��V����q$��q���~NH:F�C�����}uӜ�Մ:p�òa=&�"P�x	��S��wiP��:H��C*����v�d�?��h2�)��/B���Y�䵧f��j_w�Ɏ�	�ɓp_]0C�(����Eک���X���D}�����6\�R>5�4�4M1sW�ߖ-��
)Lm��=-��l�����-�B�Wz_��NJ�[����i�|��(�� 4�
��ɱ%n`��0��U�� <Ϫ�m��,�S����p	���Nx�G����&+J\�]�2��%��L�&pG,����8��[su���rO1���"`�Y+��%G��V'AW�G:ig#����tʋ�jUy�}9*���?��F*�MaT%'L�1��p�f?}#�$�t+rՎy܌��8�2����f.��-r�\C��"�>��I��IqL�o�I�ϔ�j*÷a�� �k�$0�҈by�B�5�t�l*��/�c�z������Ivh�x��۩��`^�ɂ��8fj�q��ǋ�1�����XL�D�������A���L��R���ebKVZ������W�	���=��Q�7_���(�風�H�@�u�/�V�(u m��������=����u��
gi�$X��`�s���^��F��|�!�h����5�&T���6�^RP�uL����*��^:�!sF���?���e�c/��l��8ȷ��@lI��w��7���rٷڔ�g���8��~ڟ�qe�-1�(��=�xzk���8�b]��<��޽� 7�x��������n�He�(	'��R���J�kO�a�O�6r_����j�?���Z��]��	b�gr����w�r_�˶���؅��Oh:.LvO�z�[W���ǝj"�m��9����fR'�<U��bC�҉��F�:�u�Kq9{���{Q��4W��������)�?�Pf�9s�[禑�MQꊬxo���W\�@�y�x xf��@�k#~��7��vJ�@���`85�nF]gF'-����>E�ǙB�9�U׫l�0��" �3����@��mR��{46�����u��j![��<n^d���.[|y��W{��Y�"�`S����JA�M[��;Yk���蟶�:�! ���z�G�a�H¤B�4=]'ȿύ]7dF/h�A���R֫h���؈�ԓ����o�U�J��0o?ry_��Ң?�6��Q��r�}��i�m,D|'	�6��9֔z������k6ȹS�y�f] dh�q�X�Ntao]=�y�N����>���8��<�iM�);���)����ha@��g�z�ʬ��g���$�kq��q��&Ȉ�m��S1ˀ��=������~Κ�������z����{6&�	v�R�W�(h��fǃش�,n���H[��cx��apI�L�����0".s�^^��mE�X��e~��s�u����md�Em+V1��5Z6�0�Z]�� -�j����ǳ{��u��vV��+�f�X?��J1�@�·r��҇����]����5�c���Xs����jh�g��e�q�;��T;(U��o�~ͪ]ɧ?�3��D8�)�h��g����Ш `��o4����Y�>�t�Q9	�^e��� �OdI�"�2����m��(%Jc���t��Pn��_���m�y^�i��.g����[�CX���l�� u	�0{�@�Ó���td�q[cܝQibGR���u_�R���*���u{��>'�f,�d����h�8"��7;:�[L߼090s��SR�>�t���|Qp�^�U/e���l��(���"_���ʾ��O�k?mt����������42�q���Z_er:�,׭��7F����B]vٿ�͠BTw�l��/�	G��D��0O�o�EPj}g���_;��*{�8'�}��S�Br�6^�4���E�2圅w�w������H��I߲  Ό�;n�D\�,#�b�(Ϣ�H��̟`g[/wI��C(Su�kو����kS\�qt7ٻ?h���Z�Ń�D>�T6K�=@�A����'��pS_I�<���ưʰ��1|���Bt0��ԝ���#&�N&�j�W�$�Gj����hWKS��]�}$��A�j��i����^B�Ǒs�r{���6eT��c�NLz��Ь"���׮r.��\����̋�];Pq)��]�Wed�/~�V�=z.`˪j?��.U��M��/��3��!�PL)Ŝ#!�A<�*/���ّ͞dZ:�¼���x,�A\W���H����/�)���+�R�N�n<ہ���8�Цp��DI�5Q ��+�K"�-�E�ޙ�k�ds]���
O�3s*�b��Ǖܖf�H�yn�by�ED�F��p�<Ɓ��Qf�c�8�ō؎ҩ@�ɝ��(�%$���߫����Pu��V�W &d2G��:�J�sp�Z[�:�R�爉���΋���-�r��A���_�[���j���礇 }�O|ߴl��Y�d���OD�K�=3������%I��p�e;�/ߧ%�!$&�x�M�߂r�����*�O�zr�������Y����@I�'|ȼ�/����^�(h����elw��1\���X� "��U���7�BFy�K��-��W�����^��)L�Srf� R��f��[��ޗ �o���c�dի�'֖����S'�1+�->h��ξ��ޮs2|��e��D�$z��ޓ-}y:Ėq�]�Eo��]��Ws0-"�3�h���� qmC�D���P�>��e�\L$槕�pC�OA�]s�\3o�p�h fZm��$aE�z��Ԗs����+����ϒ�ljl�ǵFd�\X%2 )�纼?�i@
і#�UI��g�P�~a�v:����QU?��I�������*m'd1�9������!Q%�ew�yb����{.'؋���;�ֽ#2J��t��ƨm���c��Q�2i��@a�\�e��-9>a]�貶�8.ٻ��TK�)	�"۾�G����3uyy2��T��5�?1��W!E�Y�aҫ�8��'@�/i����ȏ�����\����k��4��<+_<���E��d7��u�y��Z����n�G:}�gI���pU̑� P�Z�x�f,X>�#��2j?bp3f�Ѿ-���t��3�Wx��*��0�ʑhS��<YI�Hܰz��jg�"=��|��J��i�<�3~�/ǲ��K�b��d/��|��g;uwA���)\{��@�8�|�0�~��-��z�d��$Q�+�im-��n+NeWĘ���M�R��	��ڂ~��Ŕ����0 K_�۰�`��?̘\CU	u��āMf6�~��N|A/�x���xϙ�2(]�쓛5�7�mE�K�E��-�(@l��M�������<��ӞXz��n�&�4�g�)��e�V���}{�h���)���z@4٤�hx8�@i��OvC�T�/�]�q��(�(!��~��~cLsGY�8��-��Z:H��E��"?�	pٵ�˸�o<��7"g�.Ny�H�r��g�7�)D�����:���T�_�G�Yy�V�ʞG=m+� ���덖���_�����Ҟ �XR(�^���1)�s�$������%�6��8u�
U��/���N3�[��;r�Y �pŀ����P!l����0;j�:��se�����NI����Sj�Y�;7�{�m\�9#����{��%i�=��26 9�MY���Q�ŨI�5~T*�)�9�c��S�©oل��(���fr��g�6�4'�<5I\��_�#���K�){�Y��$H�Ӏ��7�c��Q�O׽"����� ��t� 7=���?�����:��#�Elttj�f��k�^�ه�HӁL��W&�5���K�{<�P��
A܌k����5K�`��ߛR��Q
�X�����C�6uX�4�\���J:�9��3�LD�N��^UB�S���u�M��g)Lu^:�	��Ҽ_�HC��|�ʡ�aqG��KY_Ʒ�,a������)�H��`B��w�$�w6������G�Bx9x�]�#٠�X �4LN�[�	�N"n,��k��³����)r_?��eu���Vc�_�1�i���q ���.���gf�jݥF6��KM�����{#��ۘ�	��N],y�S߮́�H��Em����'οM��+���H��>a~���v2��&��U��6&�5�N~B3)�]L:�ŭ�5>�kX#����֞�Ȃb�w��	�	sg֖/���<\Z�/�iڡv�	^�Y��ܫ���� �K��ʋ�q�*N�r|F��2��Bq���a��/�Hrkk�f�D��X�;�^Y,
>�nka�OD/���L��S��l�m��抩,�I٨V��ʫ�5K���,E1"��A��e4�݌t�tc�������f��������"��Fv=|o���R�����c3w/���_��f��1�e�N >I@���+�P@�aMg���'ЌX�M���\:��[�Y�2��J��y��Q.�iJ	!�_���8E��ħ�e���4���V}(p3QY�>v����sM��xyȲ�PȪ���B7�uj����L��f�P�G6��А禌A���t���C�٨s����+@K���v\sW�(��f� �f��d{�|��h[���\�3-�Cp�Ԍ���������'��y;�����֎�B|߉zN6�4$��oH�H��t�֊�)�_���q��LDBy�4���6�]1��"ɶ��I5M'�:��^Y%.��	8q9 )�"}ݤ��&�X5_#D>��E?�f��	ku�%QV���I�6�� �ɥ
e�ݕ���ku��	��M�Ϭ�N����1A���]nR,��e�B�@�>.�$�e�����Le�x��JF{�l�Js�H%g��h7�G�$Gሲա�o�@8�Ay��ѽ�/���XA���oĴ ��G�x�N���4�"��*$�p����x������}��C�����͕G��X��w.�?���t�,J,"=�m�]�3��NQ�"`oMhw�0���S��b'���5ڨyy ���0ډu[c�|r�FfC�vC�n�2�92Tu&!���~�{�B�_�����f�8|�����	�;q{�c�����l�`J�G�_��.��^#Nz�+9���I��������9��~c�H�B,�.mh/���#U8;�&�@'�{�����UX�(��l�	��Un�9�+6Q���E�&%?P�ogm��^p��'�����?�48�t�	�W݈�=Ch^�pɦ	�5;�R�k ��`��w��K�������ɺ�!�%Rk$S� ��.���:�� �I�̈́�h��5���������d*�E�y����f����/��~���d�H�_�xQ%��_�5��=T	?�\��w���a��-zx�=$U�sJV�qb��g,�5(!��x��119^M��ڸ�>�	�^���J�窍�,����������0-&z{YH$������r?�`��P���'L�:+��e��� J{��"�P�y=��u[Ͼ��*��y9I�y�V��,]I3�8Zކ_�s�BYh��VI�n�Xq�)��G#0�UWYf����?����.��Q�PἊ��'��	�dy舟�c�\[�խ�AE>y���=��5%�P�7��c`e��������u�ɿܼ��0�s~���IM�04T�]|/I{��� �R�-������a|z�K���V<j�S&��2�E����J�G#���Xj`�R���2<>�jj�C�y��J�3����_ď��2�7bPF,(( �볆��u��' �i���q�J��)�D���0肟Y���Z��XFh��|kX���a�f����l���3���U*��i�AT���#�ӂ]���]�_%��p��A��a� j��R@�x�i�	2؀]�o��1��{ڹ�9�j"�U�IݛK)P���ق~cp�Ɔ9W��?&l&���t&��6�3�#��������&�6��KDXCD҃���]=&(7@1Z����Z����L�:��ʶ+:"̩��j%��p�@s�D�щv��&��jH���������l^�R���3@�%�`���0�^y́A"7@�û�v{S{���x��Ϥ��7Xg�|X�8���C��
��T�k�g/GZ�D?ѿ���{c�-ad5�)�wX�rJ=�3�/����.q�)���E�\g�Ry0�i��BI�b���t���S���?iۘk�1k�Db��bl��f��!N7z��#2�~�G;?4��>������.��=)���N�Zi��3�[�e{��Erl��W��S�a��+�z',�RL�u<1���g��/b���m������j9���e>Eo�l��FA�-���d�(�+�~�b♹A�Q�i�{�KJ�|4brU���Hְ<�@�*|X�m}��ܑ�*��>DO��[u(T�jC�:�����*�TR��U�k��߷�W�.��AS��D7�>38��}H�K�3ޑ̱Rk�
ʠ��^ZV����K��WH��My�#tr_3�͎��>k��h�6�$��Y3��%dٲ�_zÎM43o���rQ���A�hsZ�l��3t
���r�g�F��=3����1g�^�G&+�>.��u�(���`�~8ɣq�:R �׫ύ� �BT"�A9�M��uF��(0'�f�M2�+Ā���p9]i4M��'�'U��h�q�;��ܨ���ݸ��F��QBց2���Jn_��wf2��~u}K\e��ǈiG6'�?k-wsu��Xx�Ǳ>�	b$l"������7��ԣ^%ӣm�P�Zk�" _$�k��l)$�ߠ�L�wz��EW��,N�%��p��z��=1d��<~نӼqfL�[ڻe ��@�_X�H��I�u�ǍGW��y�	���~�\KN�]���tUH�s�!dOu���uμ��"��:�a�����m�fC�����̤�aH ��#'�Qؾ�)�)<���pXT#��̨�L'�ki������M��N_�s�� >
�$�6vpe;�"si�Vn�y.�$+�oQk���ȟ��^Գ���M��OC�UA���f����t'����E3�k��4�h'�og�.�&*$�.�N*�~���d}��T6y�y�����%`.�Z�xV�&6Q_��АK�����Zo�����b5�^V�����X�ܦ��:��hD�����_	`;
w:�*nۂ���Ȼ
�`$��/,U��w1����s��Q[^������,ʰ��Hynj�r�pg�8窓W~ H`��kK^��d��I���`�.�Ҏ�ܦ���N^�v�&c����-H\���[?��v�t(�0d�
�Re�̀�[0�9���AG+Հ���'Ar��?E@��h^�8i/�5�g)���V4�&����' �v /�,���LG�BL��g0}PZA���רmW+4���@�"+N�Ia��j�R�c
'l���?NE5ߞ����������P����0׺�Pd��/Q����uC���W#�گ>��pjd� \�#~��Ɔ8���لo�H�G����0��VnB�J���P���5�	����Kū.�e]��3����0����:��4��[�a�]����-k�l�k��{Ƿ����;��	�`Z����9KQ�w�> ������y���x[@���v��D�ӞuFf��ŗ�P2<���^�!��U���m"�Sb��c��J$�����+�/��I�!g�ԏX�����t��T����P���4��i�0�P?rh�����dS����/��%}���sBvL*e�bv'�x%(u�0������vj�-Z�Q�/�0�K3�h��G)�c�X������� SZ��?�u�6Z����`���V��`�����2�<d���p(�����J$6-�4�WV5:�d3�\&�� P�0OH A�2����!����w��� �/x�����\���L|�%��hd�OmKɧ�Ĥ2ON�
0'�W~��}S׶ª�'�X5�f��#�����X��	c&kV���L_u r�c�p&�~�f����9-��o7�"$�,��h�����M��Ǚ&�2�M�}	���A�ڏ��t�Ŕ$�}�&1�-�Õ(Y���;�ƻ��B��e�C�B�G�� ��4������H7�Ƅ�LY���H���1�K�W�*d������0����ƌ��V�|�����q5V���ٓ�aS*e�����b�,�I:NBgf�~���K�Ɨ�Y�}۴�aR��M�ч�`��u0 ���Q<��_	JC�pVE44���)#�4�BsF�����Z�82�TDl���U w�"KbQ~����8Ҹ�����4�;[U@�^XO�����p��o��l ě�g [������o�W����ޜ ��������@:ё���<����� ����Jx���A@�,�M�����V����>TI$����e49T��(��w��ʬ>��N�ŵ�1��Uq����-G[\����&�p�u�g�9�YT���S���z:�����v���Śz&�����Hr�f�>�O#��+APݟ���T��	 ��?r�l��К�5O�a�>���n��
-��b���b�&�w���6�%V<�� l�I�#	@0��'��]���r�ذ.�y�P��C�]�$�� ���#	6���4Ҫ2���[z7ڟ,t��B/?�	��c���.�Nɋ�r"#��ɧ�,/�#�+7��?��P��Y>�q��P�\�2o�̧
 ���#��94f�X��J�G/ޛVu"o�S�/0y&NF��#�݅�ՈN�����ş@%�><@1�/	M�*th�������w�{Ԭ6&�7�;�j��@)��@�hD�4��Dsb��];�+N#��J`�jPݖ���f5/4���2���3�`t�,?��	i�QZ5M$_U�����>��ˣh��fi@B�D�� 6��vr0�w6�OKs�c{�/aރ;QrvWvf�f�ࠇGL�dy'� :~^얺�J.c��2�n���q6�����0����McG1 l�Vn[)��8�Q�&��,f�g���^�ZR��n���5=���i�[S����c��Д`MHAΉn�`�6���gOnOm�0�~��\������[3є���1Z�)�+ax6�ѳ���G%�1�l���w�PS���|�3���V�@Cή�w�"Z�ā��Uja���ҧ6�U�t ��n����k���U���ο!^6>��8A#��{6-|@C�^4�[����	$��aGd��(A�@�W@Վk:���U���^*�2�0�8cy  O�nH%����r������&&��m��3��"�	�_o W.ܥ_��E�/�v�D	��42�C�-CTlJ�2l��L2r#�FQ�H��ǲ�ކw�K{ &��pێ2�Ӵ{�U^4��.����Xs'<��EN4*�8�TSk{��>�
����gz�����b�l�?���q�|�<���mh�F�̧Iwb�j��vgA	.i��z���k��I�&��t�%�3ȝ�������!f�`nT�2W����y!�]��<g4�.zqP�H뉄�4{��(�A��m��%���x댄>�8=_���V�P�L��+H�ZW ��ku��ǡ���������ƯT"L�4��n��L���g;?#`��M�"��)�ho�"ö�aH���)�^�AS���f�7VVG��0M������HE�� �OG�eoLf8�\H���]��Ӌ0�k�&�=,&<m�+�T�gt=:�6��m���c��Y�w��>�q�WQ��nçͮ�t7b�ϸ�M��Q�󌯦WXx"2�7�H�"�XT|�K࿨�-)��@h��P _��b�wa�X_����@�KsDв~IY� xr���q �Ѡ�t�Q�\r�j;��^`(��(^�&�[f����-�/��	�vM+�N���b?���V�фڴ�O!�����w1\$�q|AY)�nl��}<�}%#�<� ա-��eZ��H`�J�C��g'C��;YR��\�J�y��r� =ME���i416�&�*|.�aP���c�V��[�Y��A�8��iJM�𲹸�d�g��L��{���x�m����CL{�F��sǄ���P1�-��4��4��1�O�^1���<��'00!V$�b����OE&f�0/-g7*+�����+�8�����()i�_p1�o[��E�{=Z�Kdv�gWDwC�0L-�ޘA��L�O9�2A��ǎy/ m��[�2���9�wbIvXa��U���s)QyѹJ�K壹u�^�#��$��I���8���}2���&`[=�T؄F�Y?�cq��M��b�9�H�]�@��G�j���H��LdV��MR5�YC~D#���`;��j9TX���`)0}��dQ�]���˶͸6�!��5����ײձgU�/�n��Q�ج�6ӯ��Q�,��ԑ?�|�mS^`E��hTqs/��ِ�I9�c*���oN�����(����j��������Dg?A���4ki��z����j��D{���i�vR|:� ~2Ec��qo�k�W�>N�)�u�2k�jUi2��v�zџt*�� ]s!1�ŉ~g�b�խ���.��u����&�9,o&�U$�c�篭�]ܪ@�hQz��6���-B���N�8�k���P�z� �g$SX�$M"?`��eT$�r�q��3h�"bRE�d�^�?����:( 9�c�ƚ��z�"��m� ��Ȳ��m�BhU ����s�t��~!�%�ҷ�=���qkHt����my8�-��:�N�( ij�3\�ꋶ��k~u�����%dcWi�u�W����>��|��S������య�=��{��kZɪɩ]~�G�#!��J�f��#�F�S�*h8j�G�Q�]د���$ٴ�W;�eyN<GwV��u�K�)��ϥ��Nz�2���+VQ�fa`R�z�����g��+�6�$��ve;1U���X�,�VoJU��xF�L���0�y��_tw�u8�A�_*�?�@q�_���r9o����+.�@��]�'�����0#�u�`J�G���1�r;u޵lhұ_�H���?5㔜�g�y�4��t>���=B����y�H��t��v�颉��{u�L� Lݳ�V1��艓�����\ډX֩�o��r^��J�" Skע�,GX{����2�N��k-l��Òugh�Q�y��~��3���rdh>\�룼���fY�My�g�(�U#��Y��3��`z�>wM �Q׹�P��Xқ�h������Y�rѣ�[G[!RJ�^?�c���z{3]s_� ����}�O�����(e��\6ι��ɿ\)]�]d�f[��(�j��LO=L��h7��n�t��7ғ��:����]�~��d)�`K��!/,�%�臷�v^E^��"a�$�ju���f}̓11��p!���K�"Q��Q1"��З����Q"^��vN|�Z�F��zh�=AbBX-F���;���קd<�p0��`�궔=�0�_�ť�-���!�/TA0mқlӬ>kq';t����M�M�ǥ��)�z��S����H\5���ɤέ�T�ť��j鱢S}� �>��h�VF<��.�s׌?���/M�X���{&ɐ:.ǂ}!R3'��*5�X��/y�Ц4K����@�&Do3WC�O���<�5L�'	��`�#Q!�w�:��R|�&�حҼl���p��`��X��!+��sX�`�����՞l��l���&��I��i�)V�WNqE�����<��h%��C���\����_��-��zF,��="��H��C��2�^ql���n�b������D��)�/1���
�f�wm�*&<��Z�G�����M��YOB�,<^�{�.�f�Ts&,q w5�S�; ��EO�y�y�N���2<E��cE7�YwC�=�=A>A���W��:"���{�]ө�KnB��Z��V�zah-��HG�"Ԧ6�ǥ���vk�n�xe9$
�J|�9�eʂ;�x���`Ɨ�<�T_l�<�g6K��F:^�&�'��`g����,���:�ì�0�� jg�����9j�����*y5��?,ڔ�"���m����0j�w6G}�$t����徙��2�7��)N��L�$��upU��pd��Y��/m8xi*� �} '��Z�cGA�Yq�f���i��[�^� =�%��-��*�̖��H��Y�j˰21[)s�1�h�iIꝅ������mZϴj�������e˂�����!����L�2a�^�	�,�|��t�~� ���9�2�"�\aR�� f��盽_�8�P�1#��KOGi��t�X�`j�[�|ϿM�f�M�V.��k���r���uQ�7��k}ъC���8��g3��[��B�x	�sI��`s]f�B�`�ˑ%c�O`�g��ڦ� ��x�|�	ܔ:���ᴴ�
8�ǊI�Ok��~ǭ7E�^�܇W$��_��)��6I�"ӧ��p5@�]�u�}M�����S��zIo��^�I�dK'��i�B� �T9T�����g�o�*���D��^W�4�T��uGB��5�P'� ��D1z
��F�bEGP+��d����d������A�֮�;�M��	m����Fw &�:d�v��u��1>����IR���Q&�.�{;�a�P�q��<󻛷39�)7Kkur'��'#N��{��8�5��5r[xг�vF�C�U��>�zlt r�P���?�:��F���@�K�Rbd�#TN�Cͩ��;��p��;��5=j���E;މ�$�[1($���!�G|p�Y�&{pd�_�A���4q�`���I4�4f����L�������- v�ރJ�����������_d�x,D�2+܎�Z����D�ڬ ���%�7n�甎$�qw����+�mF���v| F�i`2ka���X���	E�1� ���l�,aOb�K�J|G�=��j�=8&�����S�l}҉�rH�U��~�/ndᶣ�6�X�QC�R�U������.�����j�iaG+�A�M��4&���4r���B�W�kW�r�S�j�j!�k`!?L_~d0�U�b��NKK8ڥ�6]\��������8��Qd��G�&BC���@�1�C�+�G@o�E�	���P:򭄘��12/����Ƀ�/T���<���^n�:�Z)�*Y\�ѳm�5�S�}��kCr�Oڸ��2�te�ޞ�;=HD�K��+�1c�$v� }Z濌�����>R�!�����D�E�UU*4��|\� )�u��ҿz
�^^��!H�����~��Y,(��c��$�[l�ƺ�?<����ޣ���㏀������G L���5Z�&RVU���u��]V���Y�q7(,!�����|@N0��~'���Ż�];�Xno�%�с����g�ꇇ8ePGY���{Up���(�����c4�7���o��T��V� l��P�IMw�4��US��p�V��9_?es\�\����c�ْ���m2�@�:����f,��ǣ��s��.G�]�)�I�X��5��H
�;ai	�`,*%�/��V��^��>}v���� ��p�ۡW��PN�(��U`6Ƅ��Ʀ3h��T?XF��l�7b��<��(:Q����&��>��:[�'�D=\-��o�$/@�\�.�m�E]w)�#g,�Ī` >%��(��zp�5����[U_�{��rC�_$d�~�ѱs�.D1�R�2�Ϝڧ��	f�J��fp0s�2Q	.�KLF� ��D�n��7��T����L��캻a����+�m�Z`�n�Z,���ܛS�Cݡ-c�.Æ�2L
�Z�m{6��5�\�3E�e)I���A	:ZQa'{7�rC"�b@`���k̵��ت�їz����p�`�ӌ��T�^�9�@w|KM���J%W<�4�a+���#�V���j"%VU�ߜԭ�̺O�lK�wK��{9�{A�OkF�j���<��⺸jh97Ea��=�ϙ��Mƙ���_�S�#������W[�؁�]!«=��7Mv|t����a�zlG�O/{������z|Cl@�3'��	�>��f�QN��t��+�_���erk��jWj_ �$�xi��p�Z��q/��	nཱ�*$�&���N̫�d��06�`�g���s[��:��_[�tٻ�C�;y~����i�3�[[a������]y	�`�}�vc�Ey���2�Y��L���x�1$ؕ����b
m�M����_<z����m;9��P<ҝ]���T���z�u��M`|8^!N�Ղ�Y��Q���QP5c'�����P7v	h��b@����t��9�Ɖ��"?I�NN;M�(<*���)�&��A�=~��((ޜh����I�MAotW�kV���E���d�m?>(�3����\vW�|��'1py�4]�HY�
N�ײ�(��W�ߒ3�98�\;+u_�h숁��(j�	��h�E3����)lr&�O7W>�|�ׂ# ��J��K���,W� �����5B�YZ�����*My峫k����b�=X$2!o�0����F^�ْҐRH�<d3a�,ߨ���=s�o�Ώ9�N~K냑dp* L�@�h����V#A�wj"7<W,���$5�#��;�e�;�"��gw�ʦ�� �oz�+j$���1�Ԝ�r�(�pQ�,��O�����R�!�h��q��W���4��kP��U7^1�FH��y����/̹:\�K�C�U�mI�؇jaӃB����mk]�U��ʓ�ch��mQ�}5�"��|-��X4��1i2<,DQ��!Ӻ�^�� �Lv��7�~M��Fd'���T�Ki�l��7�J�	q�0x�� �/$��ۛp����R��M�x��MlQ�X���a|�ͼ[�*v�2sSi�ٓ;���g���	"��ň�s�2i�����3ۀ�˽�"���qa��此���K�lX�ވ�Q�	��(8�KJ����=C	��G�~/ɚ��dԏ��V��'�K�;B��˨�.���لD�
�py�5u�P�*ˏ�$�z�oN�4�~�<��J�=V]���CW�3S����1h�iZ��IW}cY,�XԶ�J����s>���|�D�:�5{޼
(�p���*b尙�|(�]d${Cʖ1>�}@��s��q`Xh�e�9N��q�ᒿ���ś���d��q1�V�����R;$��s��<ՖC����|�<Y��l^���(�����E��1tP<Y�a[=`F���6�������C>1�5	��7X(։oD�D��0�p���(��ͬ������� ;3׵��؄>U�`�������E�Kc斔Y�!�d�v4�埀@�J�q��J�f&r�3y�n=0O�F�bX�����_�sש6$��'��*��P����oso�<�����"Wz��/Y���̿/��H C���_��&Xұ"ؘ�4Ę�<��Vl=ۤ��a\X�=|�Ipj�D��r��G��To��U"�C�m��W���r�S��h �hz�Z2�C[z.@}�"
h)����I7H#�s�uy�"v`ĥ1lN��1�� ]�r�4chZ��Mo1��<i�	����K	�^b���3��F���Z�cB�����R��8a�㓄�i�-�Q�Ag�(%����O��w�]�����E��:1'S����k��ۆ��8Y���(ފ��c��Ŧ3��8�����uI.z�Y+�F�Ch|oդ��B�b�N�ŕ���*s

�j�%Ғ��#�{G��8�(@�}���k(���NG�Gm5���r��%C�
Z��i	5�c�T��}$r��5o��U�RY�� x��<\�-.dh����?QA��4�+f��~B��5�L�ޢ rI�Ψ]�ĜFɼ��{��4{(z�Y�!긷���?�ՉU����7�a����3B��P�\vH:^�&��f�3<��Fm��,����f��F���P�2]��(F
��"K��j\��ǲ,�,639���~kU��X'ۂoD�N�m��>�I���?���E4�z ���86�;Ÿ���F�E$s�N�+��'W����/l1�3Ǜk�m5`�:�ϐ5b�qV9骎��Z`��6��+�<_�*1� mt����%�8��~���*��*K����V�yaF���1NՕUABxq���"��;Bw��]���1�Z8,�d}e}vK�BY$�G������)ON�  j�0�:���1��]V��f�<N�9��Yh@��O����>��`$rm��zt+Q��+�%N0���@m����4m��	4}+��ȷ(�b�#��"��3^u/�Sh�ݯ�X#���jK��I� M�(l,у-ܹ�ID0C�c_qJS��� <k��)��s)dB��G��=7w��_x �� �L�	OW® Kf��g��׸��S%wHIb�Y�>f[�y������à�	�W��₍Ǯ��6*�Z���3�������j��uEp��c���=��\��Ϊ �7%�(��F���OV�J��oΌx���u,ް9[Oh�	�"S�&�:+r�󐱍F�!��O��i�lc>�9��I%�d�\���4��}k��l�3#R��h���]z/��t-��}���9�\�q����R�u�ϵ5݅�IGh���M��f��Q0�f��4!��[� �:}�e�b�������'W��^:��lL�?%����:��4��qJZ���(
�8D8���.|����d)t���s���lC���~u��7���9#�@��ѭ̈́��r��;�瘗�q���'�H��I,>	A�4�L�s�\��U�?�`hҸ�� �Qk϶}_5�Y*݇�*����F�Y�p�Z�3rЫU�1��|����/�r.�S�R�Δѩ�����^��V)�	�9ŝ��j��b���^K����=���%
��~���Ⱦ�N�vCjT�[������������¦g@GpG���;8��V%�.��b�T�S��*�L�.��xt��qv��p�ĤU�Y�q��=�P�3G�-����.�Sp��;�#���p�ipm���G0-�3� ��*��y��"�Nӻ��;&�(���:����h=�Ɍ0�E�8�G��K��MC��r�cUh����tf��=���+��v��̚ێ��^@��=�]�����w:���e�����`WL��|�#K(�n{D~M�W@*c�<�u�bQX<��gp4�ߛ�R���%�������`Đ̦����#��4���,g �!�]�ꮛq�f�E�!����Q���kJ�A�GI�<��J�V�6H"<�ڵܹP7��� ij�V��8����\b"����0s4eǢ�}��z��p6�O���8���Q�,m�J���_8�ᡔD�#�j����B�&��_C�1��d��K�D��[�m�hi!�&6L�o�S��t pY�w��;��%�8��%yj�o2�6'�W���`���v�B�{4=�'Y����"`���#��BE�n ��U�����=�8����U���G������U1�'����ɵ��4{R��g����.�>B^��L߁ /4y�e<wL䏝E@V��� 
!�����>c	�SNKK4?�-q޶c�n��u�Zy.�V�1�7��>T�I�S��U(�xz2�_�hiP�eն���Qe�3Z^��T��/��o��Sl�Ea]1<�aͪ�v�5��ع�U�	8%ŋR��1X͌�E�G�{7S��fg��*��!B�疟1���&�B���N��������>l�㭑�?_�D	(6����:�cs�ߒ��{�n}\'$1'��4��X\����6Q����	����=��c����B{q�$�ФIߒ�G/��8]��n3hY}M=e�v>0�+�EϚ�Gg�o�+>���O?4*~ǣ�S�~�o�w ]`gƺ1�)��2�,ZT8��o�r�8O�ԝD����Ѕ�/���*
4i뽿�H��?R�9G�w� -�ž^a�i����5=R�u�w� ���ٿ�.�B��.�����Mɴ|Y�Z�lK0��E	-P�1�B?ܶ�uD�S���+�όxIa�^��Ȼ2��6�+�K�U�ѴJ���Y������ZN\��^�{8
W��{F)�
Z�e7$o�������,�r�	M������v!`�'@�'�v�L�*�im��)Oݩ���-�s�چ	��
��d�-�^R�!���L)����5���eڋ����[��3.oQn���iBC!.�cH��,DغI�1:7��@ȍ1i`��fw��֒�eV��O�u�vA����l%9��|�����!��xN�����w�̈́��N
�I,%\����:)�><U�2�-eq��|���|�]��⵾��Fc�Q�q5g�@�h�^>;+8wKCUJ��5��G_��=V}EXV��g �,F2s��n
�aXA�f"��wJ��Sw��8���Z���v��V�N�ڑT%���P������	%�.^E��{�A$���ϑ"�GW�>l~0�fB���ﵒ+��V�2�Ż�5�	<���a��S��g��Sx�F���x�a�p�({��'[E��u����BH��qÈ��Cr8�ŷ�[��~H�S��tOl���!��~���W6ޠh�$DB7X.�Y>��1�%�E��.f&��df�	�Ӷj�
�e;-��:ᆑ�x=���3:�@o=2k����$�
�4���xy��r����҃U�x�~�pl�!L�_��dd`��a���{�V+�o�8�Ι~Ý-q�?�b&�Ftn��Ӵ?�B^#�5!�����s�͇������7EO�'��S\���*�m] �B�����D߉��a��4��M��˯\���2��pD��M�l
ͱY`B3�����.�"�wOC@��=��M=~��l�Q���X-��$h�k�	"!,�5�v��Ϯ2v�l�,ӨP��j����a0uo�C���'�d����5�JMG��{0�'%���a\����,\�0�G�TVZ���)���G۳9��(��a��*���j*�&�o���;�u���I�q�yF�n]�@Z�fA��!�f��2N�!Tёڙ\�"���[j��/��_����q7ܔ���9OVσz�(�Ъ �C�����5-o%��s.V��r(�W �.�:��%'�������&�%ld{H&�-�o(AzDc�"����Yn�`Uo�j����~���aYP� ���)������g�^Б���uo� �g��`��Pg���ucV*�� TZh���}��f�� �,�P���T���Z�g����L��S� C�aD���)wЕ�?���"N�ZƢ���ak4.�v>u�-�0�-��50)U&cz,7��y�K�2�5y��T$a�?ø��;����|���)~�G�C}OzO��J+v���fF;��xէЋrv�t2T^��p1T�`k��.�@9�"2�d����bF�+PT}Q=�h��o2
�k���6<E��FD��L�/���E�{
��eb'e�L;�6����wh�$��(HF��}z��n=���(�{��Ʒ����K_�hV)r�ؽW�lR<3�uS-��^'�)�a|�Ռ<:�-��.W��o�s�I}��[�Օ���s-�W����̋!�/Bn���?e_�-���镣���@�&滰�c��5��t����H����q�
���$���76�~�Sy�Au�m5���]���ҁ?����m�;����"0��9�xS����Έ�x-%�hz9�4&k��X(��;�&��Z�͉�-����=�����B�v5-z�W�"�^[���LB�684��2^�}?�P���I�2�5�Q߀�;s!�Sh��o�6���'X��nt�:M�/�<�լɳ��_x	�o���&C��S��ϋ�5���D�^h�1G�<�n��[a���zu�������j�;� I�s��~�S�!8{Y��9ظ��;^��5��M���D��@U�$�H�([���u����'��1�S��s�J>�Z*eTʜ�/�g�,,5p*���NC�0�9��*n�� ���讦�����Ӹ�T����{$�fX���X~�f�{ݖ,�BHo� >/'���1��i��\�cC/e���Qc7�3�q�U��.׶��(�r�0,p�SB��E0�`ҦAP����|�,��_�pK��[�,��5���N�v15��ʬ O,��C\ߐ���DW����Ϲ�+u�����gmҫh���[/.VaY�
�ڕ1��^-o�$JAg�򃴦 �QVm�Tī���	��㶿޼���r� �l���de���_q�u�P�����;���x|1�����ZJ���Ք�,3E19���\$����*"�0�	Ej5����f@-���gr>��	/ N=�3�G;�j�_%��һ6�c�]���3�F5�+�o'��*���0�xY>��.�B�"�2�¨�!��@�4+��ST]���Z>wury���5v�_sF��\�uWy`�ڃ����|P�,���i(���靲�m	A�e"�u����$��:'�5/�\)��dP<U��_��,=V3��e��Y8U/:�y�c����P��ހٽ:Zh˭$������V̿�Z
�{��� �G%�Ea��B�"�s@��{�����F_�n=�uZ�o�L}���.����l[�����/�xF��\�J���hC��D;���-�Q�P9���*�^�S�۠�1[Gu6X8��Q�M��=6��g�E�ͻwڀZ�c��K�B,�E%���]�NoG����ocv��fw�U#�6�kO��ꆤ�j��$5���1�ᆙ�*�m'Z3xΕ�'�����y�aT�1�X
�ǒwW�Èe�ZI�8��i��W�:�a=+��7y��*�S���giov��lw	Xy�!p�=�h�zIrZ�I��y�v\'k�d=(�bU�m� $���p�Y�8���ő)eH��8)�VS�ƛk�E���p�:���*�w�!��.���ߓ,ꛩr�sėہ�{{p
�nѩF�}uJ��{�]Ҿkѣ2(fr�E�?��j��T
��[�3"�-�g����{��?#_<���G~�x���Mlh�ED�7��ػg�	m;'�&]��y.hfN=N=X&���)_H�E'��WM���L�y���1bZ��r7Ҳ1�,�#���{t���ԏ3��NX�sA�:�~p���w�����L�D:�Y�t ;$���-k��ԓ�U�u���HUâ���2��*��`�hiK�%^��{CQ.�=�ƙη7�',<�MfM��+�Z�����"v$�~�UKO��#�``�T���&Qb��t�f8��!�Ě�F֐���T�X�ۭ���ё#)�=�� \"�JQ�iN��(�ԏ���#ZU�]�/�����]����U�����Q�����|3l���H��E6n�]�*��e�%0u3|�H�v�.��%���Z=��O�o�ԫ P������o�Lx�}��Y9�%wQ�1����Ш�u��أ�+ȱi#DՕY����Ғ����V9�N�v�^<]X�wO� ��b���F����9�\u jd^���m�öF�>�J��ږ?� �Z{�1 ��Ɉ�w߆��#�Z��BR�7�C��7��h����c�2ܻ� "��Q�D��#3�(�j�qp�_���5<.��/�g_V&�p���P���]����}$������w(�ل�s��Y@!��Y(��t�j�.�E�\�8S��V����|���	�q���TΜ�+A|n{��a�L{8q�dAq�3�ǭW�?��9��(��R�37l�C��\"+wp9��������f��cz]ě�J�o���ս3�a{�o�|�]"e6���!�i'_*/�:���Ǩ=B��(����a���	ہ� W%���!��{y�9`����.�c��1�N��!��ڭ�O���{��c�ʹ��dr�c�k���p�'�w*�5Eȶk4~�_��_�-:��ƚ�=d�49��Sۆ���*{$A�wæs���3?E��@ye��V�my�~�����8#��t���iR�Y������殯�)�(��R}haR���=p�O��|���>�1 u���~@������������D9�N%���f���B��¨�yG�v�%�Z,���G�(N��׭v�Gͷu|���7r輀+��f�HWg&���̓/D�T7��b��S=������Qd���IL`S��}�^I+�6L5��
�������𫖏dɎ�d ��m-N�����T}���c�d�?�H�G����Љ)j g�������>��~��(a���6DDI�;� ���;���<h�>�!6듅�����嬥����nHDº	V�w��x��\?ɛ�!��|�t>��^�'�H���$��ݎ?�H���ńD��_iy��AvQܘ��*�����K��,*�^pu�r����Ƃ�k�����cGIļ"�Ι:k����[/�Q�e	N�AM�"uL�A�&Kfm���wԌ*�S��Gy�>r�G��v�Kۗ�0
՛-T1Ys�49d�R&����H��LI�َ���͵�굶I��U���q������5[������vh���jDQ��I�W+��Б�Ra)�[, ��6vs
N��?��2T�'p�~��C�[��T�Ӕ$eL~�f(J����/���r+U׬4�t~}��-`��pY}@_���4m�PJ߃ƅH��ii���`�A=��Ol���aɓ�b�7���:��A����{7��~�=� �'�
���a��yֿ�������O����Ti�jb���O� ��3l�Z�,#��H޴j�r��/�f�F���n�5��U6&8 ���g(���@�%utzR�(����'���aqB	�.|J�JJਅ�TA�ӠG����괇� N
v~*�e(N�$��>y�r1��������o���k��������{���/tyW
c�����S_����9$��L�1�k@�@��e����뵸� �[�BNh�ڸ/����EPu���N�������"]�h|e����y����+�2�Y�in"K|��؁<g?�<#L��G����.Y�����.�=�hS+wL�TEG���@f/.�����3U��d�~�Q$�H4*/��~����e�іN��[�&E���&x~��觡�Y"�l��� ��՜���� I���S�=��s2�x�~���
a�����}A
o���e����)\ʝ�u�;��`˂��uxg���ۥ��ZIX6�k:�+��ׂ�w�׹v[����\d�Cj��ĝM�=�����~��+D)���a��]�vǲ�Wu��3ΕNe��jMB�A���Z\��`"&�/���YX������pU��o`Xx����Q���)Q�fd�_��03�2��7�h�r������읳>ëHg���N�c��e,y�j���,�I���>6����ۧ��'P�w��:Ǒ\�Vx��^���e�̤,iœR�Ψ��!f�x������"po��E�p�)�8�~��i��1R�Y�}X�q��C2I������x��+['��kΩ�Q�<�|�sE��9-��B�Tn�,��#v�z��]���y.�P��|�U�����'��b�h�����H�D�A�4M�ۂi�vs1���OS�����5!8�tХl��ˡ{~�-��#9xf�!�F'���x;�b�C����,v����ְ�s���btz�9e����B�rN���бU��9�7Yn�0@&r�K�~���]q�?�I`s�șl����.TL�� �$��h3�̒~��oo�1C������9=��z� �ZkiÜ���?<��劬�(����p��[�"N�v �vms��V3t��z���{��+�Gǹnd��C�ݢt�-OF���,��?T�Z��;C�7)q��URf2
uef�MQ��Pھ��3�����M���i����j��1J�|Le`-�o;_�� vt߰�oX����Ӎ�0�(2 ���#����1�Z�$�i>�۞�x
r}�6���#���Ϟ�z��k�ѐZx��$���t%ON=ת�ȿ%^wב����P퇮y�[��g܍}R�g�*E�:v��8�=*^M�ߙN��fGHxe�U�R{�c9�x�H�<r�H�F�I���s
��_/7R�w�R���e8��=��d��(oM���vu~d�b��(Hb{�]�7���3����Ԏ�PD���6@�g�مoy����f7,W!S]�~6?2��[�F�[��*��X���_���`��j�ڦ�$����l��,f�fڋr�[�	F�M�f��肩?R.�\��� �y�G��d�>Ůz��sИ��}�9d�����Z#ȳ�_?����?5��T�G�Py�[�癦ݫ�on�k�A�B�b��L�3��[ȆnU�f'؜lu����������(��QTOx�'Mx�����܂8�rP�xz�����A�%��W��u�	p��緩h�LZ���Z�n(�u��;�����-�}"�D$�̻�A��>����>�0(��	Y��#�]-�h��i^�G��~��dj)�u�Pmz�R��R���R]z��!�����vхOF���=��%���a���F@��bBd殕���]D�M�e��R���1�x@�o��Z9��17b�iVF?P��xeN�־Pa��3��L8�SKc������ �q��a����i�Q#��$�X�J���}	�����C2Wr��+ 6�T1��hiu�ȢCv8噞ʸG@����μ�Q�[A�Q�Z^Ie�)��¿*6�@�U0�0KR�7��f�7i��$��|�}��Pe�3$h]9�6�Y��E
k����P�̉�k�9�z�r��]H�5ND��b��T��+xy0�k̀���#��l� �u��/h�C=x��@���b5O81�r�;���e�����u�)hW�΅�N��*������Z�2��=����0�����=���N�J�`WfD,E��͓!�9���oA�� �q�;�hu!��}?Jg�g�.�Ji��Üo���@w>���Z�Q����B��~��Ϝ:8�H"����lV�Ŕz[�I���G(�������x�6#?��Rl����>�M�W+�A�^O�ÆDEf��3_�K��i��=��P�k]�=IPWu}�T�0=.�3ԙD�D��,:$�4~*pl����<���z�+�O�Yf�S|��~�;�d ��Ącؾ��=>xb.�.�i).�EZ��!}�����Uv�
l���p���\��j�1�Z�qS��c�I�EkD5��q�Y�qp.Ь�v�8
�#�_��	���w��rgR_�� ���a�C}���ׁqb�F!�~��s�����*QL��M��'Zm8�}	Ϡ	2�BT� J���o�swpV�Õ`ȶ��2P�o`Z��߷�h<��������F$����N\���o,?����\żzb"�f!=�pj�hB��@�;���v���hh��p���(��`��_��V^�D2D���^込\����t~�S�E�zZ�U��l�	��d�#�A���a��M_`@q�xP�j�;m� �(�.�=��Gё�.�n���G���>��V�H9g��N�/�XM����� ía���.0Ն�(�|X�	=��2àg]�� �@t�=�\�u�\_U�o�2G�D������M��
�=Y��-��ah^H�����k٪<x��d���1����Hc��-����PǪ։{����JXR�@�@v3�P7����;��xTN��Ыւ�.��b��:�O�w�{�<U�y~�F���J�����x���֨Ny�̻Qg��A�Q����oȑl���!N�v�ܟP��˜�,UBS ۳M��������H��xi��q�g�h*&�8}*�
�Q(W"�\�dCǐ����}.K/�^��ʻ�ja�n��w���Y�Dće'ƛ>�i��XH�]c�^�EN츐���<�ȫ@ɏp�7���N�/ο�`�gj�]�\������gWuߖ��M*$B�����CWptG*�
=�g�uFT���?�t!�w�P�,jbdYSdB����M���o��g�R����	���<s9��^jp4�SW�V��y�ڟ��:�2����>�휦ִ��Z��HQ��Q"#�,���g�0Z�"�P�Ԫ ,���pڮ{;�Lp�����kxLu�*��G�f߹���`�z���8頽����:���}���|�ۙ�!���3S��@T�P�Z�J����dp�h��3�8��˿i72!�y�;QK�\b1�s���xv�1ȹ.��V2|Vڣ���%q.x��*�.�C(�94��xE��F�0>:�W^D<�-�^S���ȫ��m"���	Wz{
�L�	+�O/'{�yoК�%W�B��'�N���Ǔ��J�e[�RG8�C[�[y�#�ׯ�y�;
:A�9�H4�Q�'�4<���6+�5rU*xl]����4���􃤅����לS��x!)j�`��K�5e�����>K%���"[i[-4�W��A# H�� JY�|��/)�ñu������اb�ɰ������.�j���	�_���H�r�bM-s���?�m��b�����ߧQ�Y9g� �>��4�Ӊ�hv/�7g�ʙ=d��I ܻ}bD75� �7��w���`���ӯ�J8��)n4��)U�$�G=�����Na߷ڡ~�}9��Juyn=��n��;��(-��W��<�{-h$��Qi�;^��,M\�6�w,a��U�1�h�,d��.�%���eg{�61��e>9��[v�����pv�eI�����ͣ$��:�����ƵW�:������LEI�jZ9��p|��3��m�75 �O-)�J�#��^
}K�+aZ��y�gdO�)�"%��� �r[UUj��.	b%�''_�9�A���=mW��M�й�0�=T"#��t�GH"�����,A�]�Ȃ+�M]R?ٶV�
�H|�Ma�t;��xTL�"A����+�q�օ�ف+y�%�iױU�����۾)���)���7����m�u	�MP����P��sZm��?h�X��C��bR[IմK�uE�oܭ��	�v�Q�)6;��<E����~8'�]�Q�F���o(2̦=�I�JZ��'����f^�'�愇�f����FB�hr�����}�X�����F��%�{6��Ԧ�M�%Π�
k@��$=cTP�p�P��Eş�x]0��_��ϼv�=�gs��r
�0_W�kUD%'�9�yX����m��)YG +k)(�m���GI!n_%( ���{&�T���#�;2��{�C�πzg�Ґ�B#�r� b��~�(|��y���W��j �^B�L�`�ޢl	i��⻍�Ʀ��f^g�D>�z�9Ȑ>�pj$��rM�6ͣV*Ң�(��/I!�X����d�+R+"�ė��0=�>[�Wv�&b�e�t%##C����^9ò���f��Qp��2*�7�ν�+�[$s��}�J�/A��=\{;**{ৌ0hFP���D�2�#r(l�y�����:��B✩T����Z���3Y�"�lA���n�ll(0,q��'���̑�Z��ٵ��i̮/t!�*,�-�@%�2��w5_O�����:�K7]˄	�`�V�R���2��z<����M"2u�����m�(��!����	}[���LH�ŞY�v��$!����x&�@F�ͱ����D'�@hb��&pD��Q"#F�4L�3^�}n�¯{IԚ��P�K����mS�A|ΰ���.��#�z����-�
�n�����ւ�-�8�8�A���HQ=V̇i�����!1�VO;?��D���>�
j��5��d�t�����Ҋ%�Q*���?F�Ze�r�"M����ԡL�2�ć�+G*)�-��?񞤢���X?�m�6�f��Ze7b�.M�3�����tU�F��DE����/�.�X87Z|�g:�w�WIdy��ܚ!]%�[��W�XW�@���c�E1 �W��(�\��n��y�¹�����1��[,��Q���*�K���B3��y�{�sƷ�K-$��`8at��
��f_K�*_��+B�i-U/���\=��X%����3�9eRlj��b�͓������疧ڵ����6�����Iu3{�BGۗ����o$&T�N+Յ���_~�(<Yz�̢c�Oc�|�+?�y��Z�lxE>Z�Ff�����F.�L����lq�l������
캏t��G ��V��73�����
��ɤhk-�5�J��[�A���x1�[,\�ј��-K����k�g�OB)�.����i�c#�ak+�[����?Ā�b�:z���)�׈���|�Xݹ��@�1�뼴�h���W/z��R�澋��n<+�q�UF�V8}�o���53���<��'�+w��@F1�Qo�[��)y�0��󐔩�=�y���c7>u�ۯ��� ̌�/E�>�	�t&�4�N����X FB'mi�Ta�(��N��*d�ݰ2'e�-��{�ר�r�ˆ�3G����E����=�=�+VEK��uV�%����P�A�I)m�= �"K���{�7�Ʌ�@@AUA��0���8HxI�I�N�U����i;��>�
���AJwU�y���9LN�QpObl�����:V�A�	QÛ�Q�l��0�Jv�W']8�*����~�E-���*ã����UQ�|/	�f��KV����˂8�R-�^����K��lN�q�Y$ъ��#/[m� ��eq.����s���7�m�59N����s]`�F@	���;8��a:��a�"�/o�k������q+B[fÉBw�}+��),�0�O�$+�0l�1��g}��7�f��<��W���툚)kܪ�� ���:Y�Ez垆����~H�d'q.�O��0��ײ�z�tZz�`�� ���<��N����R@!���A�T��&��E$z�����x=�9$��VǬ���ꔦp@�W�i���!� ��J�h�t�vsl`�P�.�p��� ϗ�J�z���cTZ�?���ڷ�^	��ͻm'���D�ܶ��Jj�{�ֻq���A�?�� Wq��|H�2-�#�^�V�v�E�$�u�١e�c��fm
��f�4V��x���	�2#����a8x%�w�|*4����;�x>K���ȵ�X�ܭB�|�%�6�B�k���1��ay"�='@ByU9�ZdQ������d�pMf$'�� �_]��ȼ����ȳ�Aom{������jl�p;����$���/�yT��`�S���~�1����x�H�{�����İ�Ձ�N-�����8 I������弯�O��񢥑Fl�}�,����a��1�{�H!h�����,�ӣ�$lU��/��JG�n��,-_��Ȓ��%,��_k�ч��U�5Ȩ�2j#_U0c�C`���!�(����&AsU��'~Z�C�mg��qO��5�z���H��%�n���]����4�윥9���p8{8�o�|�G1����*uZ�~˻�N��1�Z��&OG��)�`��S ���#�sG0������r"����(x��1�`)$1ZsR�;�l���*�57Lq��#�dL����8��.X�����.1����qx�@μT������-�0e߷GE��]�u���(F8��|�E�0�r��Mm#~�/@�j��e��(���P���&�]��ur�s�E��A����YhMw����O�%(H��\O:�f�_�o(%�K9�>�t�>
u����8]�=啤���6�����i��;����o���	l�\����#&k�u�LA-���=*���$sMɁ$l%DC8#�nv*Ä��w�pnc�׍)�z����W6�j��}m�/!�{�:Int�r7�M���+:-_����V��
��H�g�L����7���nid*8�0�`�1xޚ��=��L��R*C�"�������W���L�������P;hy8�(�w,��*ۚ�,.�~K	���A�9<��o;����W�Q��� �#�z"�v92;�77������T�%L_��}�ٓ�&2�[&��/䊴�{��Bñ��6��o���\�c��U5�c����		��A��3�<(Ed��N�P����n>9�1G�2��wX�[���@"����yEd��tW��D&�ơ�"�,|4� h��?`C��!\���R�ڠ{����:�:r�̢zSfĚ��HB���v��ݠ�zq��]��m����eo,�ʢ�=���0X9jg�!Ո��P���1%M-���l)X��p�U냜�&q�)�eT�,F�uij?�3Lrm(W&	ړ���Q��+u���S�1w�}�u�x�E��jLPeb��2�Gl7�o��5�rl�4!�	�b�7Bb���emɳq�N��ퟄ�"@m�l�!���|��!_����'Y��
�����)�R���_��;y�xaT����v�uDNg��C�`R�>��.1>�|��J@梛r�л���fdJin+զzf���}P�7�A�nWbRg%O��`H$����1c{�)e�п�2ׇ	Ȣ��I��Tt� �x�8a��7��=��L�JR�?p���x�'L"n�NTO'[E��q�����a�8z��a�-���N8�p�Oq��4��?x��aS��N�x��s7�'�A=#0vlQU����;�8�=}�%qE���@��P�L������H�/��bBn�/���n�F�\���q<q���Uhq¡r`�K2���V$�LMcb�p���e�j�h��s\�v��X��.�̛����Q���I���#�Y?�W/b�b�����ͱ�a�9��ݫ��-�jH];��x���\,*��~�H���i���ı���U���:���v�q�������:�y�j �QI9<46|�7ys�F�őa9I�s�xVX*/k,h�xpt�(����-qu�t��o+��[�Bh T6{�q��g
��[����a@Y�� z�4dc�l��	I�P���ԣ���L!��`5@���Sp2����Q&�_����Hڨ�pO�Y�M�p^��3������}p�h�����"p���Z3�ʉ����p������`�����cӖ�ŏw���\ѣ��a�)���]�g�8=��*�w |�Ël�/yH�M/ѓ:, �ob�W �_|�9�O�����S(	oR]$�8�-�"d}�t��p����UD�f����4&�\W�Dy�K��~Z��2�T|��8T1��y]\p�S9��kZ�?St�O[�0����z>Q��t��=���v�H;�):�MO��s>�޸��<_Ɂ��!=!����%S�6�d��L�B:H��o�@I���0/5�0�n
�����+������F�c���p�suH��&I�v�A0y�c�d�-/Mظ.��
W���Y�
Q�^H�<�Ә���W�3xb�_@�+㋝`VUi�$��nWQ��B0��7�V�e?4��V�F]��̔�[�ҥ�m��|�[�ɏ�^��t�K�8w���� ���b5���%��g�C
S�Dը����r�C��^ۅw\�0<<,�b!�)c��F���>V(2�=��{hx.6*	���y�(ɏ�d����UF3����9�/�_߇:��7��R�q���6G\��n�{�aw~�&�V:���M��6��aڀ������S�M>>4���ݵ'-�٧�^	:�İģ��d{���C��¥	�"��t�[q�t��\VYTJ�I5��h���Q��Im��Xz�;�Ծ��2�BW� 7_��t�l��h���	6d`��	��Q��&����=y�+Hc�5��.!��[����_�$��-���u����X�R<?;���i����y�x!�{+��u�z��`�*�L�ό~�nˆD���N�]���ҭ|�O�ƌ�9Due��LX㖷6㪴C����¬|� 1�+(�u�z�׺M�3x�k���vf�h���#/+=V@}�: E�Hɷ��/�0��K�vRD�ctRnD`�Ud$v�\�P+DY)xB���
�guV(u>t������9s=fu���"uݿ�,��ݪp���r���u��q?�z��R��4-�,�cb[�����j�gP�a���T�k&�~u2\� xtN7�6��������e`��ҭ�=�/m��M�����]�Z�U�}ޞ9�v2��#�x�fOTut��r�h��R��J��	V���J��eЍ���S�O�qV��0���ȃ��\�ְ�".?�;�/A�v�j't���{B�V���@J���|�g���+���pl�U �_��6�**�.�{�O5Z�� 3X�
4IQ����(�,(qW&i`~��������ٟYoL�w�'Kaޒ�F/`����LL3z��$�(�/5��Y|�O�
�qXRA���:��2n'�ac�����gL��Np;���V�4z�gt��N�o`��4��`J�ӽT�ʗ����@"���o��I*\���<�ڪ8~��R~`�b��f�Xe����N&b87 C,�����G��P.;�H5�?��ӛ�~Q'�/��V]5�g�e� &�]oM�Ӡ/�9�aX�k���=<ûy����N��X�I�L/�q�x뼦�ـk�k�WVt���@
� �(��T5���+	�Y��Pe�#w��d����T�u��k�C��{�K�'`~Q0e��ʗwhwP��jH�껡��F�Q�Y�%�[b�>���G�q�;���E�ۦаmQN���>G�r	��7�?E�`���T������k���x����Ud��~���H�w�ĉ��
R
�i��2Hd��V�A-�/��,z*���L��Hoh��Ļ����s�$�L������U�GJ���p:r����7E4���s��xl¥$4k�]�9[�:�M>���=D���(C�\���x��X��6b�\|�̓�n5CXΩ��,��7/ә8V����~��i�U�M�W~��+�\4�9����bꅁ��ӷbG�<���K_<*��U�	$�)�%��Z�����@���Qy癝H8g�GF���>0���E�3CYۚ<�Ye0����Y� ��ċ<b}��f�h���A/��y��ķr&ѤB{�`(�S�ς��iM/��������|�bR��G�L}��Y?��	�<��B�aJ���Q+#9�yH�� U҂-/N��!.|&���]K ���R6����RLoeC��a#l��Ѕ���ń�m���IEUo@�<А�k��hJ��B���y!�e6d/�1c���A%�Cg����]!G)�fW|qG���d�8"�â����rO0D��������;�3\�����T/�aP��u��R��5���V��h�j;T�D6L���@i������)S��	�^����L0$zWcf�����`��.K'r���d���e&?]]cS���mڞ�&2�mZ(�p��?��$���=�;%`n��T�4O�>�����k�'�j?ʢ��Ui�������qR��Gײ6��:�=���q�`� ��sg��2rp5Kyі6.�Խ(��b���������<�|g�6���S��?X�㻻��8@�b ���'�i�CcѴ��F]1�ޔ�,}u���r���ԏi��\�2����OtY*���T*���
�Ȓ{�]�e׎>uc�i�2�և8�-�gJ�����|��������4�XN�������1���I� �����f[ȿ���B�t��\M�0�d���;:���綊�w�~�T�6�Qu��J���>-ɏBm��w���c�K'S�5��Wng����	��>��z�ؘI��������D�*�]��������
�,^�}�m���/g8��V�v`/.3R�6��a6�|2�y�J�,g�1nq��S�=�����^�^��oP��0�U�s��#n�o2/�q3��j���K��B��}P�%���#�vI�W���!l"T�r���(9�KkEf�%"!���:�rc�X�c	�~������(��L�r���N��*H�&����'��`H}���}S����G|.m�"�B��â,r�1�N����PH9Վr��mmb���2��<S����(/�s�co+w��v��=I����G���U3�({Ǝs���7*ʩ��(�r��O`�`�^	(F��6%�s�QY�t�S�,Qc�j����d8^�\��Ϡ�d�0��L�<�����X�|[��u��[y2��j�<�4��G�$*aPs����H���Y*�.���Xh�S(\"g<����9\�M��B��1�R2��C��E��&PDby�+�M��hP�E}n�����p<�S���^�6�������A	�;�$Z�c7'ϰ��L�A���I�k����WG[�XR��|�e�g�SU�*3Ø&3��(/��(J���A�}z5��g�ᖮz�f)h���?{@f�d�<=23�E$���g�Sj6N;B�̜��7U��˦�ph�̝�ZR����SǏ֥���hS �C7����IlO%>.4�#r�K�sNg��.�Զ��9&�Ú�&��p�l����p�=���Ė��[��5��v�C|'�����0�%��w��?���r�:�Ō���&��J��f��<7���^�\w0陬��9vO�K,�&�������Z��,��G��>���:� �H��|:y�Vx@���_^K�>N��3f�~�]�Y-������5���f�q�\/@Wa:�Gֆ�q�o9c��ή����ְ�=.�t�B�7��zL��_��>(�B;s�#p�1�HP�Q�3�>5Zl�*n��-t�YTW�2yS���$�i5s�����)��.% N!��St42r�b���ס̲��#�Tc�{^����x�[�}�ؠ���pzD�?�(�w'���&�1�D���w�8��?��c ��2���-��Z��f�� �3�M\osɣ�T\d��;�"o�B\�no=OGA�΢�S3�w^��W]r�O���f@V���[RN�ә���Ft�d�'0����S.O΢OU���H~|#L㼼Y�Š��Y*�%���6�Y�k�ݿI.ܵ����BI�\iq�Q�cz�ر��t�̵�`�҅�GvW"���a&�39��N�И�"ƌT�%(�ȹ�Dqm(���z�I]����R}�O�8�b�3������4�led6+���tj��#���Y��r��n��n���~*���q�ڊ���w��.�7ƮZ�a���,S���y����in�#6[�&��'17����.�Z}�lm�"=X���-(�U$��%�+WT[��O�e�:����s<�e�}�f���@ sHp�g'_T���� :�t��܏��IRwXg[ ʴMj��G���/-�������o�;��EV�;��J�
$P����0��!m�&��[4������h�^�wD�*9k�
}�>� ��CL}Y�>��w��,�9d����,"�܂�]9���q�	?��a,ѿZN�y�v5i<2�d��@��엔� �?�!|��T=�����($�WO'�:7����f߉w{�Pp��N��Nc���?�U�4)��۵��(����u�D��\܀%p2bk�.̵g�] �SGhe�R���LY�anL�t�� ��mk�؉��z|�Ziy��w�t��(Pv��F���9}�Xت���L�v�Ǣg<���R=���J9Q�TL�N�	7 ksjT����l�Z슴��*{j^���l�ȇi >� �-�앁���������􊯓��xcJ��ܰ�e���Lv�p�u���i��
_�S���X/.�,�:�H(M�)��ҷ�5S/{�����fm���*�A��y�����d��yHē�[��ɗקF����)�
��&�q,=�D��Y-�듢ڢ���_MO�0�"�n"C@�8>�9s���Rv�,Q��u�����O�V&邆�Z2���6��<�]ƻ��Lӽ��L��R4���`�X�,�mӉ\1��M\y���9�L/�B�s�نj{$�U�I�[��w�N�$9z��M��:
�p�ڠ��*A�I�Ә-�ân]p�b/�>�����֙:r������Me�\�!��$�`w�sq��^��#ξ���K���OiU,�ºVG�MѾ�F@F�# �t��n��(��vz���<��n���fy`��X�D��@�F_�Z�݅��w��m"�=�"/��Ժ�+��4r�HY�GS��A�Le��;�<'�@kbr��cgM�6������;��cN���Ȩ _�d��VrGM6��{����.��_g7����>1�V�ZT��z��/�xX���ôQ1�a��v��j�7����~0{�uA2�cW\�s�WZѷVhqw�E��Ƒ�y��`)#�l��ѷ�������[AW)Am j�Y�g�p<�C�i!U�{��J��w��0v�x��1Q�b�u�픥�O����Bj����� '�j�'��0v�L��(��gR�ŬC��4�@Z�����ׯmԓ�� ���ܣtD��|����?��;���`�J��2�
�m[��AN.E�6�p�@i7R����"�\��'x��%�F`��R�ݼ!�|b�o�?d��.^F.G'e��X�U�����.�Q�W��3͕W�'�-L�'lZ�0���A$x,eY�E*��`�x�u�<蝡��˩�>��k�ʓ�r�i{��CLe�-1�^(�v=�NP���v���M)/�'�*�����E�Ś�n����+AQy��_���-y���1ץ��x�Ϧ��|�)eX�ܭ�x��{����ܓ�Hڊ���Ĩ!��l��s����B�N𞇧����$C���ؐ-&æ�Ś���1rC=3��L�Ex�fՅ�뾘E�/���>����D�GW,�șOoT��Y.����P��ڀ.k��X�~�ܨ�L���<1�������[�5k[�-D~k�a�=�h���6����}�-�N�{8`Xrl%ߝ��?�]��1L�S����ހ�K��Xm��� J��"b��?iPy�fr`�q�x㸶D�z�}wny�d-���c��O��Y��X�`Ԫ
���w�c�#%e �����ʈ���i+n�o�D'�I�KH>�dQL'����$?lI��+D�@��2��*�}3��f<��c'��m���r��@�$7�m�����u�rF|(I�,X�]�=z!�_��[@���.�l�ب�md��"u���ET֊��l$:��I�o%�u��D��������Bfcm���'�I��^g��Qa�팫��I'[�YK��Gh��6N4����!���?��m
���}{�*<�����U������˕_���ɞی�fZ)dI���B蒦3��d��|2�t�S��P�>D�¶�	�Nc�-%=��g��j#p7���(*LRVÉ�۞�f�`n�9�A��eR#m\<�x� ��Q۳.طǁ��s�/NȦ�y�u���S0e性��bW�t'��b�BP�6�U~t�3l�eY!	t�,3t��z¯��5�L�,8K�Acr���,F�fst �S���GI�=�3vq>t�,�$[w~�h GӘl�m)���;�.�Xs6����3�H��!���v�:��[$$G�V晖)�{�Z�*���Ж��#O*�̇��6�V64���{��/�넟�ﻎ�]�?V�c/�͞�	��Ra���H�}8N��Y�hqx\�I���������%�O	iCGUN����S�q�ж��6�A�]��G[D_(�N���1e�>O�������P/tǿ�U����[?�(1��O��n�{�"�A����W�7��H�"��H�V�	�NzǪ�g����X�Oñ�Qm�*��\�Tpx��y��Z���O}�%<����)���&?��e��bmyb�V�8�>)��Ss,u���r�;�aj�6�s��:I'�nq�0(0�_.cJ��z��j�M��U��J�F� ��֗��8Pk"${M���^��<'��IN�ꔓ�{�_�d^'֒�λ���'�]JSP�^�@�zN������ђ'�!˯qs`G?�ƾ���74�h�h��JDO�B� �
(���l�q��|��\U�N�2���Wih����Gw� �V���H�˽8ב0 nYb���k�
vV�����p�=ў;Muُ����Y���O��۰v+#�su���#%}!����DI
v[Y9������.�MҵX���ip���h}hC�8z������V�~�QM�D����*$�{�:B��~�0�\�`/ *3p*���3�=��/��|�`!���A(Aژ�����!>��a�IH�g��.G}6�L?��9�v (8��,uډX�.�_Q,��5Q�"~o�S�>��0U��pO�K�t�،wjA����aF ]v�d�I/R5�����CŲ�N��qŨDU)�X�|��)�P��=B�e��a��%�����1�?��M��ӱy���{�Շ��&��)򘰠r�%�9O#N�gx;��%�K�i%��M&�@1����T��ٷy��)W��g��������!����VE3τ�e8.EL���Y���Vn����s����@z|���	uԌ��k�"�VU.0�c����.�Ʒ���W�r[�MO�M�����X@�q�N�S�U��N�?nT����.��������i�x|�Ѵ�UIZj��ЀTw4�Z=�n�c�Q������F�įR�_�Ia��g�#���i��7l*�����v����+�rt�3EC�٣Zy`�o(<=�B<�`��vT(S���ɦ&s���jj;M'��EJG��C���P/�ǌ#���T��B��5�3�r�0+�5�)�^����#A��H>�!P�p���R�<H+v),�^�Mxnv���\7ߊ֏��׍�˨�j#FV�6���XK��k9�1=��Qd��W�(Y}PK��zT
�'@�����6�Dʹvp�0�=ѡIa�ƣ(�"��<���t�h�Z���,�8�Ra�g���fs'�*R8?��*i��9��9�f�}���:��S�l�T�� �g�>�G|�RW:��"U��F�/:��!�����\Ĉ��uB}�����.T Ҋmk1��H:s�tEa�؇i{^|�YFt�h��}�JS��\�)^�u�q�5��7�]�a�F����iqެ3�o�,���僻`��_�[����O��i2��i/��
��Z#�����\V�w�҂�9lC�p��Q��8\�I8�b��A�\%��t�r!K����_�f̃�NbR�s¯��z�̘@d�k�U��:���w�D����^W�mA"��_�O�z�jg*3�Z��v׃�^�ʜ«F���v|i�"
�ϻ�#M>�g0֌G�-�.f����7������Y�ނ[j̉�;��Yj|Yk�����E�ڣ�]�J�S?[`u�����	��)��2��g[k��Mx���1fI����V�������g��o�v���J���^��ATIt�a7k޳��=Ʊ�gTy���E����4sq�|�#VIj<(0��U��I�"� V9d���δ��<1�	��!��q�^u�B-�4&��3��'�7����mn>&�>/Ǵ�.��R�͘r���/�eL\��܃��]����֖�tg�>C�(�/���/�n�k�d�%7S�+�	�{�}㳉�f|�p_}Ba�Z�'2/@w�5'�Ep`�D�c��rOm���k[�sPH��iϤ����AR�qf���D����$Ûۣ��=��ޒ|ש���|�d�
e�q&t��=�����C��Y\�ڞ����B(s&A	Ӎ��L_߷'&�W����=ڀ�X�����鞴Xp��K{_sz/�i�A�U�;
��m��A���;6G�'|�p�%O٨ۮ��z��l@�n>����f�:�Qo�9�!n�n���>gc%a�V�3L��߃��-���=p���k��Х���"�['2���I�)�sf������d�m�e�fs߃���e׋S�NV�w���ZN�]3��'��L���)���9��F
_�iI��|i�l�Z�W��Q`ct�U,����{�|Ն���b�/b.��'�>BG
�S�e�����"t|�>�d:��:��>*�*	.�m�_+�9n	����9�/ b�$�ުߎ}?e��� �ٙTQβ��o&��=r��� KWo(��B�8�a�!��/��Y�X���B��$��G�J$�;����ChN��~�<���d�>V�d��	t�=�Y�5���S�-)��l٠A�x�.�_��ȳP�=�v'wn4�y��< ^�t|2����ړ7%3ƫ�G� i\ec�`,�K��r�,�Pr���j��;��ϱ�!�n�����_��Pg��L��3���y�v�x��݄�C;bl�C��=c�#_^�0x�,ր�Ӭ,�6% �t�Z�RQ��U[m��?��
����fN��,S���b���y8W��6#d����a�xn��i^�t��',�(�ϕm���d�R�]ɛ�&��f8k�q���C�;_�gX	��y��{�t��j��{�$��
E#�1A��`�%�BД;���os�
���h`D�2��y.<�#�[�<Ng+���eaX�X�<�p�d�[�&' !:T�M!E�_\�t�y��)��@�~�f������fG��FδFK:K�R>m�W�-ђߠ��D��m��^��-k�Ε��]����T�Ƕ���ƫ\*}jQ��!\w�KK��X�;��wlvb�NB`/�R)�o�½�{��x���w�� ���a"�EiK������(v5�(`d����ܔ0������%J��9�l�L�Al3����f�I8f�H��Gyl=�VV!)�������x*��M����Ax�O4����_�OB�sϙ�vS�@�H�B̓t��u6� Z����,�Ԫ�Y=�䱇��Ŭ�$~4�ҏ�]fDa�Z�	�4���/uė@������̃|�N�ξ~����b��\_���gWI3rF�wWSQͣ�[��!��`]u�N9�aҢ�`�J�`�QP_��nr$~���v��f/���X����$��m���c�qG�k��e��CR�u�?R�su9��0��w�54eN�����| R	U1�nq�Ŭgm\j�ߡQ�/*�z04Ɯ|x�P�w�b�؏��E� ��U�0�a_�i��VΌ�'���mjӼ�k|��[�Ŋa�n�.���ve�l5�NP�����Tx8�6�u��ƃ���.f��5�k]��'�y��Fr����)�7<��@ E��`V�}��wE��9���W������PQ��6#�$V����A�F�b��}��;�ɴ��'0���&��rkV�eCkʻ�^�����>)f�R��J��U�:B�����.�rν�W�L�Q��4~n�<�p�����& ��%�>g{��=�G>!���d3`�HA
I���I~���Bvk��hG^��d`��u��_P�5��|n�󴲋��܎C%'�9�;�>�ɶP�^�Qk�����d�XU��@two&<9.�z�^]�Kه�+�Tu�Z�=��� ^�~�������W��l��. ��V/�90
G�N�;K+���h�4�=���?����p64v$�yRJ_���y[c��m����){Q�T8�z,��8��3����M�<~K�`���.��.Rxl����J�}����\��Cǉ�.�`KJ�r��y���%��u ����ʽRy�/�����o�M�ב�V�v{�Lţܡ�N=�W�۪g��N ��F8�ǘ�c�=���"ŭ��!冼����biH�E`)-zy�^�G �,R�ĸ��Z)���h��	*�Jj�n|��O��d8"ծq���ގ�.�q��W�k&�'��7c����V~�d��l�Y��dI0e���3��0��Hd��jtB�t������m*C�'=7��i�Ͱ8e�6�����ϭ��]l���a|zu9�WMj�ě�jm�nwO�j��CA`
ߒp\��ݏ'$Łf<���Y�b ���i�!@<�x����3�3`�ə!�?��jݦ�J���l�߇Mݮ©t��ki�TrW��X�n�ɽ�qaV�<�a�2?�	%�<yǸR  4V�Ɨ�0�B�`|.�{�/AX����1�o#��P\��tD d�$�ئB+�	Fu�X{<�����������l�������OK�ٛϖJ���bj��F<!E�����,�����2I'�� D���B�p�G���v�)�Nؚ�����g��B�2�rhP%��frG�cr�f���o
Ђ�^��r%��|�	��L"UM +4�Z���(��냫�/ 'J�b �����/���`�Ԟ�iC:_�I��r �e�3c�����s�����@s����AU3��%c�ٲw�'�,���P@��Z8�YV��{��ζ�@���� �Z�-�J5���\�C)!V�a����-��̤�{O.�յؑ�M-�/�_��c�@��mԹ�B}*)n�X��.�����*n�����os�� [��Q!���DcrD������Ȼ��~�M�<
�Cu�t�}�ݶ�V�T��Y%��*S�1Y"cے�t���"q_F�ރ�b�ǯ;�xe�op��m�|/E�����)H[�C��{Љw��^g��Bog/S��y,�zl�<+	[��L�Fj6�ޱ��x>����Y��f՘�G�\@����0���|�EC�����ns-���r}���((̙����C�����<���/ץ�o
(	�#x�f�4��)�9���G�E%7^��w4�{$,�ɵ�3�\�E���I�g����4���\}P�շ2�'��^�OD)�o �v�ܫ�j�`�a�PjsP��R���k�7V+?����<ka�~��[�=��R�c�0��=}��'\��K��js��4D�Y�R�un�GW^�^�vA�R�Ky_뀠�#���{��]iv_��A7݋<��ӱ�me4[��K٫-B�ʹ�n6A�FG��e�$�����K��@���S��B|�jn$m��3��%�
�i3�Ž_��*��~�s�v���a)���4'S��	��:^Y���f{�,�v�e�G+�N!�(����i��'��^��dO�0���%5�?)��)5���?� �.�\K�Sw���� y�Ax0x��W��ބ1d\�1z��p�o��q1���=j�
G�bk�Rƹ��`��)�'H7����#�g6��<���e��E3Y������߰oFt�R����� H�ў�B ����5�[J�|�DF^d�/����2�	'Icv�8�q�J0_
��b�ըt����Sj.�6���yS���s�t�7��|�!h"p���o� �W�RY˳��� �Dڝ{�����#cN�W�՜B0�''ꢂ*9Ѽaw�D�,�1�U;���n��<
�jxґ���*�ϝ6J1�ck��g#U��@��R)4�R^�S\�d���trА)�C	5�N�I�0��{m5���~Ћ
�����f���"`+�~G��P�J��]s�Wa"�8�発L��&Ϩ���e���0��:(�=�!2rvK����h��}G'c�u��7����ޓ�^����u�l�^=P.��a\���U�|�>*?&��Ӻ�;��\uc���"r�p��!3�)I�S�g�U\��eYH�Çy`�u�iMUL�n�Gg�oN�ܵw)�,_�x�2�JZ���Q�o� p�]��f��.��r$�MK��3S8P���	��!�:}@����q9?��|<KQ�{�?E��v��V�c�6�ӭk�b�jS�̻�Уim���[�:����t���� �g��As6��r��A[�=_L$����ݺ3}�o�?�w�e�΍*vµ��|�b�|oj��1g�:}%cFS"�5�  ������8md�1�ܦV�_��v���&���Bg�|��;E�i��$X���$c�r��1��F�6��JF�x	���g#Pi̥Q�Y� j �s+���"k���+_�wLX���:S��Rk�}$��"�-j��<~�\�x�=�g�
�%8)��Ǘ�\jjM]�¦c��1�9�<Xr���h��bO!��5_S!z=D�$�'�.�x1�v�7�G��*-v��YWR��ŝ���k��f��qP~�1h.���S��������s���#��R�sT�'�����v�����F3����^O��43_M5�i�;18��(��K�	�+�C�F*��!�eP\m�Z�d�|Ј�B�7�v�ҕ^���v{5!�tP��')�ꛕ�kΟ�Kx���4,�8��*���6��o.���_����"�n���_A��ф�^��΄�.%�3��f���͂O�&�mz���lt ��OF~v�Y鑓p�`���΃IZ/�Wƣ���R�D
s>۱�#��$�c��^D7T��� {����)�k#��~5b�ʗ�����@X�����j�绮2Ǧ��"Q�w�� ^a,��U8:h���Ǝq)ü��ŶNnu�����R�a�{��"��߯����0}d؈�T��*G�4��3���r�FS*N]�#��o���q����9���pZ��w]w�Q�|վ���}(��+�ㆈ?9Q�W�U����7��]�V��:XL^sfe��,DHSHTGL�a�{�xL��ίx<>cƞ$I�8ؤ�-�����O��ԥFcw�	+�f�ǆ�ר��v@LCV����X�+��@��<���(�K`3�Hۢ{��B�F�
�dg8���ZR�E`�Ⱦ� �ڠn������^X`���\=��2���-��Ȉ�|_bTc.��&?ES7D�cޔ�Єc��)�t�`i|U	�![i醣�/~�r�;rɓ {Kk01A`���X�O�Jko?��y�P1�ƍ��1��|R��A� Î 4�Q��K�Y���T_��k���� 4t]7J%����D����~������!���|pxTd4�pA��aa�[V�}��r��|��_l�3�fe������}\�>!ss�5�q�;�!��۵[Or��⒝��M8�Eh*߫T�_x�b{ˈ�'���(&���`�u.�-��1�F�B��5�i/�hf�n4ꮇ'����D �cmI���T�o�e��Q��_��4y�:��[&n(��y����5�f�
��	C^Ԍ���5IeL�� H��(g&�D��"�@v�׾�sB�W��B�y���``��:��*����s8�E�|���N(2V��H�ׯa'�zM�Uk�W%}��57Z�N��&�])Mck�r/\��m�x�Ugz�2��$�,v�G�M۬:�։[wC8dW��0�z���)� 4�?RfX�ס|���8w
j��Zs,��d���EFF1�]�f�k{�F)i'لU䌵:�MA���4�ͼ%͉L��e�ZN��x��R����+�L��zS�,�(���$��p��~rTx'y|����9xU1��}�z9߽���K&���E\'<:�������{��Fj��zenWAS�0G�����j�a�O����J\E���bpe���E�H��:2�]�|�?�iK2�^ƒ�;���]���cx�.	T�P��nD�ؤZj���3W���3��"�����(�O�X�p�a�����P�t h4Srߕ�|�&��j1.�\��ڒ�w_ύ�S��h��vt��N Z��u�ZIc.%@��i̵C���=�׉�D�<�CY-Ȃ�-��M�t�������~���Z���;ON�w���H�����d��{��l�����`=B촂�K��O5�S�򼯹s��y�'8O����0?��7i�='� "��<zs�����~�Q�����3���Pc+�����S�`���c���T#�q�I��P.�W�FbVt@������IZ���W��6J�W�+����%�,�+�׿�p*�Z���!o`��.�3���A�1ţ2{f%�P"y�b�� j��zc����y7G�c\o�r����bTD��Eȯ�Y��� �H�i�X�z��82�ѧ��5#��6�N�c�Q��-Y��+8~sWѺ0]�4�?�D%G��Y���j����'Y��Ekv���h�����!A���O��?{�o�4kXS�h�N��ſ��9U��C�h8��oi�r��@�h��d�o���ӄ9J�#��r|�,����2=��AG�<�w�i�L�N)�����.�5�r�G���[$�
/s����b�D�xem�����ZI����YI>��僎�������h�+��N�3+/Qٱ���Y���AW�����6�fMt �3���9����e#��읜���Ʉ�{�e�C�X�#�D��8���=����*�~���؝C^���o4O5�-�(�_-��S)��ؾ]�vb��a,L�i2�(��(L���T��t}B�4?�ui���3F,�����
l��4-$�7z���u�~�z�1-M�ʠ	(wڶaݴ�R*q��0s�ԪO?f
�tGq#�-˕���\$	L���J҂Z"�@7T�,ib?5pʒw2͹��r�29�E�/�����H��֠�ԟ�M�$.Ȝܱ���/�1|'����t �V��~t��2"���+ɞ�sn�?֠��]o�n8JmJ�>.Ԭ���E[P�f��rnn�c)��^�Nw���k��nK��2��Z�m�����N����Io5���F����˪��������d .B?h��ux2� ���`�$$���uv�`'ْ�1�k�(��y���u<)�vC�[e�������g�y��H��z29@���t�!�M���1�0W�L�)��ˋ�q�C���"������:o3��n(C��[��SIB���ϮɵȲ1�`� t�v:�(/Ğ2�d�r�V�EX7}r:;ՕB�<c"��O>�� "��z.�Qo0��q�d]A�?���F��2�{���Z���*N��si��$k�~�3�:���L��6�Z����>�`���Q0V|f�|7J��8��o��[�es�� c�B:5&)3,�����+h���{���Ӣa:��60#��I:�=�Hc���x�;-荔mI_��\��`�Xv�B�	d_v����1�qS6[���e��W}ͅ���b���3�	
^-�}�Źɾ��,~��K�x��rݪa�h�=h�6��*�B�(��"~��n�q[B�,ezz��r�g����;g Q�c_#���q&
GX�tQ��x��q����������ST�{��8.�A䯫j�ل@�֎W1ᢠ��ƾ��	i|�ꡮ9�-)�[�?���:����K��W/�E~��~����(FA� �H�;c\�<>u��|�4O����Q�+���H5����.�(h挲Y�O7��fx���$I��!k�����1�1�,�]Q/�����R���*����Pg���:�L��1F�1��Ӟ�0����AT�Q��Z�QVV?I��d<@5�{j�Ԗ�[�$�!�ǽ�B��:�$,s����c��gV�V�=<m��YC��ꏢ�BS�}��Pk�>�n?N��:�8Kae�Uޡ���������g���Kp�2���`O+O�6�Ϲ7?��&�����O0H��&>��f���/�h��P%&��r�I��*�� � ����bn.Mń&gd�����^�h��w�����;�n2���L��Kg2R�-�����PF�[iW�@K¤��D 2n�����h�_�T+�N.�H��\eg%�a
�}�ԗ�z�U���,¨��a_��� �Q5��0'n�r2>�Y�
����7�X~~O7!pҹ,��t�D�=y��$��&�r�c7�L�je�4�m݁�r�ݜ�Tj,U&�D�sĺz�y-b��e�N����j���NR߮��G��}��Ch��@ ��.8�^o�D�f��Y�ؑ;� �T �+f�C
�#���B��WA�A9 ]�)Oy��Qy=u�]{Up�_^`Z)	)��ͦt�#8�5��UtdS�������Faҙ�$K�~�);2����JkFe�ub�f���� �Gf���+���|C�Z����R#�[�X��@�#�A(�/��aZ�c�!��GBœ���˳{�+�9p�(�~�^7|cc�[�����u���#�<�͓g"$����6f�����+���s�����~?O�B񀮰��1�r_<�(�z�1׶��H�82BH��Mb��1��M��?0���lm|3&�-7l��c����6��i�	��`�}'�-qȌ7BR������p�Я�����=G$�/�����5�3��� ����� V�a�����E�VX��^�ٳE��㏪�5@T�-dJ���IR�6
��w�4������t/@���A��y;Ly�	�E%��p	\��خ�93A������q�!'S�گt�av��Q���j1蒝����wV�"��g�O�I�l��)b$jS���z�/��5]n7��1+��'�0I�5}E����NU�($a�"��i"�FG*�d[���o�T�Im�/�8���cT(�
�6��?,B.P�/[�����P�|XZ�;�^�x�'��N ���V[Ҽ߹qA`U0)���y��)��!�L�W�u�Y4'cr/$��,3�Fʚ�����&��O��<���V`����`�ߨ�[5��O)���N3&n�d�^��=�J&�n��,Mn�ww��a%Mh.6Dg4�)����p�xc��Yj����vb�l8+)/fs�>�im��O��f���K����A�҃���Jl�0AtiB�t�+�����<wYR��Zȡ�%�@�%Z��F�-���`��� ��nx��\��=m�n��jcֺ���,&c��`,�9W�,�]��Lq�H�]�*���&v�����ۢ���_�\�^�pVh~٥�"Ն*'pi
��-H#�s�B[�_��S�5ݦ*ci$�(��aN��&�@c���|�*kޢ�?�����.q����T�w�$�[���e^��^ܓJ�2�"��N��h��dעՌ^r� s�Zz2-��-�������,$�����:({ⰲ5-8�kr`=NT&Ok��_������t�8$4kӉ'�o�/+�.��>WQVh��R��[����]�0�W��â����0 ��A%�8Z�
A��VF;���+�[�-p�8�\/D�S�?;�%��� +�?���:o����˽I'Go�La2��)U����CʴI/-�w+�!����N�e�O:5c�MI������ϟ�]<jݎ�J\������ �@�8-�!��n|��� ��Ʌڝ��'�%R�G���r��SmK�j���H�!='̑*�rc7.ݟA�_�
���J�V�^�0,E������`�Zl2�
w5]~���/�lEf$*ʜ�>�1���U�4���l8�=q�����:���LpksG��o�!�rm<m�Z��~�dRl%�g�Z Z�H5�",	]}AcI{�vGZQ;Y�(�Cx0����*7v!�(fփ��R�m�pq�l�C��~k2�B�0��3���#��g�@�]`��9Q#��� �L��|�."ei�P�o����Tj�2؝(���2s<��#.A���N"��&��R���dz"���)�����xS�����o�55Y�e�Z��J(�� [&�&�z�����j�{}���Z���2��-�S��Q��=!���k0@<��lk
9�G3,�T���M��15��g��O/��x�8��1��-�d&� Z�1�J� ���J]�3��}��a�T���|��|'�����	{��1�0��=�/�l҇�h
�V&��hfT�a!@�����C@*c�[�'������q�f���(tOg�;B$�p�Wm;��Xr���f	�]F ���=$}��ϩ�cΛ�`�qP��g;�tm���U���f�k�V<:�:�oiI�2�0-���FXt� �0R�u��@}%'�'�,� =��If
7��W��7������ҶӋ�o����6�V���ԫ��y&Ll�#�`���}�� �z���;�Ń��c��b2�xgg��L��㋣���7N�MCʌ��������Zi=��jѽ�ip��׻��LMѻ��sgn�d�J#}4k���O��a	XB���lK�����m�8�-�^�=��*V|���Sؕ �g�
��C�0��&�g��B�Iz�enOq	x9;�q�Q+�^0��K��Eܥ�'x�]M�Eוz|��Ah4{hȣqwZ]������!4L�XՍz�h�Y��:��o��q��5�a�"Y�Y#f��}���(x9���	P���	�f˹�2�^��O��L+�a�I��A��C ?*0��|�L��������&"6��ϧ�:"�w��}ʅ���tLE���U�[���*2��[��uP�� ���+iƕD�㶮r
F�3b�W;�j|�Nz�y�� �6�^ٰ����f�d��Y0_r��BN�Q�M{f��Z��j\}z����jX$������x"˗�8���L�����uV��+�L���4��Ӆ�ݣ��{��5��q[�p�GWȈߺ��g|觫@Cc�j�AD�r���t�/�v���B��/�ˆ8L)��P`-�o{_�7�µf�Ń�Vp�I&��l���m�-�ňi�9I��Ï���D�7��@q�V��K��q{��ؓc�*��"0R�4���6�S��gV�hK�zK���'J�($Q�[���a�$Z��Z�|@��w�1����nc��J=	����K�ւ#3�JL=�%�0�j�v� ���w���w
u�}��#s��T>��	ͭ��e�f��*{� p�1k&e}��ٳ��5�)�������G������a�U3�w��K/���0�67@�od�kO�H�B��Gɚ��i�c7��,U�<�(B��.��h��lan �d�䁮�xx\��DS@�;G�����9F8�ߡh.vmB�k%LꀟL�V�OĔ�+z\u��j���A��&. ��@�̴������H`(�
�sϞ<�LG��9�%���3���I�'�sť�	�=����܁�m�Vx6����<��V׻D�x��N�j6cu����gb;.�Uw��7���B�J����̖@�{(�h����K���ms_b͂t�ں�h$V�.6���DN��x8ͨ��x�2�v
�_��Sy<>�~�ݼ��`ۺ��蚹v����݂PR��t�꼣���l��z_6_��U\#</곎���+'K\�x�;0i�9;����pB�iU�]��q���n��Q<H�[0y,�M�}�[+����;��>�6�1�L�4�����jܰ�G���!P��9�.�?ѭ� ����9�-3��j��-qp�ͅOy*�4
��5y���/��B}'.<���h*~p&�d�oj��b�7�i���m.��P6@���IB"*�W�u#��$����5U"�)vMf�̰l>�����aqv$/[_hBX�75ѩ�Nj���W�#�zS��rbLhD)d�'�fQ.6�>[���VA��W:u^������ն��/�F���}�|KD$죻j����̑��>��
;������J��KYǻ��\� �?�Xy��G����*v��|��4�Mj��E�v��G�2LD%a`�RZ&�b�� ��'��B�J�ț1wنyr���b���6�$��@w/����a_��ϞI�Խ�4�@KhyMa)�%69?0^X�#LH�������!�f��q0um[�+�'UDv-��Z�_oy��VK}�7i�� ��?��ߪpo��k<$���tרI�НꂡΪ�$=�Q�;���3޼��h���8�R�"�x����Qsys�f�ΟK�:g����	É���Ẁ&�A =�#�3}�?Z�����	+��S��A�1Ou�[>~�M�����~\�	G
�~oOT����~5��[�KO۳Ȅ�$�U��qg���d���j߼��qɒ�1��T�@Ϟ�Z
O7hl�/�5�N��.��(c]a�M'mJ,=wC8�TA��b�)��"q�=�D��^"��'���'I������`6�O�$q�R)ۄ��L5M/FQa�bHy'��֡���j�����T퍤��!�����@�����ȶ��Y�a�u�I���ך-�/P�_T���4eԱṄ��I!u|��$W�U��en
*`;Ý����r�����0�D,�f홅KK���3f�'Ϗ;�a=n��P���(f�A��l�)\��@FW3��迈,A�4�a6���t��	��Z��J	��w�y����1C�0TRͩ6�|xT�F8����=b�)c��r2�°@͹��u𳹚!ى�*OLZ���EY	�XɴH | Py?��CP	�	I�ݒZ���D�{	\�p�=eb#r��W_ {�eca���i����i��Q����{�Mza�Y�~6�K)2KX%*پ&�� %� [�s���ə���_)�\���i��k�F����EJI�L��T2�a:�\-;C^��W}[:��Ȟ���9?l��~C&��H7�o��55��p�S`{�+�O�W��d��|���"�,� 9�����J�Ę�����3���K֩7*�-���� #�'� Fa�>�w8PuՔ`n�������3P�cӯ�2u޿���z��,̿�ヨ�n�i<�I��2ߑ6�[�ޓf]j��������&��%,�_���Z�/5#���M��|������um�ܝgtJ�7��^E#5`��`'Y�ىS���I�x@�5�V5GvF��~�WXL'G8ٙu{+R�E.�=����)���G��$�o~���M6���I����#lrP�M���Va��{�D�֢4V�T�M�>��Æ��(���G4I�MF6e�
 �Z���%�qޟ ��v��=ٳ�0�:��·�P5�pZ����C��οq���4��r��-��_�h��!��>ӛ�u�z��`kPOi�D�87��N:�={��I
:�5����z�>��2��z��p�δ���#�A�Ob��tz���τ�N�6��_��)�H���A���ө2��a�G|��L>�/�񓶬
����R#&����IJ�!<�5,ZW��M���>�	�K�w���.��߄%T`��Ό����Ӷ�k��-� a� ���h��Ĥ8�k���Y����R�>��\�!�� ��y��>���CQξYP&y�3���P�Zk'\������Hw&j�'��uV��O��\�!�mp�b����%�y���H'���2?��P͌k�Րi,E���5P��[��n5��@.����8-�1?�_h��ć_!HC�6k8Ń��HS:�$���{:�o�	���镘ba(7�?I���M�L���TүW�̡��=���|�y���~���v`���sq3�6��vN#�����d�����u���D�D��`�2��묖V�	[�
�ܔn������{w}�u��U@����g.럁�B�"uKH�qh�>ܧU*8lY���&��+���NO��gD��!�߶�aZH@���*nt7����=�6��T�g�E�G$K6��'ebftZ� cY|�#�_z����)�8o_un7��v���Sa��}L��\�H+��`��$�v�,��e�,��G�}{�c�ą�n��1������"��M�*qE-���2f�����y�df��ՈN넴 �w��h�w��)����>+`�n�z9�����?Tc�9������^���G���Pa�:�-̋���?*�h%��k��9�ct��/�G�/=h�Uٵ⦭��;�4�7��ﵬ/EJ��8m.f����c?�Rq�X�yl��Ƹ�g2�p`������ډ��|�q�J���6��9�����S�(�~\Hj&�-���V�S��$� H-.�w���J������@�hz@jt���lT��|}��� �1T��.���%%ժJ��
TRMs�/c��g�.�;�Y�'cvD�ol���~O���
���e}�^���a²)+������ѫ��&V���#ũNG|�@&Ů"�h�������yu�E_2X>� Թk3DN(�Iͳt��}m���1�;�Na\ �hg�au�	�F��+�Ԅ��bJ�?���dmGu�'~n
	c�a�� �?ɔŌ�§��][��Y;�!h�����m�[?�r>7����֦��v=���F�j�qw�m��ΏvbI�wk�YU��r���]EK+2���\��rơ���1�d*�/��X�Ȑ����#P)6�o�oݛ�q���A�("]R�Qֵ��fa�|+���~��)��t��*c�2.Q3R��c2º�X���ˇ���ѓ�����Ɛ���%wo�Aƪ���	��������w�J͵�*P��N[�ݲ��Ά�N}U`�عl� �
���0W� j�qBk���
:z��L�V�歸��ހWP�Ұ�
3�EYP��#�C�KzA�<dl�n�V��&�k96�����d�� �Z)v	��`��|Nx�abC��_i���B������_E�O}^�\�&��,G���z�A��"�L*q#bLq�ߴ�g��W���iN9����r7�eQZiI|;O�ŏ2��*��Q�4ҟw��y�;4�x��p�F���/���c��f���Sd�H�8
���n�Ӫp��x/���ķ��K'4��g+��L�'����u�Ȃ��c��B�u�kM�-�c:�cRP�Kgy1#TG����l�X%(��" �T��ae�c@���)p=��L�8n�eOU�5�G�Y�P�~���e��i�{7=QQ,��>ԟ��:o3��HAPԳ�� 3���,�0� Dȓ��v֚B ��$��r¨�c�Z�6�^F�c���#xX��.�7ʋ6E��n|+��n���J�J�kA�G3vS��U�=~h��)���<��o�'���6,
\T���l^a͑c�[F�@I#��K��S��*�O@O�\qs�|-o� ��Y�}6��1����7�U�7�?w�����R��$��^c�X�j��s淌����F��h����)o���S�S�p�Po�'��RU0M׈�1Pi����Q�e�#�~yϒ���A��%�8�Xz�]�K�wm����)(J3�{�"���S��AQ�{@���p��W�S�|-�"g��y�Dę��N/C�J������ǏD�X��f���C3�'��f����vQ]��+��M�G�+�jx	��i�w��>�،�4����0�W�)�1��]<��d����z����Wƻt8��J�9f��Koq�����D�
d<�ؔ��l�Uh��r<�A���rL�:�)@>�v$�����!�Ø:M�9H��UGV@%�鴻����Ak4��Ʉ��9],n�}��p��j����k#(��!|E&yO?(���ҏ�t�@ >�V6b�%����A�f3����s95*A�����mV>�4�&�joG�5�
�@�� ���'yg�_gY��D� G�|ʜz��	���D�T�T�E&U�*_q��R�0����Q�N�>J�RSEaᦵ��$L�k�$t��j(FӔy���<�B=�zX�����Z��<){�ou3�Iݙ��Y�A<s�Ρ��H�=f&��c���]�S����/t��&�KY�;vb�]L�s�4��$��}T�Vyg��eu8���%b�|�7��r�^�"F����ܤ�zxH�7<6+����#Q��M���䫂���2�����-�ҵxE`=�̣� =迆���qÁ�l߹o*��*[f�{�����4��=(�=k�
�����R1�E�����9�@V7[����)�O���B�[�x���V� ���B���X:a+�%�Zk��m��I&ŋnY�IY*����Z�=���heH�4�̯�5�?ެ4r!3/T�������wsZBh0�d���Y���-��Z,�'c�Sg��e�������Y�:�[+P���'sw̵����K}`~�����!u��7	�>��7	6������f���)dD����/_*Y� U�S��mx��T��lT�#]��ڑJKNpt�,�UMP�T��K�����Χ���̙Q �+iq��e֭��R�޾�A:v&,S�#!*{��y-i�Jv�y}��qz��ž.=[+G�]���ݓ3ν�0C`�n�Mv>�B6��z��:!�]t��/U���U���8�J����TU�"䖸�
��f�g-؜�~g�������Y�sg��g���t�ʷM�i��+�3� iv�$K�l�b?@J��V��E>�}]#!�Oy8�u-����9(�||�Rݰ�>�u˛���k]]o�)�ul<
�}7hU1<d�b�t��(��3u^wy��o�2�E���	�䑀��R��q�!��ʨ}��y¹�q�#�O:ޡ��2&"d�s"^�3�����e{=�=l�����VX�蟅v<���������"�b�Ju�`s���`�!d�z��!�mH	��j�:U�1��|����Ѐ	N(�5���S)��_�����#�0�~lz�3�
R�Os�_Z��FH�	�0���х���`���˾�e����{�����Y���Q<��l�`����֌�<DGo��YՕ�a��]��fh��]��݋�K�o�pډ��޷F�,�l�&&t��R������#h�Z�{�'�YB����_����L#�*�Q� �{�b��tP`W_����q���1n���l ��L|k����\I�p�ǵ�+K����:C���˭H̨d[�pȜ�d.
��%,������nÚ�I���v���a6*s��#�-0����PL�q�+�S��oX��W���I�j�y�MV�P	T�h�A]�&J��!鍲�^�����O-�����.�2�XI�T���B��H�/ʋxZj��{aKӕ��F����xY�~����J�cE�����{������J�&������ O���"�|k�m�*r>�{��;	dTQ8�@�t����s�	ŻP=�^����ynԴ�����	�^߁�=kA~�p�{@%��4�^���s��Q�=.J��%��8UC޽\�)���S��=.�0ܗ��O��f�.ǈ[e1��L��`.-�#[�ϐ����R?����X-?]�t���4y��Az��7�✉��b��N8��g�kKG=�u�����gspt�g�\g8��EIx!�ղU��Af��N�,�P�"+��8�X�{��r ��4����?d�ԶU�ˡn�����k8&VW>FV:ly����70��-7�9���Ug�>��xw�&��J�Ӣ�19��5�CV��E�I���
�9�#z��B-m^q��	�?�+Ϩ�ob���U�Ԙ�A�}�S7�d�ik��'0�@��������6e��_�c�E�_2�f$����A2N�\}_"�4�	��}%�7�6(�� ·�J<�7�0���J!g�*|��&/���8&�����67�C�}�f�_�"xI�2�P�jH�M���3.	���E&Hɏƅ���Dx�����q��%Ob�L��N��̢������Ӄ'o{5tub�kEy~����-���NۿC�C� �v��׿� ?��=r���j�
�"�C�������h.��s����?��eB����3"� 
=f��"�@OF� �6�]�N}o�1��Ms�v��MzMS��l$"h���qvzU� �.�|,�<���;���#���aA��z�R�cg:�8�3�<+��/�n��-1	�fWI�f�<��4uj�Ej�6ET��w2S�T,�П���E��`����ރ�:��tS8��z��<&5���� ������l��x֩��@:&�����P��	��%�FM�6�7H�/�K&a�aO�lbz̤P��'�~�G���r%n����g��e.�k����E^���2��(�������:mGD��!m�2������<.~�*4[h�{}\}c@��� ���`q:K�fW��k�U@�|�>��|�"N�6�-�L9&���)U�$0�L��u8Oy��'���"�)�!�VGU��JՑ�~��PDR!��p�d�A�������i\5��.u�mO4JnB*�ZƆ^���^x�>o3jd�szs�6D�w>��ܿN?v�`���Ǌ�}@I���~KC�8�<~%���qm�h��h� :^�#�eF`'�f���v����7磨�-@���^w\�����q$��u���Zo��ZHXC�՝��+|!Aog8�̗�r��>IA��Ǹ�f��d�B7zvG�ڙ<�m�קV�=�-I,��e%�!�5�0�D����9i������Soe#���+�)��,���D�s��f`��j7Ɲ�<���D�o�#V��X���'Y��V:\�{�#�[�t�i�pi�eʸ�ݱ��p�BJ�C��*π=_��B��~X�
����4�U��H�qE��'	����Y:�_У���%�_}��'�p5BX�r�o�Ȭ0�ȳ_,����4f�r%�zSF�(2^�Vpޕ)�ȵ��ho���BG&��%�����kb�bN���v�����G�Q����h�_�`�:(�A�N��|*�Zf�����jyg��;R� �$#�]g��C����	s��KA<ŘM��;ao��җ�dw��,iՊL8b�\�P�豴'Ut�sn��-K��\�;,�����P�λ�0 �.�����qZ�t�7�A��	�]����T�bTl7�8�a0��:yq�2O�"��{ؾm2Yb��'�v>��^���o.�?�^�||m���&oz��	��~���ߴ"�&Ԁ���,�D7՜ �\'j��6g�י�e� _��0H�v�fc:��VN�!R� Ix��]��Yu���{�橫-��\^X��0IU�g2�8KȖ��>�E�6Z�`"P3^���[wI����1�+���� �n�v�4�}����BǋO�7
hK�����ϑp���z��W����M��wWX:���q���wb6��;��m63H��;�*I��ً9�����*{_��呮�D�����\�5G�Z�?F���=���V-w�j���U��Q���3(�w	��}�f@*Ħ1��\�~�������le>oH&�;~��ҍ6~�p"�a�S��E������@B�/0p�ԛcԗ�]��|HE4���^�DER�fR�w2+B%�i=�����J�y��7h�����y1|OS����Iľ�oge�O�q�cS�}u�q���aD�*E}�-��0C��_t�n� \�,�zP^�����-��0B��&�.��œAwz�!J$M#y�8�I:����v�խfg�g�P�����ze�n]!����=|���<N��Nq;!�J������2X@��3uP�~:��+����p�KIA�3VU.�ߟ���H�Pw�ַ���_f�
:3D�$�b�9��#�o�� A!{��O�������9��#��҂��H�2�(�;���Y��Q�N��~�������1I���ס����oޅB�����Ddn�SȰa��0(�� �Ƅ���i�Ϭ��6�2���C	�XL�L��o�{Q��(8�/�n.���F��e��o�>[Y�@� +�(��N��d2��#L�?� ��&�pZ�;W�x��Z��3�ϑB��3K@ia�s=���_-X�������F}绶���ĉ �� h��8�[��g8"�A{E$p�.O����U4�3��r05������W�cn:c�cx@�h!�+;o��8%�$�� :&�N(��C�+OB3<����c���4�*A�+��V)���l�Lb��b��v��vc��3�� Zn	m�<E�/�b?] ���}?��դ�B"�{��#	��N���x�. �Y��X� \t,��i���@��A��%��S?�����h�Ua^Ѻ��*��(ފ	��D��F���s<��4�'��!:�q��e�6���jD�+SH�ݧ�jU�H𭃘���Z���Wz@{���F j�[xR@�lAS�LO��ٓ�V ���9y�HZ-�߼���HEu?>�a��X
���H@,M��5����5�%��a��8��lL�S|Q�{���a�;�'�47 �"3(e��5 l�'N�L�=�q׏��'�u���,�Q7>�&���wu��T��v]�LzQ��|;�W�ka܇�>���d�!������Cѳ��"��Bu���L+~��.�t��J�Xc���iQ�r��{Y�.�����a�'�@�������z��n9g5W��I}�f���g�|z�����Йs���?�ldJc(��3O�5����CӒ>a����jGP�B?������5�<�RVGc�����n?�_���h_�?�����!|u���;f�%3�`I�S� ^u��5�hجϒ�����=��&S=KB��8��wd	��K��!Ҟ�Z���/�>Z�E��y���P,�QJx3��.w��A"`gg���j�0!*P�!���vYA���+cg�����2�w��Ӹ���u�`�-���g�!BO��#�t4�!��¢o0�m�J�+Vҙ�I� B�.D�t����w��;��
��24(fZ�iD�y�\E����\��8�Z=�;v0��~���,���t����?�����f���L�-�_l��x�������u��Ϯ���{#y&���':v���y Q�4Q��g�l��j���%�����D��)Co�S�˅��]�Ł���=aԼ�Wа%��*�s�Y�+$�TYw�Bݝ��l��M���&��a�S�g2Sk��9^�8�N��'9�T����J����S�6~zX��	e#�$Ք�g#�a�
�n W�.����������29⍛dܞ;����aq8��$�bN��cWz�0\ ��e����gM�`T���ho�/Ic�&���7�h���	$��.n�L�G��S9�MĒZ�r/XT�E�W�xx)�.Y�A級�!y _����͌��U�C�i�.���R��c�bLj&�h��O)���"��F������+͟%H1G�w>dҌ�Ғ�
+2�9w�-�_��H�����ĩ?�H��:w�ݕ3~��{c��,^(�c~���?'y�����q;VI�sM"�z}�ɺx	�w_�
#��I�$S��L�>Å��&T6o/^�w�R�q$~T�< ����EjN�7
��M��B9�ֲ�Dϧ�ܐa�к@\ٕ�4�9/=Π��'T��f	�k�J_Nc�?z!e�<�Oԥ����D�v�����ݻڭ��D #�gT�E���}����K�Q�=������y�)� ^V��1G�(k�R-`(vꛤ�AF�~,�h �_ `$|7�	=����-?]�F��*{�q�&���!��}K-^��|/:�D�^V���7�M��hw��@Y'38�G���� ��Xp��G��� #o=Y���}�\~We$l�!l`EeX���9[S��z�A�r�N� _����Ze]>�>�7��\X�8�e�`���ı(�#(��1n�����E^,q&|�<��M\�0�X��!�2<z0]�XMP�K������x�avU�ep��WK�Pt]��o��P����$=-UU �&������DG�-f�o�I���3�q����O�����5�0��a �ί�--����n��,<m�|ܔ��P��_���=�aM�DR�4�{�]]q[�eb�u��g�����C��C�j)��ظ�C������Mbp7�G�L�6�7�����rw�����oe�If ����B�3;�L?��ֻ5�*�L(>�M������d����)_G����r"ҫ�߀>n�&C��cS���͐k4��i�<I�!{ZV��2S)�����k^�\&�Q� ����'���o�Dw���=���igj�5�������ߋ�IфUo8�2 �iqe���_ ?�ѯF�I��h�8�q1�����J�ZI�'�MO/��ZP����c�T�Y�ꇵjSSv�Wʔzd�PY`x#�>�(���߈k�	w*��Q�����w~_���>��v�`�h�gv������hS��	��#��6��!���T�Q���6wW�\�fEFR�x�u /�7��w���ȫ	�"��Q23��_!:#&Q�N��ߣ�۶��'c<�S���kq :�QT��gȌ�4�8w�э�
�������\F՞���,�E���tq�?}�q(e/qk�e��Hk���VV�XO}��W/M��/�r�8�i��+��Y�p"黫�!���8k%�ǁ�^�r���L֫��?B�k��"GI��sL��*l�Z�v�TgL��qb5����rf�X�{�u� xe���40@�Ipi���R�ծ4���*T�C�ѾU����J�۲z�ч�.�.O��U�+*��	݉�՟�Bl;��	-$-��{�׭�3v($X:��7@"�%�]9ʄ�c)��V+����kE��)����dQ��d�{�r)����]6	&nׅ��Vӵp6b�*�Xch�W�Q?�Ĕ�-��&3�7���ǵ#��U�D�7Aݎx,�l�i�YS2�!��!��2�BE�!��yYWktL9�?�y�)Q�芡����o�j����<1\l5n/��X�H���CO���nE_�dh��B.
9,N�\�//�zR���t=ߢ�ID\}�db�Q��Z�ڹ�v�*g���E��,z���;�JԲ��j/$Oв���y��R�FV]�jk�
lQ� ��tEkM��^�i�3�H��-��R��)P^�k8�[O(�d�"�J��Z$��)�l�y:D�p���c�r	H}�}� �q����|N�!�Q����-�4���g�R4�$��<UMӘ�J�v`c��S��A����kR��쵑�`-��	r����ұ*��"���}�AR���SOhq�`�+���]7�V��\-��+�C݃���4i��r���aqe4�p�K��G;D:m�l��W�b��ź>�� H��l*�͟5B��K�5L�!ۥ@��14C�����(9��?a=���3U�s�PfS��n�A���Y�� f ��� ��GM��Oθ p-��,���5P���[�l?��+�R�D�t�:Zģ
�&W1&yO�J�fV��YN��̻�����d�D�$>��LZޙ��r��F�p�'���,DY�T �p�l��(�
�W���U�:����$���1�mj6�@[�&68��ԩu�i������5�Ϗ��I����y��*��Z��PӁT�ۊ�_L��"zoO�u!@f����wҲ��o��nb��a��I��H�����}ø(���[5"���g6�N��-���?����tx���*U���0�j�I����Z���@�1���Д3�¤MN,y�o�9��'�$�E$��V��İ��}JGܚMc���ƀHT�W�	�����*ڶ](����a:v�q�..
H�?H��˛��%��Pz����]T�SER�y�E�L�	����tp������}p0}��'�#���AZ0ؤi�jQ5��&�i~�o�A�%��X�p���7�N�t���m�^?���ޏtfw���
!^�N�[��Tp��bz��|�%B+s,�<�Sd�5�������o��Jq]�QeW�Ր`����/ i��_��8yk�	�1!1�
���JF����-q=@}H��ͦ�h�s:j�+ÉW��qJi��n�u2�����OS}lg�K�#.��q4OZC0���3�iT�\wVC@c�@O=��h����Y����\
��g��H��]�DS�g��/�0v�P��фȻ�/O-�?r
%�����\J��{P|M�������<5�b����E��HzB��Q&9��-&���n����X�M��}��p���M�~�T�T����<"ԌX�#��*�B��Nl���=�¾�;�nGrY;�_�An$�p�$�f�8G��VE��G8�^��Ad�K$�����ǣj"��������J� U`���B��h��G�����/y����$u����N�[��M«�%Z~�W��9��_g�'��8&et��ELWf��������A��/ϖ
��o�5[���<mh
�����v	�(-�
���:�q�{�\
Yx�}*�_j	(��=`�UnX����]����>�^Y�w�$(�b�m���b�Ytl�GK���L��O̰��h�0,�]Ór�iv��%�唆]N)#�{P>~I��)_D��h-M�"��L��Jȥ�-�3�M�Ȅ���y-'�����B�͗���#1�B���󩅾LK��;r�E�K��D띕1��٘�@���F-��;�6]�Д��)���$�-mEI�9�������%���u�ˍ�O|v���,zZh���75��w��{��(q$�þ���z�R����	�X�Xn ���͡3B��	�\9,��a0i֐�^�)$T�oknT.d25���V�IQU�Z��G��d���d3�����}\�*���ψ1������L�\pO���h�n@�cK�C}{0�eN!��X6�Bƞ=ܢKa+x�GN�w�,K���c�ƀy���t�[}(���A�Ƴ�*�<��;��t~�T�m�O���� 
��P�_�&�Q{�+I���5ךWP*��� ]��	��@��i��"�~�T,}ۂ��|a�UĚ\_k���U-TCݥ��d��x=��V��܆�K���M��.���X�ǳ��/�:p�#b�JU9�Lt�!4�CWd�ߣ`�`�'����d?�(�;��5�d�H%���z��ʇ�]�nk�#LqK�\���٭E�i8��$����i��u�^_��f���^�к8��}Q�l���ym(hoc������b��Ь	X#F�%�����J�?X,���BKs�
�_��*�@�@���|�ߜ,��UarR>��ZAmn~�����~��Eڅ������!�آ�W�N�Y�? �S����Zb��sn�RN�tUƤ��c<˫�S�֝����7
D��4,k�-;&�
��Q�8Gŀ6�(@�}e'[����e�%�>Ո��(vf[L_���1r枤,d���
�P�L�(}���q2o��-�&�ġ�kP��mGn)�m��`������3�j�+��4?�O$S�G�j3a�{�����`��g���9�P�r xr��;I!�����,}Yr��o^Zu�wr��@�M��ۗ�f�z��Le�a}�`��f{������?d�zP������/�Z�S��o_7��A�d��*U��x՝�,c?;�2s�6���gz��.EՔ�U��a��`w��^����H����z"Ƅu���9~��ր��T�q�y�:��<k0�U0���j�����"���9�jb}��{���ѷ���A㛻 T��w�۪:�=T���G�>-� �����OP�kxv�\�f�w͚lT� �X�T<L.)�/X�*t慝 ?%IL9ZZqy;�0���7��V��G�,V^M�5fx��p����׷΍�y����j��6�/�R+�HP;?(�G���U	�1���7�k�EjEJ�w��Ֆ.�uR�am�����S�C2,]�1�����^a˶�Pp�K��>�C^T����x}�<�7�,< Q��~����Aήw:h�x?!���PV;s�n�������;��ebɺ�,f�6키W�n��YT�~�>���

a"+9Ҿ��G�~�=\�N�%<lEF��g�2��|�"_L{�`So�C���.T5�I�f���g4bTQR�z*�N�w"c��ٛδ#K���>��ao.w&7<<'��Fy�L�l��j�s��O���	�_i�nwe��[be��Ӻ�<�s[�Xd��Ӂ���7Jvc��T�<=P��N� A!1H�U<B�_�M����B�(��}���M@&{&����Icz���X	��$�򴃍4���C�H�ꮺ�(���x�`����E�k�ƟapAA��^������{�i=����:0fN��gca�ס��r��g�ڢ
%7��x�;��+�|�@�ؓvpWk���}��U���=��K��-�N	* ����i���s�$.�HWҪ�*�B'@���}�4��N��Nb�=L��T��+���@.륹�����.�����%����i�����c�P�'X�`�ӫ����@,�,?G�'����.i�����,��v
����#�?�.y��L0�����?W�1�� �{��	�k/�%Ս"��m�D�mB�6�[���h3���NM۪�g&�"g�/ek���D���$7A*�%u���/ԍ�37.rVI�� �-�������S���Gf�9܆��� nX��ɖe����]��ɾ�͏��%齔�j�Y<!B_�]:}�"X��_�!V �8ƛe��E��+dʡ��3�26�o�G�<�;d��K/Z�̠V�k�����	�h`�]�1�-+π69xӡ� Pi��ؼ�(�+*��|��s�"盞>��%��^g��A��/I&��B�/�{W."��&U������iAD�)���L��8NT�@W��*#s�<�aS���G}��Y�t�*���՜vJ�θn��4<�6�F����f�Ċ��d(x��l�-	
\����������3H�t�~���F� J�mջ�J�������h�-8˲��á���`�>��ED>�|������o�u� ��G58�o��?�`_<�u���&�+������=�6�.R��Ϫ��ߵ]��nH��Pm}'Z��Y|�l�n��9eh��N���V�ӹ��%�����BU�`}��
 �A��h8���ռ]�!�&��~˥���c>�\�X��x����;@�=�`�YyX�		�p���,�v\�o �L:�ihl��s۱4�ј�g>�B.�A��'
n�-��4��\�
�"�(e4:��Ҝ%�R��B��I?�� �C��I0�|�w�YS��?��%�A]K�d�K%^u�ke:�;H7���lb%��6k��š`G���prVt�
�npQ<�p�Y�4AlM��
���fZ姒+u��N�
ʘ���HĻq������2�7�ů�#�`Q�5}�^5򿂥�=��i����X��+k)������vɈ�r��,�2ܵ�[��
��T�@��K��}/�����GRxbߞ�~���p�*�(F�]�삿�ɐ�r�mvuJ���}>��Ȟ�e�[+W�p�M��J|�@�JrM4�L�y��y��+-b�XY�t�� zo������L�\��6�����:Ջ�g��Vc.}$|̇����S؆-��߉U�����`	�C��X���I�Xv�uH����1��m|�Q2pm���B�]l�J*dQɻ�le�@=��F�om���S6w�(�W�y5���'$[mL��bX|$�դ�i���ب�H��f��-�4�ߥ�d4�� ��mM��E�\R�ѭ���Ca�艟��^���z<`�q7���X%�Ϙ������Y�_�)i` �݀�miZN��RΦq�����D���W��z��Ą�7̔@�����  ��G6�.,V�;K.q3�N&u�Y6'%^��'��߷~RL���̸���*7/��<�Um�g� b�e��z��+�VM���׉6�Nx��bt-�Yw��ᰳ��{ ��A����d=�i��^�����]�����G	\:~C�g�^t�Er��������b�̂J˙���x�4��L0B%J^�O1�d�=�_m�����B��i�%���q��*,�MV��Ga��࠭����xu�O^ʀ{5d�2?�)�c0��-t�ړ��IO�l�6f`Խڤɖ�L_�ӬDxfi.ߑ$���g��Ʉn���*���\jd!O�M��/l���3��?�=�I��0��x�
E:)'����R���<2	o�Ҫ=�`_3�/�;������@sM�F���Ϋo��t�f:.Ԭ6kN��$e�z^��	kv�у|=�}�z���,3��`��Bǿ��a�g"����m�Fx��0���
���S��|e�T#����:*����|=�h�o�YpPJ��#�"�$�|�L4G-�IZu�Mws''��}m�r��dh�����_�yO*Z���j&���1�hw齄|�eソ����Z�'6ۄP�Gk���D���<�m�>�y�\f�L�YK����wh�K�����'�.Bل��FE%��H[�&,�}�J�q)��~:�?� � \߽���ED	 \�Au"�G]U�$��;fg˱���e�x���Fw��
�|2��:D��=Zd���	��J��{��)�/z~�޴�ō2���l�(
3����q��B���9;(K�G�_��T�(Qh��ڗ��xJ�Pm�H5D|	sx%�&4�����Gmx5�wjzSq���2љ���� {�^�-��#8z��s"u(J8;y�����*ݑ��529!H~}�z��i��@�%z��c�I�#���{��R�M-�C66��W&J)�#�C$V��e�{�4@`Si��)=���<��pu��C��E�"���~aW@���:1�'��8�jYi�k�-�BZfs�T7QӖ�n��I�JF"/
�/Ѵ��g0i�� �]E�_�w��6i�U��<	{v��O��+Yӹ�_E���Gl�>c�Iʁ������R�{&���}0��<ynS�=�R$Ȧ5+��Wz}Y�km~��oC���!�km�����������S���#�BF �R{	����/�P�4�^�PC� ����y�M�R�1"/�,/��'=�F�X <�E�<ĺ�	����h9��;��-�^��ü=�l+֍���
'��x�T�c��V��Y5�2������:h�8v��<q,�ք���k�1���oeTU�fL��3ަ���Rc��)��(tu�����_��w��b��j�Rܥ�u�Vu{ߦJ��O���+RQxx��e4 �b�"4� �-d������ָz��<�!��G�U�b�\�ȱ�+l*���6�bK�L�ϔ�f��.7S ���zx��N���b�7�����b���{i��޺zC�� p*��DE���KPA��J9R<�x��ƚq�^�ǒ��l�##�Q���*)���B�v�t����iA� ���^���ly�&�7>Ng�������7���f]�Z3d�����r���aL	���pG��Z�g��}����+(Z��5zyu���<����|`�����������3���I�X�D�LG]U��^vx�+&���B�۲�%�[����k]W4��F�Rz)T��p��[�B~F����z�N��)�b�fD�#� +`�5�#����WD�U-�2�	�~27��Q�Bw�6�-r��S��0&F��K#t�1�"(��*0<�æ����}�"���E�ڡdL�L�n�*%����^����sX��U&6��& �ƅP���y-c3�f��'$�ܦ��O1�EJ��l4(o!��u%"�<;���
��l�a�f���s�������4�����V� ���c�f�V�G��=�b�����=��B.<A������aB_
;ﰯ�E"�m,�G�6O��;䱁$�Y3�U**_D4���KمG���ix�5�����&s�����(��Ւ�`:�����'��#�t#��T�Pr�P��-�jaY��
��|���
�p�˛7	v�,��X|q����L>+u�ާ6�$�|��������87���߅�j�۳l`:E�z��*�[�$g�Σ��Iy�KfDDtr@3J���h�;.�;�)����[�1q͕~�N��1x.c �2m�&�x&�Z5�7`�R.�*�M�m���j��ýu
���0�s;��6��W/��~��i$;x����*�(,(p�I�}枀��`�cE�����v@͔�{�1/o��� ��dP�c�1.���ET<��k���
J�5��D���fM����1�;o���˅�E����
�^��r�E�8S��:����o���$�A��M�Z�o�X��5O�lş���� ��6KR���$%Gm��#-����cc��[�����֯���2�Z�y���;��Z�j���{]�%J�t����
�T[ ��H�B�6�Lɹ�����)��p��P���l|����\$�7���TF��༰2���>��O rӚ(.��~�gi�ş45՛����K�'���1�k}gRmdv_�8���6�� }sDhM��KET��E�����c�.��O�qտj�E�q�����h- ��wY�.I0��q:���U�6!���\�&�`>p7:ٱ�!������a@方=�t
��?�L��P��gj	�
�6�걫��):�I�������f�N4X� �9�
�>�N�!|>���\w��6���CV�#$pM�������EPq O���G c��qP�R��pl�# ��~�0N�d���7��5�Q�E�wxFa5��_0���q�$�/�
�
��~�#;"^A�5*v�����ST�q�P�:?��ߪ ��$0����e��}/�G�`J�����<Y��<����+���ϖ�r+J�鍛��=�~�|`�'"t��U���z���q@��ݓn�h�~�[[���*IV	��p���w�Ndl�*�mY�Q�TLAЁ��>��bs^!���Բ�c���CF<�6K(*�ۢ��G�ҙ�˨��_�Rz�ؽ:��uF��g���<��{�9V�u��eo�I��J��}�C'3�M���q^-�d�x�� �a,ߋ���2�~6y��U�q�οj���tFD�[��Mmݽ�I|ߩ[�i0[���F_gg����d۠a87�8\�u_�:ɀj��ڱ.�T@:ؤi�4��(>�A�Y"����{�׵���l��J���/��2q����p�I��;��O�+�ׅMJk�A������k3T�1�-T��+u$�xzaԔiy��{�FЌ-�h�ӥSZ�@(��ys8�3.�1H�6���$��R9�i�xQ�S^�Qq�vLF�MO���;�R�G��}�g���s!��
�"��D﫛/���qB�Q�I�ϻ��C�+L��"r���Lj�h�1m�_VS�w ��f��M.�ռ��[T��bJ�/�c-�� {�/M\��s�x!GL'�9��Z�ڜ�nEJ�P<`���u��i!�8n�j<�����-�?#�	�Uh{+[��S9E���?�7��i,��A���?}mC�k�P��K��b�QZ|@8��)6�3&A����J~<=�8�4Θ4�w�o��l�t�ꯊ�t�y��hf}Ok���n�r�<�A����=!��+F�B�a��G�>�����Lj����ҿd�X���f\��ׄ�sQ�{q�i���,��u��[������P��Nj߾O�m�}osh�`�wi�W��o;>N��(�!��-��Q��h���5|N��{�[Q����;�� ������.gq�9��o�*�lA�,�|gW��T�E'Yyڑ,I���D���T��^2S��i�v�)����ɐ�c(!D��&�0h��ڻ�f����i��) �˔�FL�"\;`�Z���	8N��Έ*Xu�f��x�x���W#?�=�lz�}Ye'"�q�uke�=7޻@����ш���A����we]r́|̤[�l���%��X�ϻ���x�	"���8]���T^6F�;�\���x�q�K��x����Pu����爮�Hܼ�g�ԏ��_u6��7��Q�M��rT�����O7r�ļ�Oy���vq"q�mӰW���om��ګ(n���и3��69,�;�w[\x$�	�m!'M�k�HL�M��y�%��}��K�|f\�k��+�6ql8:�*�����)�l���V� ����w��]fql%'I����cԉ���֧�ڰu�ylrO���m��0Wj�Q�if���ta�U�OM�#��l>.Ն��]�Ur~n`����olg
qS���o����4���ܛg�_Tx|�	ϘF"SM@��5�E�&��k�O�<i)0sG�v��K0ek�����K+-�ފ���]��朗	���1dJ=R]Y�5��|�R��EMdf��Gv3��I��W�mO�o;�1�8ө�Jg'��{�6I�XÊ�ů^���XkЫ�qA1������	�"	��h�Ҽc��+y��)��LRYj�����͚����#2]�ŏᐢt��ul��)����@����A��wJ���k���� �%
��d<36�Y6;�3�3U�3�A&!�'���o����΄�YGz��]�A=��R�dq���H�5�f�1��𽏏�t��$Q����w�����)�sr��pe`�J$L`�"�10f��Nց!VnMG
k�z;Y2���#��|�,��j���BYOC����W�lxM1`w���v�e�b���~K/�l���a$}� g���J��
�I�?>+(�N��^¶�}Ҳ#oTt=nM�d���?�!});	�M%4-�l=�3`;'[>�[���'����ϼ���_:�������3)D�~��T�;�oܚ��F�T8M�����O�2��B��K))��QV���'c�3��$	k3CR#cY�]R9�	0<��"�ce. {)���ةn��B�zL�,�Hn���. ��(��O�P\Y�'��c���+�U~,�}\s�=]}�qLf{�@���
o�$\o~�DCfO�Ŗ��(w����`��'.�=�d�ǂ�N�Y�yg={(�1y���y0��ӽ�C�:V��㕵E�(��10#nƈ�l�<�F��a:Щ{?�}�8�����K$�%�-�����gR1����A�����T�`:t���`'��> C�Ev��]��(���I�ϥuܜ�g�����V�k�VW��_yHP���D��Hrd�{�e%	�e]�a��g� ��^�v�N�-@�	����|�g��8 mG{��\<	ie+�F�L�L�TQ�ƄQ#l�Z�$!T(rB�N���	�|�X|Y/��7rb�%�����Ȳ�Q�X��~�5�Mf��G$���7ܪ$ۖ�LY�l�����"��o$�����l"��noM��\f��fJ'O�Hq��.~|:M�1ϕ֍�������2l�)0���̦�*���!�}�u�����#V>I�
4S|,%5"��Fe���W�b�x�F��Y�i���u;` P��05�U$*�;���~������z�>��yk9����\sn��4]pwx;�$s��_�0�6��=?��td��r+��Mk�B�d.�tƲ�ʭ��`�	!V��.ĭx���;�Ƿ9����n�/`�7�z��rVW?O�6|�2�xH�+��斩Fd/W�)�����-��Ah�	��r�i�$�U���%1��i�Y�"�%ɔwN@�N����hf�#���x���Q�d�N�\NfFOJ{l����5er�ଘi���O���1���&ʐ2fo]��I��O���K_��/r�[���	��Ӝ�$���+\l�6��/�7؎��_�0��Ź�tv�T?��P5kŦ�����Ay\���U4N�Κ����X��)�eT�e'�}}]�N�A���X"�s��e�a���M��>����5��zOf22Ѐ��0o�F�����[�PK��_a�M+Ꝛ@Wu|h(����Y�X��^N�?3� ��E��o�����w�D�]��иv���&�P�DS�����_.����Fk�yd����ۇ��-����mW��y0���T�����_���,�F\�1�-V	��3���Fۇ��+S�C
�7��˷+P$E�$?<�Drh s4�P��]�dP�Ä&��"� ��(���<^�k�����7���֌W��]�6�ʔA2aͶ!��1fXL9��C���&Ew��Xu�Ɔ��03oo�)�l��\9������J슙��*yl5=��HB��V}�-8Z��]Y���$�Y9��C�CF�C.����S�A�0/_}R�O����<����?	-�S:t�p��)ٵ��<*���Y%A�]�wS!��KMa��j�8N�wA`�
��D}>��N����1�Q���� �Y���ņv%/�s,K#�à�C�䘏i�-���z�v���$�ȱ)�\qc���W��<6+.{�tZ��J��7�a܃x��?}
sQ{��,D�I����i՗'Ul�QO2uU�B�qc�G���n ��EcCU݈頕��拉c;۱HQ�a��i��@���]ǩ%�����ݜz�v�Ϟ�h+��Oy���(�B�(��`S1T��@�$D�g^�B�(�ΐT�
������1�u�#�f����u��A�ZOR≃�?c"\����$m,_��gu��.�SB�ʊw�=���l���l0p��}A�5ិq[��bngJ�_?j������-�Z��H��U��Jud�7v���XP"-n�nP��׼�@�~B�ug���0ob.�E�=�s�Z�(t�vh��	Q�X�����S#�+���X�=6)3�9�45X9){Y"K�"�*�.�{/D���rn������o�;���9VM���t�N�#������BN-ׁ��]	��v"n��Y\����6]h$��d�^�Gj���Z���h�>��e3dW-�Aj�|r�9�x䂪33v�l�d30���>�7�*���u�:���	��ar�'E�� B$a$g�~ْ�5��/�FO]�3o�ȶu��P��%��$(hN G�s?�g�n�E�B5b, f��
�wI5H�@i��a�?L�;E��O�Tx�e$,2 ��n{�Y��"a-���``������z�k���y�J�}H��@��s@���;�:I`6L�N^�|�1���\%���d�6��EP�>�]��߱� �rH���÷�ʁ��8�
����YX�;)��A���u[S���S`��U���Ya�;�*
VR���>���-�w;�>�Q�j@��w���l��N���+`�[���n�G�(����H0���
#�*{A,�<�՟���lԺ�s��V�`Lʛh�զ�U�-j3�r����C��M{D�Xp����`@b���A7���w�WQ� 'Rq`�;r��N�?��F�y�����DM{��^��SD̵���?f���,g�.�����!����o5�g� l��QK	��]逬@�F�3�o�{����@�FX���Z,.�k�`n.�v=^�8ۓ�cx����UW����ꍧ�_J=�
�];�A�PFE�K�%����ع4����Qxo�qʃ[��2�4Z�U[e�/Px5uًT[)�4{%Z��1Y��� y�{��t7�9�/ٜ����B]���[%  j.u�8/> lPt����,�Ws�H |��4l��d;"3�U�����*9Ea<V�{=�8�Dˉ�u��#&�gw��mT���݄�t
��l�/1�gVO|��)��e�Yr$�N�)}z�܀j��4�O$i"i%��*2R+cwUY+߅X�Ӱu�����۟ ��#��X
�9
@˰"2�]�x	���{��B"�F�����!� "t@!lEc��3#��G�����u�h6!�z-s&#J�.Z�p��>�3�t��F׬wE`�s6�b�h��_
�9Ɲ��\�Ų:
� �Y>}J�#sY}��Wϳʸ$�9/�K|)3�OJs�o�][?�)`�i|&l�D%y�uX�C�js!H!DޔU��[f	�a�I����"�^2W�BH�-�CO�S�+�V�SL�����A����H��9H�\j���.4N9����������{B1�JeG�5uD\[ux
�
L1�0]C���f���E���w���d�����K�9�=�A�"����-wb�),%oh��;��o@̿�i���(�A�>�)��M�.�Y�������6�W"D��5`��~�q���;�k���	:�p�塣~_���i~�q1�u�����g�!t��ry�,᥽���^�J��v����xX�@o8~b9 B�<~G_J��I��3��uT��Ӏ0~!��*;|�!�H.��XG�+?��HsΞA)9�^����a&4��Q���p�Btc_���"��"�f�HJ�19F���93��3�{C�g������t���c��#��o��qm�o��q{�K�[�@c|G�n�ل�y�;!��\�y�j�?�L�YlǱ��~�8�K(B=� �@V5�i��ǖ|�E]� ��a��.|F\%+���2y9��+%����Gt8�S+*t����ʼf� ��~���S;���y�Ɲ�o���/ˢ�ڊ5�;���z��S�s*"����f�^�C-���b�j�4x�w�KB֭�_#GAG^�&Vu+�p�Z�v���84�w������M��^-��&�  ��K�8��z-
�����ī�0k��C� ���A,k@�a���]?l^GI��� ���?>�����v�����0�|�ӽ�� �iLU2Bgְ�D�d�n�Iu�>?qkjX�ڬ�=��O�����Y:�s6�4*����������1��	���m?��C#����%��S�=��UF��~C�6c�x�I������@W��Ogz
�킽u\�!�K�Հ(s��c�΄"\ �z#�c��8p�F���;͝�#�R���5S�bo��\�%r��}O��cG8�h6kКu7T�'K��Jm
f����H��̼+k
_�#��RU'q`�NP$0 V�I�/�k�m5��#��*��e��,�C����"�T^e;��i	���s(9�,��2�"�n?v�0sU��w�EdP!���˜����F"j���#��O- ��$*6EQ��"y��|���zD%��T^��F��E��?2M努���h�mBF�R8��]h��;��DW�I�Yp
Z(�,����f�&��yᄯ�kc��>����EA�:V(^,~�����䎮�S��P��	��/�5���@_H��Ӑ@k�Q|=���²���wl��hA/����� mC�Nr�%�b�$Cܼ"����wg� d��ѰFN4(
ʬ*��ǲ��K�OH�)Ĝc�����y��1��<����z�	����ud��_<Eƒ�C+�D�xּ�5^b�|���7hlB�AG&��P�i�?5T���zp*���o�>���/΋�W��v9ٺ�+ll���ɰllSD�JX-�1���<��L�H�3qj<Y�ǩĺ\������eB�Պ�ul�AďC��!V�H�P�4D�X�f����buQ�:ێ=�총Q��9l�x�#4�
t�pMN.�y�Co�����CJ��I��3c����s�]uˍ����F��p+P�~�U���1�lݴ0�K��ѣ������l�	�Mȧ�H�Dt��x�����TW��օ��Rm��tZZ���r w��V�^��R���φ�.���Zj6�#��j��l]��񗱨�5Ͼ{p�9"U����Sex�&E���GQ��^���1����
��I�M̼�C�D�"��`ىm�ڿg�~���_��_��薝�Zx)��b�s���io�Y�6���'��nI���_����Y�?a�(Ot�3_�B$�H��f��ݵ7�C@63�ʋ�z�	\Ѣhߠ��Ԡk�� ��/��8Z�1m5Hn*�o�I�?A��K��(Q֑�l�E���g�G�����H¯�r��u���o�E�]ʟ8��33���4����m�n�"w!_���H�U��`?�r��	}�z���V�38ぐ_g���o1Ԃ�x�����5�؆>F'�c���#��s$"�����@a�0e�nC�)��?Fo|4�%M
.��L~�O�7����47¿J5�l,q+J���:4��/��5�1�.2�w&Φ�8�<�:�҅�c�����ԻYg썃D83�N �;�h���� c�������LJ�G-2Q4�%���Ƣ1�O�IaY�É���B	әޒ>v����1!\��� �s�"�S�8��<�9A���ʑ§M	'��՜S��p�f�wm�䣰��D��ogh�^�v%}넯i0�������2T��``'�9���gzc7SEd�'��.���aŦTc6i�ok����,�p��REn�J-5�Bڣ�b�n�H�Ȳ�������C��mzX���J�%��J�Q����MV��䞄�����U�@�{�$�R� 	��_��
��f~����<��N�B��꿬�dU����߆���>,U�����1}+I�;9�H)��`����P�=yBd���A��18�!Nǫ�B��蔖o7�:BLM7"���<ĺ��,���Q9��N]In1^�o��S�˚�{�����'m�:U���K�V�}������n�~|Ծ1ľΝU���T�W���Ћ�!������A�!��U#�2FA���Nt>�����m[/�j`D�}�^)�u.�X�Rh'(Ӌ����F��r�6�`_���r�o���:;ǡ��x�u
ؿ%�.�vW�BZf�|f���-#c�&t|4��2j���T@�������v��qL]��朔W�OʶcF=���G^�KA�F�w0b�d���=~�>/ee�. � �@�]�G�"�2s2�g���W��R;*�r6���-Ѧ��(��ƞ�C�|����}[k�tN��d�_K��R��T%5�
�7�e�%�c��*����k�XT��!�5i�-��^y��WNW�&���7��aQsǄ�'p<T2V�v��av~�Ǘ���rԈ0�"�f�rυ�/�jf�vɯ�뚕n�Mi���\�W����������s^&�ԕ��9���N���'�(Y�J��X�	|+G���&'4LV�-�_OJ�-`��h��K�/�ǝ~OuTp�!E�=x����G[�lR���A@
�I�DB?Q�EK��Jq�����I���N`�$a��+7��%�z�
�>I�y�d'�L�Q%��O��h?�p��m�A'Q�Asx�b��� �]�&��֊������8�\tdU˄y/��_�� ������ӣhS �ç�8�0VtC'��朗Ϫ`�r��0�P�i��M!|������L�����I�'iIrE+nld���g���u	�ٵ�� ��� �,�!NP��.C�>m���}V������'V
,.��q��ٲ���pOR%�A1�-�P�u�
sK+�ε�#�
A<��	:F�g1�Sj���73:��p�̴ܾ��u�p��f�j�#7U�)��)�)�KGp�5y�tvܠ�{?n(r�'��9_���Xz;�3on�)�a �5�Y�d*�3d�T C�� ���Ykr#м��w���.��>�)����L着��mQ�hӾ;V����U�����8���P�^���W��\lg�n4�Cʂ��Y�q�R#RW�)�x�����I�ɧн$=�=X����E]��$�x^�5�c�I��-F��T����ڳ�>��L�ǕP|�"<L��ǃ��U�Y��)z7-�������z�FU��ر�$������gwo���73zw�2aP����DH�ʙ�$U)P7��!��	+7���j��B�q�;WM�8h~�� T�8B�I8��a��@F�2$���4l<���硖�H�	W@.(�3��^�=1�D^��D��>��Ė	�M���p���@�D�|��Z@�����������k��:|�%Ǉ��� ���UR˱y�]D�ߘRa?_nu��֏R?!%�5K��$���*�#�z#ϩw!<� 4,\ՅS�S��5����F�I������_Z_��2B#ta�Όfo�'�l�������)k�9�F5�AӒ����"�U�Ipͪ$�}�k�W�X�����q��Qkk��
b�K��K��+����'j�_@�3�j�E�ҕbOP��U �cdzSӅ�{^L�
��Z�ۡ�Ƒ��)kf�m�_X�#�E`I�J�6Iz�V��M�d�N<vU

�9K�l�B+�ߣQ�2�d��4��&�l[YN���C���R�{�j�q�A*�% ��y�ܼUwY��5�������W��V�8(�qSi�l� :���̜~�HJ4���O"Q�!�g�k{��y��D6��h<_������� �� ��ڻ�B�vGW�ş���HP�X�x���8�9޾F�y��"��Q����H'� �;3���b��\�����e�U��s>��mf,�I8 ��+�n�j���T�,���+��r�w�۶6�A�ĺI����}��-���_dœ_�����3\ݫ�{�J��Ә'q΅E���� �_��0�"8��U<���C����L�v)+X*x�)��Q�ه�dPNw�"����frQIstH��]>�Q�bS�o�&j=�R&Ѭ��A\A�ЬsЀ|b�W��Ѩnt��/F�?z���x��_7�Ք����us��	����ZK �r(ba�v.�Bޕ{�?lX)v��{��ݣz��P��c�P���`Y�s�as�M92� U����H��2v~�L&k��B\��&T�5dR�=@��:`W��C#1ܐ����@��|߰�:X���r�㡱�,��ktu[,H:�2����XB�����O�U/Q��b�5mMB�hV�Z��V������EM��B:B��:�g
�4$��xh��QNG�#����#��-c�pRe��
���	9�Q4�"��,8��Q���&�U�$����n����37�������W�g'�!;<`L��nPN�#���ѯt<.#4�Xvq�g|��o
����U,'�'H�/Z���e������iʒ��ux��b��/���ґ?/�>\�X��ǭ�֤d��z�V�pmN�5��g�:*ph���i]v��$����*_WFZ.V�%��Gp9��*M�L��\w�����X�/�̟�/���7�Pg��!�x�H��D&�L�U��En���\P���7��c��k�N�n`6�d��Y��2Ҹ�b-A2��_�������ƙ�]��A���1�� S�ч�w���b�g��g�.���݀(D3-zS���	�!�]l�A K��BBb��@V]_B�&���I�!�q�Ǎ=e��Fgf?�L�j�Jx* Dw�H���*�}1H4�^憤�"�B��S	���W�!�s�3��K�w��- 㷏����O�^m7�Qd�n��(��R{F��U��w�^¿$;�I'���2Zz-�*WLbY�Z�CE�&j�"������l�z�sE)�y��{��v�K=Dr���?I�[�#�UG�F�	��L�wS���Vrk�5����j]e�ӊm*];X+�HZнw'�|�R	r�� ��R��R��זczBH�+��jBɛ�s�H�;��6������C�_/ �?���5����Oײַ%��f��AV�ʉ ��?PA���<MOMaS!躽������l6�:���se^G�@:I8���[c���T����W�ռ���3jZ$��gLla$�o��!�݅�i��]�)�p��HfV5$��FuײÓ`���#,R��5	�D���`��d�ur����
D@�)z h]��WUdPd��G�i�s��̸qFܞ�=�Lp� �wW�O��}�Gr/��Nw�����C&HNO�y�v��>mܷ�Bܓ��!�ޮX��R?~Кn-vy��5i.�])�Ak:�s�gп�W�
Q}����/u����pok�)LU*s>}m��_\�@�=�nR�H��"��V��T\�.���M+��	�`���`<�I|��3�NC�r[�FW~��X��'����V��K�1u��Q�A��6dJ+��~���FT�$��ω�`a�)��t���hI)w��������Vݼ�[�I�Fq��0L����E}0�T�-)��'�k������b��h��=���ݙ��N���G��%��3b��k�t��h��j)-���Ӆ�����.���ɧ�$9�Y�=�� �s��^��n��x�ט���G�It����ȁ��Nf�CM�NPמ�f�	�YMa�쳲$So��Q���(�<�|׮ڍÈ��Oj�j_����`�ul'���vz�?һG�E��F'�?X����������|��xⵡ��Hψ�Nу������&4�hK=����!m�����h�5�:x��0�^�O�@�R7�N��KI�ҁ�Ft����Yi-����Yb��wVޘ��s�4��A�),��^�'bd���XvyѮgI�FAK���\@H%�6d���a�D/�8 xL�=�69�Ob�.<^�v�jt��Et�O�%�H`v{����Y�����=G�J�kG��V�Q$�	��W�X�m
�+� �)Mf<�R�ʜJl�9��Ǌ�
���d@���3Zp�v>R���T���ʭc�·B1d$�>
�]%�=���H����d��C��Q֛فՅ�n�%�33h��l�d�Y�33�$�]�����4��e������1۝nz�?���ީ �~U�d?�D��q��QvO�0��%�;�+F��m��s������K5m)�ܼ��L=��������pOw��R���v(+�@��_dpr�|{r�d4��l�f����XZ�u�d<����R��.�J�@��,��K+�U������T��"�75PzP��'[J,p�WH��P@I�.�<h<���)_����j}�]�MBQ�d;�.i���,Z�i�X��ˬf�9��BmǤnES�"��Ô�=T��ф݋����O��0��.ۀ�%[:���ۃ�7	����xOzW�w��݀5��Q�l�oWa�k�<W��Idz/����\V�"�I㙻���氺�s�ΗWĵ�nx��ﴣ�o�ْP��d9T�2�?��'��y��4P)A{u>=Ơ]Aq��4F���kr�F�"t"�Q���B�2�{釈�c�Y��W_�`í��Dܭ�(s���W\S�T���|l�{������Z���%ͭ1��e���=�k	K�Z�Ւ.{���>m�#��u-�.�{x�˟��6���^U�.^ʻ�~��>�y)�E�1{�Z7�@�1���A�e��ۀ����F7t� �C䛧9�mTr{Ϝ��_����8F��X'�K;��;gw�<?���%�.����H?������*�Z%e��v���r߄��NI������	�(�(�7����f��G����Z�����w$4�&���t�?�hi[��{�h�l����4��4��4�8�v��J&�`]����������3 n�06h��̈0����V�~,�g<H}���P8;��-�Tߚ�Ձ̐?ϑ�� 䮓	Lɇ�6w�1�ш�hP�0_Xqi΢�����h�ₐ�s��ƈ���$��R����IŶ����������%���Z�t���{��x7�z~5��'��.� 2�������r��۸%�,�5�5L>��R	��G@tS�xJ�l̘&e���松��k�]�x���G�Ń�	\����f�b��`��Y�G`�gAzK��/UfN��`dg�AF�dPB�ǋ�!~���4��u���I#�&��d� �LF�+̐�H��8�c*����u�����t�7U�6i����� tYł�E/�-bHO���y���=�m����_pez5��e~�ܥ��Q���|����Wܾ��0�
��j�(QnpC<���z��?��Hz�k(����qt�����n�E=��&�$��C�ڲ`�W������(7��VA�����O�������%_�c��uBj��䵒�vh����H����=��6�_YO��Z�y��l
mv6c�ҝ~�˫l��$�R�{��1�Շ��U^;?�)���N�Mg8�Ç�6��=��"/���P�ާ�������n>f'>r�)��g�o;��\Ԉ��<���ׇL��!���C@OL�d���fe����;��o_��Q��3�������� �칃�Dz����,������T��+r�R	�DȐC�#:�a潳�C�s(��Y��:C��"z�M_�����JvҒ���l��&�x��=�e�)�emdO�W��`DAdr]����=[Mh��cx�d�N�Z���0�L��:�Q#�W�Zx�xj���Ȕq/�/��P�N�7n	kW�Yӏ��g�;�ؠm�E�$����J
�s[�7qM���"5:��6Qi{q�g���W�XШ� j���f�b_���}�~��k��:���4NV0;C>ع���Q�]��O?�پK{cy39�r���4����&�?�]�5PI��<�sE�pkE��?�KP��*�fǖ<�Uʹ��oTu�Zx��?�nhi�B��l�5��j�&����9���5Mj̨8A��^�+iL%�Z�R���j8��mWm�F��ahWf�w��-����3�_�!�DR3N�V�NLy� ,̭�=	$�����͝wd�wϡH,�;U���Ө`1�/ډ;ڈ��\���:Lr�׮$`�hJ�u�ܝ?U�#E>@�}���D^g�7��R�`wKO�>�/3��7��i��?�DxO���A�Tm�b	��y��a#U$�~�PB0���,y��*"?��*m�K�}$_�nH�Z�vIA�{iFY��f�l0�V�!F�r2Q�h*��\���j��܀i���qN�]���(q��>�=������'��ȧ��8��Δ�mr��@6��eog|`��t�i]�0dG�t���	���)�m{B.7�"��c�'� j��o��fe�w|)���k��> rؕ�R�	u�Q	m^0L�Ez@LƁq2Ga��1���3�)�9#<��������W�~d�+6��xo;c ����rw�����Us��V�áV~�����e>I�]�$w����Rh]�����
�V�惨
%.pZ�j񖡜�%�	ݻ(5J��w����a �=\�=ߡ��1���g��5S�aØ�����[�ׅ-�����������N]������D1'iLfk�h�,p�@���f}�)'}Dr�������+��v+c)�����������x��ۼ_KC�%[g'�
g��]�f��\'b�$�t焷(�;�*�ILJwl�l݃�X���0�(@}�h�!����p%3PYw��7��K����>C�o	lG���>�(����sΔ��SLc�w�A��ʱ��>qhtj�`o�nUD�bjO�b�z��"ɲ��Lvd̾�j��c���dAF��s �=w������<*e�T�b����fRv��B 
xj�24��(�?(�4�k���D[�}�������$0t
�����e�U���S'Y�ʷ�.�V�R��~FL�}p=u�.�(R��� �q��%�į��NuK�`�ܔG�_t׽�^*�8������I���'�� 1q���w<0�z9J��u;MҀȻ�_���%b��kr�m)Z�D^�6�Y%�F��>�i?��}��h�L�/yܜ��wy�z
_��e]��B\!5���7j��H-슄�[��GO�-���ѧ��_#g��?�$���U>���<"[�A�t��m�v���OP��lŇ�8�;S��Dw$�ϫTS���H�kIcBuֆ��5��%�B^D*k�B�'=>�ХU&�p���aNG���n�L.@��5��R�;,�*Ct�V]*��$��
��9o���
<�Q~f�Z��x&q��f�O|O���c��$��X1�R�~r�5L�m�v����n���n7��	�[���*�V��*ul�K����j�~�̺�B7��k��ʆ�*o�6�u������^	J��L4H��z�[_�}	xʠ������R�,���(����'�ΝhH���p�^
���|�@a>���Z�7�7 WGf!ӄ�Hn������~=et�vKC̬���fld���.�K�?�i��X�%U�.��a��]N�r��G1@��TX!q�.�2���.���e��Q�9��O�҃��S���|���0�B�J
�5����H	9Ȼ��m��vc.��=�(�-x0Pg���ڡ]�H+j����^����?WY��&�ڽ��]���N;�?�޽������9�2��}"���+si�E'1,���H���74���>��$��`�̊f�J�xba���R.����w�#-/@u�/k�M �R[l%��?��2L�������|h뮮O��f�Д>2��A+��~VѮ?�jHij���<wu�t6���4�	���з��qq�C�~���Aþ7��~K���'�����{�!�L�,2��<�`x}qo�|̍Vf������d�T6�cO���1��[Ye�Sjy����J�*A]�zBZp=���W+�%��y�a��}�2�u����a��b� >ku�?^���پ�����HP��Z���_��!��pϝ�������T��Ӝ�h��V���՜I���u�g�9|��M���8��2�6V�^'�M�*�wa
=δ~�T��5��{�t�}�[�br9��|2l��eq�[]��4�b�)+'������̳����ef���G�.����J:xK�Ͻ�R䚣\�q��B�E�ы�����z�g��e���h�������tuQdZ��~ٳ�ܳ?о���۩WN�U8��	ܩnCy�U�}7�AԯjO���>J�ۼO_�������'I��_�ʜ��� �}�;xR�:1>9$�c��_�o�d���{�G:�H��g���䚀hL�c�ﺩ�:���>�� ��̺�6�Pn���ڥ.h��P�'J3���88�V ��%���_;?��r�}Q"���@��`�9~;M��&xZ�?|���t���o/�L�(V7nz������fJ�z�w�o�#I�Ĭ�7�qsMVg�6-�iӱ��	J��tXT��T;�5F]���v��~���Y��� l&��a�3��o�yiV ��+�w5���5��C��(�&���q�DN�`��L��4dŚ=��G5�<�a�<%64��(@]�?++ڝ��܁�j����Z7W+.��/�\��]���S��g'��A��-R8�v���!�hi��	K�L��b�ԋ�4ָ9���E� @�/ų{��oV"]���`���U�F�A���re쩵�5X�������\� ��RR�81T��}��9|.=��KIPߗ�c�k1*�x9b��<\4���ũ�V}iD������&e�� ���E(�hY0:�v������a���$#����7�R�Z�j�)���Ь�f\�K��������p��'�N��g��\#9�k��([�L��F��e犤����4��ҙ�KAT.�_���4E�
ݿ�?gC,�-�NN��������lX肪�e�h���3��i��N�`N�����"Z^j: �~�B��06�D�Ǎ�� �{۵�K��,z��{H��ȹ!��g�$��GA�!�8#8�-�OT5���v�eW#c�@�S�u�����#�����s���|g@�XIY[��$S�8;`+ϐ[�S�����M�A�FX�5�/#S�����PUi�n<��!���Q�@l!ْ��דPW���1��,A"���3}�k��:?��6p!�@?F�1�M�;L��Ǎd�(|>{d��ɘ���� ��:_�*0x�`��>�K�Pr�Ї�%I!I0�f����y��Ȋ~EK��mㆮn��Y������9�8��5d�� >h��Qf��I6_���-���J�-
�� �%��������NKdg(��s���$C!�q��|�^�295R	Ν��Oԓ3'>=���}��#�?��
9�`��JW�z�X�Nń��H���&J�,����n
���^��E�FO9�v�5�*M	)����fQ�Vt��1_��=db{F�x��l����{�F�ܿ�Æ0��cK����2ͣY�0�A� �hMZUk�h���(�G6��i�i������^���F8��0�h�u_�3�)�d������ĉ�MZ�����g-�+�T�B8!B����{D*&8�S�ԝT#A�Ԅ�эb^*�m\�����K����߱���0i>z��,�R�����I����9���̇xh�&���5��{6_UN�v�㪠P��M%t��d�~آ��:�n�K�U���ն�ܢt��Ԋ-�n���}ǚ�]�����c��O�y�?L�o���B����$��L�lӨ����|	Nm>|i�ya��ܜ���ѐz�|���V�0f�)��E$6���*v��Z�����nb�e�x���$�f����Z_�7M���3s�+��3��\B0O֖��_�p|Lw�dh��_Ó��~$�!,ب}-z�T?��C�:�1��Yk�*M���E�b�R(���s�"�S�#M{��
�G<דż�#�'&d�5�R��\|���Wt�m7m�ona�}��i|�dS���N�����Ǻ8���a#p���Ѣ�N��B�M���כiK������zz%�?>ȍ���,vt�K�Ri/���1t���IR�F��U�;;�.����3������Q������G��;,v&���h]��XU:���
j��XJ?���{�@&u� (�l�O�S�)=^��dǡk��\�"U  �搛I��Jtl�RK����|��9�>tBc�ݵ�&�����T�md���,m�����e���~�����;_��:��jB\����JP'�4~/���wg��L��y�=ur�*��.>��v�������C��@9ٍ���-�����=�M/�u'�$i�TCT�Z�B���$	�]�������&�대� <4�b��~�����}h��N���)��V���Z6���a"����b���:�O�����f�~Q�����g�%%.[�T�n�T�)�O�7VV)<�|�қ��6��M��JwFeUb��WBM�5����A���N/����3V2#�]'a=�^���˥_�҇2hK�mG��)\�?��$mt� �}c'��IM(�j���W4Q��;^����;��.�Xt8xC����U[��W�m�[.��]��3��bK�.YRR3(D^Q�{Vo�C*�,��:�-NA�_�X�ZՁǧ���V��"��ge)�I�L?����Z�u�3�����jl.Q9W��E����´[$B|�s��(�OF?�1[��+"~�!*;����q�m�X�fV���%���S�OS����FJx�Z��%0V�Ĵ�oQ}��o/m{�m�vB0�@u�I�C&u0��*h��}�^#�UWo|n��w�X�y�MJadv�;<�41�
�0�5�=��g-Kr�6��c��޹ܺ$dƻ�X�t�em;P9�f�?�4(j��<#��l����m�b
����Aj;����4̤>�au+%|���L���xI�0��N n��g�ʜF{g��JS��O�ö��u�O�Ɏ��qlٙ�#�2�6��+�������s6��b7���m��B%���$;�{4�g��\Bg����ԥ�⤎^�����cF��Ӽ/���kG���4�;Ӻ/W�=/m�G]��^�1w#@>Ҵ���	�H#�Ve���wC�j���r}��B�eC�o��U��Ia�'AC�)Q�7ë
����e�I=m�D!�c|���P.;�WUk����a��u���'�z5�?[=Ru2�����\=���eBA��>�+_�{_)v4���8/���y����6��xa6����˦O$��������/��3@Z�����́��.��Hp52h0���4=)�}��?$��׷䍬)�}%��#�����v(���u���NF��s�����~FT���v
���B�3�p?lĵ?q��<�È�H��-yg����r,фћ5h}݃I��%���A���k�N��EP���W3	R���J%K9W�P�O�����­6I(�I�XJ��V�[}�Pa��KʶM�PM�b`r�C�f������fU�����(���W2R�6�w�x(S	�&�Н���,�G���G���_���vI�?��)�=jjT8�ל�v�[��L=[@������m���` �d_�0��\��6��%c4�v!j��r	'9v�UA(p��8Kv����V�*�vN�@���L��d4��������ˏD�<��<*� �ϸ�����ǡ��B�[��6i�Oo���
�Z�d�H��N�1'ֵ����Ʃ3�˥{U�� ��"U�Eln-�G�ۇzN���h<���A��R�}bN �$�����&�yO�nv'�j�[*���#UZp�ch��k2���x�ڼ���!I�A4���֡= �}dF�w�.i�V�9�ܨ�1l27��]��QR~��s���5Әn�+���$���@��	�i/����*���V��C�x����X{ڞ:�,���l��K[�rSyol�kJN����lnϋF�6�wܶ��=ȁ+�nE�cE��+=b+��~/<a83>���&dl?�c�8�d����~E2.��������ג~j�YѤֵqN��s�ig���}C�Xn�I��3Bm�(��E��ER |ȣ��q����n)g�hO��RR�av��XH<%\"�ձ�٘�p�����2CIZ�66m�P�:�lS�j�B�7�\�/��^%zť�r!��
 ټu�C��(�h?2�C�S�d�g�Ŷ4^&�W�C�/�K������31rF���q��~�g�_9�x��UN ��lX���]!�`N"������Sx�,�[���t}�Ճ�WC�X�78�W=�	-^����毾g���ʍ܁�H�;i0w��7X��F"a�x��h�ճ���k��b���႘{���f
=�O�ᢕwiw�*�FC���`i�Y_�Y��zJd��G���Ys�6��!,�}?�?�d�#�V3ܩ��p� �{����mm����	;�}D�0���9U����tL�>�[�V+��Ƥ�l��k(᮳&���5}}�8��-F�҆�$LՕ�9�u��`Q�U�|�M쫮�Dі�}���ˡb\Cn�Џ/��b��Xp����� g�����u����?�a�@h��O����ې�xDe�S&���2�#�_�/(�iL�$�B�ψ�P6�"�9�Mz`k1���jo[{0]�	K�����F�!)����h��\�K�vh��(~Ƣ��w�V�>�6=;��90/ֻ����@��i��������k�)>������d���%���a���Yǋe��$c�1t�@�P�t&�Fԟ���[�E�o�b��r�b�֤�Z/�@�ޱP�q��ӎ.Q��\��	ܤ*����5yZ�2/N"�!q�9:��g���%ʺ�&��mE]#�oea�������w� i��������Q%�v�p,��b��Jjކ'��SS�d&~��l�bTUUjjˤ����9�rQǕ���J6ߔZ6�����#)��g�Bi�{����}�����Sy;K��5I!�9k< 0Eܪ#��C,Uս�ɠw�3�n1c:�dm��b�yx}L��"��4�̰1�����"���
(Z��A����i���o_.�m�
d�p
�x�C�U3��s���A�s&r� �(*ʶf\i"��s��{E*���~�1��m 3��#��~6�t���h�=o(�6����<ɱ>y�=�X:�yuTӹ���&��q�駢z,�\ްr�+МbD.͑PoJw�@����S��������wm̟:n�
\\�+��2ٔ���Ln��!K����RP���9$:�i]��oĹ����vk�%綏d1 ��T��A���4e
i�����>�VDvFj�u��~yI-�wX�Fd=�á���!
��0"�D
��թR5Ma�̏{ӹ�>%-%��A��9���F@��l�0k��X 0B_��Ϲ/j�{�фA-hN�{������Sj�(-,�����՞�=��Έ�Bq�	H� �}�SO�@ Z�~���U�a�.�īDW�:N�����é���������ʮm^PF��~F4���i��ƪ/����Qm��b��Ԭg����l� �rkh��;9C�9���s������p�/��S��<S�=�6�*W1�L z�X�3郳���[��c�;��2h)v��'1C9�� ���e���0�D�)!V?��TS�{�G�I�ܧ���<���߲��GCyY���Nz�9��]��x/ Q��v��j|�,�A�ZG�N3Ŋ\{?���Ұ��"֓�x�
U���e����Sp����f�l�9I{�cT����!�*�-�}y��V��Kv�2���6]��:_���(���^.���$��#�dd��z�0���Qw���d/���?�$�!����%�}��>w1����z\�3�$�о�����n�ޜғ1ڨ��`��U�祖3�qz��<������U�眉G*�6��o,��!)�>�k�Е���[��g�Q��w� �f�cw#�㣆���s���y�4����`���%��C�P�ը�Df}gHz��ԫr{6�g�Z�?��	���;���X�<H%HΜ��k�1����Uq�۟RD^��AJ_��er3�1�$S�?����T�����K�z�����,ws��/�j������p��[����JB���Rf�����^	x��g<��+�y�)m�Nl138���}M�P-���ʂ��.��OAF�!��F�TJ.�*�Ŕz?��Մ��U�˸K�^�cf���k�V�3Vڭ�(j����Q�6�rK��nE�v���"��^�%� ��E��T�w�$�!��Y��/����u�	�1xx@f��H��������kF+�K9�k@�y݂хR�}�k1�g��h� � �ls
`k��h.�d���]v/Iߘ� ����C
(�F(���{E%q�7j/�O`K�>Ww������i"��L���gφZ�YDs���Qe$��CZ�Р�l���y�
�[6�;У�?FZ,�P)�R�$k����SH�y���#���^�+o���/l؂O�K�.E�&g],s��:S"����8���v���w��<��Ӥj= \|E�U�̃���+�*���q�=�S�F�ݩ�~���a=ϭ��4�&̂m�#�a�]�3���P��-��~,�k=��f�]M�O�Y�t����JGc~�aGW��-q�Q��d�,@�j���$h#B��N7��sQ$�F���9�V��b�̧��YZ�N�7ï3ߚ�C�1*A;6u���m3�Z�5MA0�R���&J�/������;'�D���q3W/I�KY;bF�?Ǩ$4v�X���)F��W�e�@���F�5q�����y�/�S|���5�Q���`W�o��[U��C�*����1�a(��Q��/n�^oG�xK8$��w�@]e<��Gμ�ϲu�2%�{6Eٝ�N<�O<����ح6h�f����Kx�ǲ9���1�DJ�컣�#���\w�_�#�I��|Q�1�*�.��?oF�]6G9`.��#�aKI�U���k��s�s��C�O���+	F�n/,`p�q�V�����c�8���ve:t�|����7x��brs@���X{�E������
j�9I�G��=u�8ޗ���<٭��>#Eu�SO��^>Tk�R����ӏe@8�������M�����$>��W�!;�͠��m��J�Ȧ�b�V�zo��%K����Ma�v�xt�ǆ�2�����!��p�IWm ��%1趱�!$8#��d@��H�z��˒C�]��F�qmY��,��"�Q����8ƪ��r�-^ǹs��������;�#�Ƿ=��? ��9-&�Q��|���Ա|S	�MD���2_�JΪV�� �>8Q�L�Z[3ŕ�_�����v*��*r�ͭ+ƕ���� /���Ϗ�b%dR����CʁF�NƲ|��,:��Q���p�}��=��=y��?;���wG�,�������\�hBM@#8��(�M=}Rʯa��s��$�mf���P���o��. �)���sf��p�㕔�P��a��_@�Ec�\�3�D�S���8Qc|��$h��ڽE��B#.Ms%�*�H��uT�s�3���$�M�E5˫a+i��
��œ�B�ue�Orcg�U���������<��$,@�("��R�)�n�-;��R+�t���g��J���o7���	�G�Oelt��|fe)�������ﱏ΍G��4����w.%M��9'��.:����h�C�D*w��TuyR�KF���fH�,�n��A%��q����rnyA-A��Jk=����)�_j�R.�
g�Ǆ��E&����3$�vb�Hh�%�]���_��#�Y��_wr
�:#qm�g}�8�T���:�G�5s���ѰC�u��k��LQ�a)y.����ϔv�%��lX����;~�?%�A���y��W�[���4� EZQK�,b��8 '�ǰ�7/
��C�#�!u���8$��. *R�K[C
�"/3&d4��� P�Ll�E�H_9�>��c��e!�-L&=2����5n���r���2z�s�3�!�;#�E��T���&��U�*�9����X��nn�v&��E���{G�hl6܁��C�T�u_f���,œ��D7�2�l^7�-��|���t`
M�:_����K�sY��٣�_���c���K: C�x���!�\
�nv�����'�.�z�k����.�/�=$�`Mx��f�z@�jY�cV?-�$=o�����L�f�SN�ːH�4�$dmk������h�5��ڥ91��u����ӏ�kk�\�k��Ĝ!�#OR@4N�n;�+V�8�|ߔ������v�Ȃ�[?/%�	���h{�婰�"W6�I�#;�C�q�ޘ��#B�����G�{�Hpֿ�0ю*�7��k%%���V��ϻ?%�a�fD1g�z��9$�
��֛��v�2��i�hee>�I7"����$JN��o����]����wB���2�y��WSN-}��{�smk^�Æ�x�4�?ٻF��ʾy���gF�	�z�W�~��s�ܱdֶR�(%��X��#	SEa�6�6�7��[� ,RW,˾+��kз�4��I��(B�N�gz:��%~�O)m���T&�����	�J4����e��4�.p���}Y'�г�Ɇ/�l��

��J?03+�����4.�*����~�;�ԑ�v������TC)�A�lv\�)���P�����&G:ɨ��o%\:Y��0�?���~�#�_^���~?�2�uK11�J�?F�n�~	�mPj��$vs 2�p6��A��1l������'~&�]#�����8��ly����%���E�r�٨1�f�;f�m�Xj2v.�����L4�u K���D�@�n����ڢ��@��N����P����^���.e�9��ʹ���Jq��a��Q�!��(�7?=/�����yT�uz�.�!�M�~�m%�R'+�F���5�^6��Ѷ/^��J�$(?k/9���3F�:ڈ��?���!�5Bݴ���wF��L�z?ɆՒ�ŃߞD�%�A\�缵��Z�h#.�E�cQ)t�`���`�P<���JL��P��D��drpT§�8��?��8�Å��a�K�Ә����a����)a���l���ܯ�w:�F]zE�Z(.���
w��/�!)<�Q&;�����3H ���9 ��O��màQ��i�Ws��~eH]0��u1c,�
��܉a�s�q�[6C�����<"���?�&' �����d�>8-M�ڟ<�o�M(����N"�/owà�Ak�DZO�i�B9�)�!�����2�����Ʊ1��Kp1���׹�R���h��:O�R-oL��9_*K���#+H�-^�-k�T#X`w]�P�L�N .��5t��8{(F����L�ZN�E}�ϕ�fN�qT���%����o��C=���`Axo�iv�	�����'�sH૔�m)�y�.m�6��9��
�bM��ԾYt�4�-Gq�;���K�X�;d3 ��D=`��?��y,��4ulp��ŘA+��җ.������&�H�V�9�wl��P��C���.��2�&��g>��x�0u�6|o@��\���.}g)e�:}�L�^�਴Σ���_n�&ᆊ��9��y������c���*?��Px$�9VD���~:��
���x[ka{JZy�"��G��	�ڲ�}�Y�볋n8�j��	菢xoWNL��$��&bY�OuT�;�R�cV�����ؕ�����}���w�-��n��N�L3��r� ��>u!V4��R<=N��r�����Jč֋�E�o�U���k��K	[մ���=8����qGV�����?+�����pCkl�A�"��X~���A�4��K�y���E�~}^��t�8�\D7�|K��	��ϗ�:w{��F�|[� ,_y>��[G0!l�R*�C�������Nz�c8�d���G��=I_�H	��Hո�a�4a�?�e��}|4"- ��CG��Z	�r���A$GH�3!��.��Y{\tb�A�L�~{�q@���qnL�]jU4�#j�/��'jcZ�������R��z:on��O�����}�c��Y����я��Pɞ�(.d"4���	قj�8�LnA1��%�[FL��g��\)�������V�d�.I�e�9�L/ؔ��}�ƝXu��"-�+�k4�:������}"�H�������E���걤���T��	%C�����m�Ndj>��[�@�L\�2�+��[u�~9�j-������Utg]9|�~�F�[c3��ʬ�'α�ϜLP�,Ea���m%ikl@$�@ٕ�`�v��6
Ph�u�4��a���㯭�6�0��Y�$L�?wS��ZqR�En,]��~��G3�`g��K���5-�k�J�Q��&�v.���FJ��3^�\f�P`�gݽ�6uS��F��;��;S{P�P0�3v��5P̻hD�K*���p���{��Uѡu��U��E Ҡ����yT��+�@4q�	ʽ�V*�r����t��#���
6MT B��Ɔ4�_��#�c獣>bs:m����cD�W�xRi�`@�%��oAb9
��}���F�A�Ffg9B齷��G�u����Wu��ѾA�e����8�ŊT"Mt�'M�5ՇN�o�˿.(;?P}Km`ψ�ν�0�i���;��2�%)�߫����=�7��M)�Gܐ�����Z�	�����_��7'}���M���P�+FCX�+-֋�e��"�ۺI�*�
J˖����,��h�K,on?/�?�̬�x�q�kHp�{k�[��;h��?��b)m�!�B�`Ma+�i�]p��״Y�;q���������{X]B�q���b�J�!-^m�87�����ň����a�U��-�Ɠ��Tw`AI���d|]�5��X�tE$�ҎV��S�(Z:E5�ò�^���Ӱ��'��b �Lɺ�Xgp�\'���a#+m㛟���{��zu�<2���R�0��r�r�o)�r���=���O.��\�H9c9�b�>����>�r�;j5�CUi7�W��hE�4S�Sk����ǐ�k�9Փe��0���:M�l��T���/h���w�d_���M=?`�H�Ϙ�B��Ȼ��� BFe��5uQ�շ�ߕ�H�9��$
"�������N�ib}C���z�M����k�I��\����^^�T��T��Y.ܷ��8-�J߼	�O�O�����Ěv����L\L��2�R���*N5䃊�5"�2����YO	��^W�����RA��&�-�
	���sʣ��S	�ɹ8LuM��l���0M�V�֪����G^<;�.fB'�;�� �mk�-��f���_��.[0�JL�7�ߵK��?�e�V����I��~���n:Sr"��_3_%ߚ(@�&�1�B��V��J�=&�[O��@����7�tj�y��|':tP%�-����x�˽���9�TY�K��q��Y�� @do'�t�jM�!�j������B��b߳�,c`�q�^�?������4��$�V�%L�x?��f���������M��rN,.��̌��Dy�G��|�i�)��L�s��y|�x-C;]�r�ty�3��|+�W�;=mbt	��k�g7���^p�Ջr��MB���&>���SP&�7���v(��s�_�G�e�YT 0�YL�kp3Wt~h�迋�zf��i��G�u1%���L�@�0����"f�q��4D�=A�>Hi�p��O���X{�K�vj��NN�y�_4�݀�y\&��Qv>����	��'���1��U����kMt7�g	��:���\���֯vV�Sf�*&��)���%S�E�é�?EJa�!T�u�%�D2et+h^ U�+�y��a���P����:��N4|�	w��~
:��N���@4��܋��):��"#_s��s昌
p�+:&�,*�I�=���Vi��,����%X��D�T��}K�D� ��#�<3�]塇�E���o%@�oø�ф����^͇W�1m����4=�'��"*b�t`К:%K���k�E�kWhv&&^�̑x��d�;�t;p^t�Z�r8�h�/��aa���]����>���y�k�ɽQ���PyʍЮ��
�Mn�_�_@�a0�mv�%�\֕}s�E���hW)�������d0h�ȍlY����NP���A�?��L��+,����R�����>�������A��}�DBC7}�֬��\�gGL���ߝ�F5��`��&��u����FX��k}��j��U��Vs��ؒD1Eb/�[��Sg#j�kZ�9p�Tr1
D�q�$h�����;9�~$K���.���7n�i����P�@b���)��i}ږl�2���3f�˭���6g����^�】0�ψ��XEm���b"�>�TZ隟�ul��)Yp�/Ut��3����gț)��ߒ�=��7�)�{���n��Ò6R�=nz���F�9؊���é;�	�v�\����v�Ga[�5��A�>#��f.f�Za��Ϟ'���$��%�Vڈfj�Q���m���N�X/�����!�{Q��GP�l�Q�U��o���l�t�}5_�h��V��P�	���izCǐ"
�AW�c�gn`9���RY��^!�o�ZI��T�h4��R��tu���nno�x�Th)t�Q	��2Cĩ?Y�I_�xB����F|��+���d��>�Ew���U����:�yŠ�u;X�+I��5�#О��/��EՋ��W��И�ޞ�|zk3���-���r��yԌ���������MXBc�������T�`�k�2V]�F����P4x5�f}1~q#���Ru.������t2?<d�b�@4����Ι��}e�H��`h��a�אaB�Qj���*��Ҧ�s.ԦA\�8P�_��,���+�����R�_Ra,���n���i$�R�Vp	����"(^��g8���V��-��\�N�ݔ���YwSy�_u��7�	��2���@�(�BƸa��Q��i�Y�Ѡ"���]��v��U�g-�\����A��bj}[��ŀ�	zdczf��� o���"���'XX�z�M�bB/B�򎋱<�}�ރeVѰ�8Kgq�(�U�\YKz��8�H*�a�(�ZE�_��&{x�?��L��>\&J����}U&"��`��DQ�a��$1y�z\��-@���c�A��b/2PQ�򻟓��S�X�SV\	�q+�RF���@��܏��>�H\����$f�����ݵ+feL�2'���rC��a�j�� ϲ%��)/�3�d�mB�	�T������ f�VԮHZH=F����z �����\�2����2�M E�m�C��L�B��Vb��\I��]������h��ÙT�&�Y���A�^��5��b�������!����B���:��s@���W�.��0
�����v9Eh8���	�V�넼�uD�d1�u{�n���8~m'H%�O�!��ag���*����Z���1�5O!"�����N@�?����(��9=�d�ͮ՘|#����l��\P$�c? �260?�p<7[�b-�oحY�
���o^Ps��DR�G���R���䐅�3��������յh_q�0W&�w�`�iE��5�_{�t��8�naMvZZ&ߐ��Z�R�"�Vx�Vk����8�γ���J=[e��|
c�44�G\N�pk��$���=�Ig�U#`c�J�U�� �+ּꮰ��[�h0����6١�8�-OjLImS���IO�(=RO4��vSf�!�e.y.��|6A�"�� j�"9�|��p�=t���9h�G����+��Rv{�'c>/b��J�k����Ă]�.��w��y^��ت�)�Gk�.W�7�͔#�����r��#����Ʀ�V�k�wm5;���VT�� �(�*[�JL��<4�4�g�15��VnhN�Z�3f�S;�9�����"�1�'B\���k��h��˪�T0�����+���+Z�O}��b�0-MC�|�{���Cn��YQ�+M1������������-N����[�IIO1�<=��G�|ڏ��J�~Q�ZlQ0 8)י���]��jQor@���!ie�a� k�j���� 6��^�h>�&�t�-�-�<��w�ݔS%i�eԳe�{���E�]�]w�T�_�%���t��Z����s�Ζh2%���ւ�
1䳁;]ks�{$�(&�
P��enS9K�Т[/9�m4$��Ī�%��ލIo\��	�e�2��g�^G���&b�;Բ���Y{6�s]mN�,u\���!̥����M��=�$��0����|ԣ��!mO��w�����[��oy�H4��6 �3�и���N}s��SS��3�%?@<�¹&�� ��k��e�⤩���FcgK�L�
! /	�_������r�,R���T@���3`5�7�jA���:����G���j��U�ʻ��z%g�������d`�� �Ĵ!��ʪ�.�sLRHYoc׽�:f���,�y�<:�av��4�I��d�)���U7�����kƧ��l����6v��܄N�ew ���C��^H,?���p��޺���0�W��~"`���a�b�t��N0�,#A�^P�"]��]褤���΂4a��/BҺU�: ݒ�4y܂�1����M]�0e��7X�PӼ�x�7X��Bᮨ�+���K��%��2`4�﫯E�w�?>0|Q���y��>5���F�l�ǔ�o��-w��T�eO�Ԇ-K�������N=͖)x�}�.��i��t��g�3D�UM�U�0f�{~��r�[�K��T��>X�!�p��!�<x�I閳[��c�k��`��9��=Vv#;�8>�E��!����B"t1�ß�l���z(E._ ⼂C%A��!B�:�i�f���Z��n�C! W��.Q����Qw�A�4L�Z���1��hO@T3�V�e��J|�#���� ���'m�-���#�1J��`��}
���/z!��7I�w�lk˶�u"y����^��h[d�G(.���;�ν��.+ꖗ@��g��x��U-_��ѪP�XuL��Gْl����i��F��E��-*��_$^�e���Y�q&��9�z9��z�/�2D2�N��bI����O4(�R���z���C�.=�s���Z �f�T��_�N#"�ͺ�j�/QB���e�j����b�'.	����9�EtYvo��o�m@��Q�K)���I�1p)c_]#(����dP�Xw�u:�\��6��W���A_��r93�o�D���Ʊ�~N���"��T/�"X*���Z���C�~�<|S���l�S�^ "�C9m�HQP"�����D8�xf�ʡt���\�&�Ѐe��S��1��P���dYL��B�ژ�G1�,>A#/.C�:�V{��J'ƫ4�t�\ �Z�8���z����Gx+�!x�ظ+J��`o�p�>�d6�UP�����g����Y�r���/��K�X�'Dr8��;uU^ӁTt�����'���=��ː��`W5��~�m�I(�ĈR��y[!h�1�GAɌ����T��SŌ?��X���p%��є���+��MOO���+c]�p���m��_h���+Cr]��ԙ��a;d��nD��FQC�J������P�bXp����8sСwIr�(����j�����/kv�\�/��ɕW�ĩ
�,O�>y�c��@Ka�d�K	��p�
�!����+�]��:�aQ����yS+���^�"#յ�,̈⼘�$�+�-��A%�H�F$�t&��g�R��Ԕ"��+r�T��U��
	�|�W?7���������$�o��O��$���uՋ@R�a�ԛ��A���b�.a_��2�[��Lt������@k�	p�}U
'>�*Y�c�+t�����ۺ] ��~�m��#��h8קٙ^G����9f`닣����?t�&X��;S� �z*�Ƨ�2�=T.�5��*�+�X{S�!��`��W24��b�Y����	�\���	q�F�(��hl-�Se��-ɰ�ڂ���횓B�69;� �-��9��]�8��(�[x�%�/<���8_�T���;���3�-zw[nE�[L��q���H��'֡����1�v0|Tw��?L#c>�{$dWt�0VX�ϧF�*��;B���y� p\̡�8��AG�!�T�0�34 �Qu�����^�ve�!�1^���:L�Գ�N�#0�ʛ�.S�d�f��ʽ-t�
��� ��OR�j��&lk}8߉ߵ���es�e�6)M�Βx����/ �P��rwx;W&^k٘�}s-��;�<� ߋ~*��2� �t� 4���`h�5�����-HE�$��Sc�s`-o��w�Pc�O���M����\��gn���pQN'��~jpf0m&�42��&�%"���� �1�g���+��Q�D:0o7}��E���k�l�H*nI�`����h��!e4'��^x��ذ�8�<�~*���pRE�����e�!`��#�������yh�r�'��U ]�S �kбW����k�oj������>9Wg~�ǲ�u)cӷM&o�ܝa�}�9�N4�o���b�CU-	D�7長�,RJ��R����3��7Ą�~ҿ���2	��$�S�>�EE	�ډ���A��'/�{=��P�Ig�Y!�O
�W��NЫ���}���-�d�Ͼ@����1���g���o��a7,�E]�]�]��W,0�Sך�"��϶��(�Ӆ�����؏��;��A����v�.I�+�~�u[l H;����C{�������)n��g� qx6v\#SQ�wE��_�c9"@Ǽf���C`l���,*l_&k�Z�&)b��$
#�A���2{�a5l=��p�%����!�):�4O��<��3u��6�/�<���	�����u�$����8��3�����O%����_/k��ɕ�>By�\n4NZ�f�f#!�%��s%<2T�wЉcn�<O��h�K����Ŕ"��^2I�'�7�Y�iW/=�UL������]�L�/���\�T��ѲH��B2=p�P�ḇ�H8�\�Sհ4{�&���}w��~��?������k��n�s�])Ɋ��"�ϸ�!=���ޡS�"/w	{��#�n��+���R'�sR���S����������f؜n^@ר�P9�%�K>�C���*��^��L!�tf����ñ멈q�E4ke<{l�Ї�*��/q7�:h��Jv}|<w�hs8���=z5"��e����q��y8��N~sg"��0�ԝ�)��������|�¾ Ŧ��`��x�O0���Md����E6��'#䘩�vN�8!�h�&읿ٿÖ_\m�7����pI,䀿0s�ZT��f��=B<��z��� ��*�kQ'���?r���]Lt㒌���x���3u��Af��$z�o�n�7��{3K���	��������Қz��\�����M8YDsՏ�V��|Rw��z�(ZmsfsM�ފt�w��T��a$ҁ���%����o�_\>J��R:�N�pj��
i���|��.[�8z;��չ���^)A���a�	3�ó�]sXC{�Or���6qC�i=ovSl�3�<yĚ?�L� p?
��q$��Z1�\�+J�hc��|���07�|��K�"�g Aƨ?����-D�zE?�\�ē�gd�������N��ߴ��jP0J��4�t	�sZ[�?�q���(�����/�]���L�.�U�H�}+�S2��ߔ梅����C�K����~"x��J��y��W:��[��N�G�b��P�#s������*7/���C��?!Wq8�Q�Ft����N� .�C�z3���Œ��j~����0"�83�Ȭ��#�Q�0MxH��ah5�Cl�;%gҰ�{�?nZ�����p.�ɢE�E�R�"��[�d�ؾ�;��������/}��XW��������x�"����y�}�Kغ��g�/v�վ�e�r��-�g���ս9����5�Zd��l�y=&5���Ȁ������	R!�ο@:&�^W���A��?M�q�ۆe4�q�L���׋�h��0�B�� RM�ex:�����#삓��~�G҂K��F��0 o7�%v � N�0�N�����35���0�2�g��wL��~/����y5�#4�˧��Yx��x"�<i����d�A�4������a��>3tR:#����#�x��#�`s���p[3B�ZvO�O*H�!5�A�a��/�o��G���i8���#^&Wv-���o�Q>���.�Fw>#3+���h@2�%��J��`�fQ���Jz���>��}�m/nJTO��lX3Xb'��]��7J�����vd੒��y&:����oePf��
�|�ms�fz_EE��,K�0M6�KҕC�w���� ֌+n\��-zr6��h^i�K��/�0�C�E����Q�S���7��4י�L|�6D�^�qW�Y���&cq�j�e��Q@�h���5�Iy����}�	aW������jB���Q�@��ٽ��:��!?������~.�
�O�G8�ğe��=O��_���c�j��Dz"k�P6'�lT5�^�E�.ĥ|9/�߆[���H���V*�5Q�>�����Ày�y�l�>�!�zA�H��ac1���bu��0.6B3��:���|!�O�e�ô}��)g�) ��KJ���h|Y�f�m%��R�ߕT+Q��Ez���:��MC�H�n/8d�NY�������g�;>����Gȥ�]��P�)$��d.��	��ھw�0c�eO��սf�r���o��|��	]��о� �Jx��t~{N�]��	�Ɂ�#��Z��`@�.x:�QAIځ�qW(�=\���_n�@o�䴔�<��&k'I;�w�S�"�8��X�4�!|
O 9�<���y����YSc��5��u �oZZ��y�>����g�bH���JI- ������ư�([�p�de��M��� f�>�ct�}��w �]�R�Bo� ��x$�я�n���'�v`c�rڪ+>^`�C�7��r�m�D�|�ym-i���	+�G��� �ɇ>�����w
��� �j��Ҟ��ը}��d��MxMaƱ��ZB�r�1��]��^��)���[�!�!���Dàpu�K���j�iĳ�i�*���?xәh��q�jb��1����m8�K5���<S��5
Me���"��x���3UI�d�.O����.���V/���F�$�9��8�v�[�S/����Λ�Ѽ�L+\X�$.%uDc�\�ݟ1��A�EDgXX��+!Xݨ�N6�a���a�A�!��@�dl�8����Z$�4)��t�pɮ2>S�������qQ�������LUM�r���f�,��� �������3a�W8��ϛ��l�� ���r�h�YEC�>&�G�ؚ�\g'I�g@���U�7_�������pPD��)�����^�J�pN�N��ݑ���d()NMW�w�D��l~��-[;Ed�RC������j���M
 K!ȫ^gg��Ag~���P��	�V.�Po+�&���g�E�T����,%՜��u�[b4,\J�Bd�l�F;Y5"CZ��s52�j	�X	Xg	��1�B�n�')a�
�ya��E���y��~�p�{�|-�6L�<�_���Q�ڱ�_+�ǿ��8��v!����6;w�#8x#2��,;!�(� �O��(��R�^��c?����.�����9�-lo�V�W�x��l��� 	�	@�f�#Q�iC׎g;IA��xWP�jsw%!�f�Ԫr)D|�/4F&�7�lG�LAF���<}����pk�=���I�P�d�Z@ԇ�85�)��2��Oe^�2��e����g�r���0w�$���h����(e#�ơ�n}-�>3�p!d�omX���i�.��u%*/D~���ܫ���܀pM�h����.w� �i���WP��u��<�3���O�[6*�vӹ���^��`N	����<����sG�6��6�V@\V��ߘ�d؄����Q@�4I�`�-����.��/%����'�1ռ.@x?���\�b��+�e+3]���:�8z��ή�m#ϔ�Ð���`����d���q�VÚ�>���u��+qQG(o�n�F�R׮�^��rn��X���0Hc�4��b,]`���G��J,hK?n������r\br���y!�y�:�'|��K��4OD��h{�e^���aNρw�:Wk�H�˥=��FΞ��3��>q��b��;�9dK���_/�+W �h�0�~l����<\4g�@���,�mJ�i×�@u����	s�N�#O8z���7�|�$|���cJ0õn��Np����"c�>�-��#�8?����^�P�u�O�d������ y��蠢��������E��m����d��sё8�KL�U�~�I��W���f��7?����̌#1��>�Ԩ�3B��^��W�QW��s����#��έ�*8C�/���ځ$F�"C�+2�P�b�S�b׶��/p�v�!(����1c�Ì���1���T�p�ڏ%T�Ro)r���!MH�1�jl��q�,���\���]�rX���t_̱������/I�T�����Vʧ����B�ԋN2�͜!�9x\�:�~��
�+��%�h�&�K{�1�g��A��(,�ǽ+^D,��w}_�Z�ʑ��u|o8�&B�ֆG�K�'�(5�����Œ )�E3u���$�KE��a��`9t2xr`�Z��+�!�RJ��-`�%'�Æ- �d�X�������s�/�YU+�k�sP��!�@*�֕��:�}@Iu�(�7�X�B�H���L��,C�^�,��,*��A�Md8���ֆw�g[)���x��|E��(�閤yO���X�����oC�sed�t���eF�h5!���{��&�g3� ����<���nR��E�׎}���SXyu(o�[��� }gfP	YGm�<{�I�] �?*��`��|w�$l�:�f]sQ"�%�*�|by�b�)Pp����[?A3��/Î���k��K�Ųo�KTN֎�}��E��#�7��ԛW�P��w���B��	��\rAQrhA�3�E�E�����q�צ�]�hm���tn�ա*�n���1���߳�h���5돷V�F@(iђp#��+��J��E	!pv�I���м�zbM�d�2���>W�5&Q"]����~��xk�r��	>�-���N9��aX��^�8j:�Α�ʹ�"K�j]�iJ7��Z|��:�-8Fݏ4����U�o�l��gikR�^�l?�͸ӏO37����"�I�V�<^c�4�l ���3"@�/�M=8�TH�X�� �zƏ9��ɪ��￞��L��Y�[��Q����O�ZV�㈭C�h��À�ޜ@q$�ڛj����<C%s�sWx8PUVV��EL�kW!��V��C�7J������DG_=2��*�|(O�Q�� ����{o�%��K ��Ja��P��;e�p+ÀN��yO�.����i�1������Ϥ�G��Q"��[�\"ꥏ��,��{��=��w�h�ߴ]PH�>%����P�g�T��~�<��E<��f�F�_l�W-ֹ��[�^� 怲�q��[�3ڃi0��8WJ:�<��@h�`��m7紸a�@�{��您��{�U�Z�ۜ<�#�m8rm��&���\�\yG��[�s��'�[_���f�"m�CVjp{�>m�$U�����tc3Q  �u�.~���]4*5�&M�ɜ.�s>���5A��WtF:��v��\�k�6�:>����*k��m�Ø�qKJ�h�i
���ͼ[�#x"�ջ����5P����Z��[���ܘs5z]$P%� �g>T�����T3����-Ŵ!d��m�{�2�����֋Lȸ��2������O�s�U�-0Gm�C܀vMI����Y��Q�)=�J�
&��<Ko�>Ӻ�f���4ˢ�M�ob	�[0�F����	�i� YtĲ2��+^��'N���M,S�1���ל�/04����W���)'Г�p�s�Z8󀹶e6q������%;��g��T�Rt'U��͖��0)�;�ɸf
4��1�l
� s�\2��1��FF�ݬW��߽��9�~��v�R��6.Xץ�ɩ��(c�o^����J��YTM�d����v�U�p��yLw�,�sN�;���"�B�W|�P ���v����)��USi��9��g�#�@:������8���6[`����-^���p��f9pM s����d�M����
��샍<�+N���>2k�������Zݝգpl�)w��@|�UE����/�P��S?`��LX�=N�؟�57���Ǌ�h����0��e�Gfi �!Q ��2��,)D�фr�� ˢ���s�I��5��4�!Ĩ��*N�6�)E5�ʾ[+1%3�Bl��@�@ʧ,1�5��5�u�Z���㖏-+kZ	����5<D�	�@�y4�VUM/�D�,����t
Q�MW�]=���5h5�A�������@��-K�H����<���D�s8?�A�Ό$ӔӸ�W�ꪲ7T/*�z\��/d嵷��%��}o�{��>�U�ͯ5�o_��/��*��B�-�9�K�)n����15XUyfH���?F��#QR9R���# ĝN���$�Z$@U��.R�V�?<�#s�8fu�q�:}=�����x��g�o�\�u%{�� ;�ei\�e�r�<q3�x8�s�l��tgQ��>��"� T� �X��?=�8�%��E'F	0$��$� AC}_'�c�ޒ:\�f/r��}I8����)DLJ֪Z�^N8���z����j�5�p��SK����B~�t�U�7�`�_~P�5=�g�tʒM}k+��IT�h`�s$��X	�.^�{n�xz�g�!	1������Q�= ΢л�o���9#~�J�E��X<�g��k������f��?�+���`�B��h�LB�v^�tp-����גV"�H�2s8�+�d1�<r_��u#X��I��t�!��w1>�-�f��I_f?�,H�ȷM37�bw�o�'�gT��Pњ�a*9�^ZT�ס��<�a�w���`[J����풏G�'��?$��'^t��(��oJ���Aх����P��LL cu�[a%H/�0C;$��_�<ȡ���oT�>�f`�	QQ�9M�V���n��X�S�8 ��j��Q�%p��%��н�(M��aݪ��9�&]�1���A|4}��K�տ 
7(�:���ظ����K��]$������:���t����*)�/ơA.81������������0C��Vm��j�U�wl&1�N��U��Kw�B�C&�eO��<�#���YM![��mו�$1������A��tx�W���]�Nh_�5*���aW�5�~�т���{�a&@�h2]��t��lrq�^j��p�/RrKK5"���"p����a}S�'� ���҄S�suu��J��%�$�O�۝�`�ޛRI~�a1�,WZ��m�����ٱe�f�CNBO���Ъh���K���S H�M/N�<C�G]D�ȇ�%O��B����u�M��(1-S���E�_�4��R���>z�G�YN��NϠa��
ڎ3���;xs�Elu�qh0�t�u��'���j��]�9#��=��A*C��
�^}�*���2(�q��g!�n�mO��g6��4�e*U��T�K���r#m{�QDD,�R�L���b�4Bq�x Q#6�H|<��*Hq�/b����K"���d(�u��A�83���]�(H�F�����j�A��s�D���߀���6%�X����a���J������������C�$0���s�}�s�9+�P\�(c]wr^������]�	���E�����L�{n�-}�������f(~��
�7dm��Z�{��fѭ����r�o�3U�8�ӡ�E��N��b�7|M��Z0F/ �?��C3`�ύ��((
u����9YŸ�Q[��7)���	ٹ{;	x�U�|��9��u��dtę�`����2Z~rȠY�����\e�t>a#������(u�����-���T�;@���?��8�E&����ĭ�1��v��>A�ҒU�md�h۞k��{�Y�F�`�������C��{��E��� 3�a)�ŵ{�����L
:2�j�<C����&��i�LL�x��jBf�A��^���!��fI�T�Wrǌ_�9kLE2�3{��Dy,�G �P~6)�I@W&j�f�_y�nȝ�{�k&��~J�m�5�S��������j��t���E�y*�>��>�������v��@UxI8���-�m��qW��2.����}-xʎ̝��1�#�(�>�%ʈ�,wM��Ts7n���@A�:YF�R�#���k�v�t���s@$GX���	zk����؊i��)�wKA�,þ��E��L��^�v��� ۴�z��_�GGꪡ��\�ţ��%�������H��wHC�<c�\D�i�,�^��A�ͬ
�J���x�:p��>��TR��>n���D<�y��\a�m3@"�4Ic�ݞ9�*���DK$o�0��.�1D��*��c�zu��8K����*z��>s�s�m�JC��N�p��t� �{ŷ?�-YZ�1
��E��۸�a)n�|a�*��BG5UUUCb�1>��>�+�C��:������[���Xm<��.���d�T[��n&�;��Z�m4s�φ;_��B�	.����(_��{*6�@Xǈ�^2����G��/�8l�f&[qZ��9���δ���O�����Ľ/hʩx��V��n�ħШ�o&W�?M:�d�ޒvџ�W����q<��J�p��a!m��({�膇Z����"�Ui�Q��?���T�����s%J`�����~������8�+H��ɮ�{�4?u��:@�����z#74��L�j��}ˌ�%���K����ұ���Di#�^�BK����v���A�"��.~ ]��u���H�$?i� ���互��űcmJF_+ �#�)w߿(mBk�%w�,���l��ƀ1�b�5��.C76�i�n�}�3�އ4�$���� Y
��u��U�|�7��G&ڲњ��JO0�q�:��u��I�A�M���"9;/�?��S��d��dH�Q�U�ݨ�cS��:�ז��N��&YreM�a������W<1����x�TؿwT���]\��Y�#����P[��*�����I�a	�|�l��	�x�N�rh@ZI:����Z&�4�>i81x���&�h����d����D����~(�n��Fs���(q�;�I�*E�ŝ���&��Ǝ)��g$2i�I���ڒ8��n�{��7ԅ�x��}�C��>qZ�N�[;)�y?��q����~ ��%��:��J��.k��c �;����D�u'OL��*�llY\2���n�)\گ7Ƭq�]�yȕ�(ú�q�X>͡��ꂅo9� X?l��^�l�W�q{���[^��,���#��`��,[ӿu��?k`
���ÎU�.7@<���r�̹ȧ��C�#�� K��Ȕ
5����}�/��@Q�w�x��Bf�{�������B��^�BV�q�V�pH�v�#��H��4A\LI��ڤ�n�vE�o�ж<~�N�̓�I�
�a{y�ȃ*hF|�UF�u@g��>$إrW�6���d��i�dQd�����I#�w�ڿ��i�� 8�Y��&�Z`2W}Xy#�����iO-M*����J�/9������`�l)���v��	�%D1?�v����8U� t�K�3�Wb�����;�~t�3�UX&N�������,d�K�
��1�cB�e�k�X�5��=jc;v���gs������꾆0�E�Y��"Z�6C��y�3�yIn�i<7B.���/%~�9bl�P4��&��{�S&e٬`�� C�ؐ|[z����D�_D7��WZh·#�$U@�"f:_R��P�4.��«�Y�6�@]mI�$^��&�v��l�utB���u��`�����;�F�xd+�N�����ݾ�#�D0��N���AY�!Sv;��l7�P �5IϓZ��>�h
-`����/�8�
`��Z`�B>�Ew_Ԑ?�I
^�Ũ+��L�I6��ɪjtm�v��z� �.���F�}�����(L�;5Y����QK�HW=`�_[_;̉|A�L=�̿F;�}�x��y���x\�����C-�� (�;8c��9�4+�� _�0�I�wl:�C���9����_�w���&v���,�3iϝ]}�/�|�%�Z�$�sᐏ�j��7��H;�6D�
�a��3 �x������y�?���g��Oi��N�di-
u\O�dZ�$&���%�<���_f��O��W@�o0	��x���� ;��#�Q�y>���jv��������~W$��"����~����Ӑ�}��HS6(a�����ڟ��i �����xMޡ+��x�<o�B�_4M����o����� ��z]�ב�� �(-<��wZ�%T���I+�e:V�Ч�`[�:S\�6�i>u2�������!�5��� �)�c��ǟgʓ��~��,��#ߪ�29��!�Gx9�~�G\�Edn�`6� p�����YQ�`SE����}�)����.����$G+��-����V��Y�QɅ\�>�c����@�9 �5�f��H�bD��</]p���d�a��i��(h������V;���j��>�MWG)�ȾM�����F��я��N�f8;`7��B'I(ϧ_�����Ti��1
���Z]&�q_���-�=Ԩ/��jOv#+Ȟ�� |[�K/�!���p<�G~�\5�����fZ5:z�����	#h>ŮG٥wFsjݼH��{*�j��	G&��u�2æ�K�p���g���$����/[�lRM ��M��o�K��%ɼ юϋ;,��P��S�����v4�3F�Z����HՉÈF�R!�{f��"��9���k9b<�z��U��|�;R�	�
`�Р,�f�M=;k�ӏ��rk��m�Z�3F_΃�#�PZ���8l5�Qc��BtdY�a�iV��MRoaf0C�
���Pr�1�u���@R��'?L�K���G`����q#7%�O��myǲ�T�H��ꭝ���#�5kI�SQT�+ՎL���n�FCs�����~'R�ml�Ą�
�x��(Ȁ)�	������5~����\k�|�.
�5\q�%�npt���P���4�4����l�u�^o�>�7��e�v}L觓��T�X�r��6�fS�X���C��t=� �V{Mၻ�|Rx�$e��_�	{_�����{(kG��Q8�L��e�x/��g���e�����1��v�A'}�� 3)�{T|(I~�ۑ�S	 ,D��`;ҝ͠�"�h~�c��6�␺"�r�֟��eԏK/̯͊��~��!�b���g n".<���B�4�����{I���N$t5:o�,Ğ+����N���%Ö�9M&㛒�l�g��!���]����{���8rL>�J�4�!�װu� �6+�=<���CBv>�<r�<T{�����cC�rs*\�pX'n៪v4�^.3��K� ̅u="���Jnw��wn* .'ǌ�H��>k }����x5�^��֟N�K҆h7'�zj�20���	J���3Y�V�s�;,�li`d�����+����_2������EQ�;��;���'�<f6�˗����P�yS2�,��6Xo�N�z�Ī��a.R����f ���#>hϞl(#��k q~t��h�H��s����d}G���PLwq?ã����5���l���2���`���>.:�b��ՎPn+#T���\?p�:�����J/H�E5���F�b�Bz�}��������B/)ͪ`M`�3l<��<9���ߥ�� ��۸^�E5���"zp|�L9�*�J��ևL�U�i��1�{���ݣf���?&H�>v����"h��C����r#a61��G9C�0��gґƤ<��Ĕ��"G�AX>�L� �A9(�o�+��2t���B��WF���D-�����]���-&0��۹��Dad���fIO�)�{B	�ZP��ΒT�V�@ඥ���V�7�s���?9#o�҆��#V��F��a��^ť]7��Ǧ�i�t����.��#�v~���>�9Ζ�N�s^t�m��Us��"��S	���n�+G4�pw��ś!\vӼ*�5����Dµ���nھoC�r]�Ti䡙�ږ�PM�^��~���=�-�/��aq�����ѷ|��%9sLb1�k�wTl'l(�X�M!�9�JnI~i%� }�RW[�3]��LL�����o��-,��z��B��� �H���p�#|�&md�k���Đ/��]"I@B0�Έ��L
m�v�����<�^Dn����e
�r�@�<�B���)d�>!V4�`���3���ñ:�ڠȥ�f��5�x1}����#`�+P<�4oNؗ���w��(� ���~��Q΄l|�q����������
�w�Έ�y���\�G���w�X-%�^�FC���Gt��id���*0���l��4�e�bM*+#�9�����B\b��9�5{����D�E�? &����m�'A��k��!|�7�Qhxz���v�c����v�,a]u>��i�94Q��u��j�C"ئ���)��-Hh�0���=�md��i�B{�|�l��zc������	�hr�� ��ܴ��t�ɒ��E���/w��2�[�h���}OLx�:�C�n8��zб�^�n�� .\�	��#RO{nʡb�d����@٨�v�(Z4.�}onG�'N���|�䑜NY�=���u��!�aT�]�p�eHc�M�Mp�����T#�;�Ӟc��z�
D*�#}0�9+\�k��=P�ΒK9=x �c���f���S�7�j�.}�G��0���o���ؐ�C�����wZ���Ձu��`�ڰ3ux�
e��:��1�=H����"3�c;��/A�^��7'a�4��1,r�l��%�j.	��뵢j��1q����HCx�Ƀ|0pPp=K-�b#�}�ZR\5�eҸ��H��k��.��{y�1�v��C��{���7��fDR�ۤ*?�Us.��!�D_����X�����@��-�Nz@�٫�mL�bs5�"%Cޯ�3�
�{�U�@/��l���p�K��#���Q7M��TD�kWY��5��Sv�p{{O�>�r�d}ݺ���c-�nQ��eIiܹƱ�x���$��#}�j..S�Ǫ��6�^AhA���Ε�=��6�w�oQ;tK>������J���D	�����»ГA&�
Wz�?>�
�#w��i9�4el��\7�C�X�uhw������F�>2�7�&��.�����99��m���$-O��K2�����\}��y�&ņ6��)$�?�$v�:��1��[�T�b���<������w�_B+ڦ��l*��QS�d@����{�`G�I�ٿ�����P���Ȣ�MR�i�Ğ���}�q�H��R��j]R"����0N4I`'<Zv�����z�n�rp�������V��Iy'���k�(V��.e������*_`:K�H[״	��ڙ���J�>��cZ�Z�)�uSվ8����}f�`=+׹P�
c�C2e���@��:q�)�C0��鼼��"-�:�Z0;���`I��k���	7�����u��h=a�4�7$��-��!K����&�f;1"���,ˋ��,�p�-�T��0T�=,�V"Vܕ�3&��R�q��Ezx��R�80��+�����ِ�Ԣ�pK|���:�Ն�J�k�Wr�g�S���%9̡o�-�@Kڢ�c��H/�,�pXN9�>. 0��g��i����T�
�ߝ���YOˏ0lf�J���	a��qZ��-zل���;��Ȧ��}��`�������Q,���&|�:l�"���6��t��;�3�PAM̕%�b�+U�M�zh/W5��J6�[S��ڑ�ǔ��|c����O�A~�>�k�9u�*(\ڿ)�v�Ơ.ڑ��e	&n7�ǳ�u�ͪ��Pv%VS�qS;�[�}K�$�����V��9`���Q���-��N�yE�4���0��ޘ����q����g���@h4�o��̑�~d*RZ:�)���
l&���(��ژ�5cb�{�ר�iZ͂���G���%�w{�	������eX���×z���n�@r�z�ӓI�1�(8��$�2�S�-.e�����7eT�F��@j�/yJ�TWLr-���*#ޕ�0��܈A���8�8�.���e�W�߁k+f��M}"~~ˮy����v����8�IH#ƍ���~T���un�f�>��ܱ�:���
3��@$6N����nu���B�z����<w���9��J]�~:��H�ҍk��_�v�Z�k�4�<��c���B�ȫ�OR�Z������>�f��qK@bk]v1�]�CBʪ�9ӻ���e`R��M-&��m�b�V\���� Vm��R�Gj@ԃ��A٢�C����Ps
���k8�S�NZ����o/2����OV��|����/�mE��m�p���v~I��G��߉�/������#5�틘Y����D�pVv ��N�1�6�LC�o���Ў����..eT�;� ��A=����^5l�'��P��]v���Bٱ�?���0sF,h,q}�D�����f�њ����E0�����)����y^Eh-��@�+E4L�fDV�#g� �?�r�9_���0TH����4Üs���EXJ����hK�'�:x����2$7��z<��5J�#$��kN9���T~��w!�a����k�3�s�&^��o ��z� e�~
��-Yp�[���Sh����^���X�[:��$B���{����v�M<��%��[���='B(������\?�kMA�������3��cB�0�/Bj4B�j����E������1Ϻ�9�ؽ�	����M4����M��O^�`�`�7X��#N{��LG}!��)�[骧N�SN���]]�_����_Q���H=3����kX�f�V�!rWVZ�U��ghÔ�t���f҅�/C�a�_�I�����tlYQ'ʠ��
�\]?ŭ��0��9�k,�n�ӱ���5l��
{8�KW|ƀ�T�����F��?��ip�U�x�"~n�Gn)�ӴR7�/a��� 8���1��9X��i<�!�#e��!���ѳ�wh]����^��ܽ:w ����oH��.��<��=鬪m���U�*?CWb�lA�1����YDDM���|S�~�b	��2��,�*a��!���=?ς�T���k���OI!��1�ױ5.�6��я�C,"��M��&ɀ췂����v>R?�����x��<�u�.�� ~O��$<z7Ӆ���ЌOl�Iz�wׁGXv�ˀ�G�GE)��q���_�&��O5��CW6[�r����"n{^@���%$��v1gb��!7�輟8�
X�zR�AG��g��S���ق�d8�QOr�u��p#�G���a4�0��&"��4dӕ�����p��Em�8�U���_���]�nѥ(�aKo�w�a�G%�s�6]F�3R��&�:��U}�B������䙷s|��rk�W��Aur��f0R$�h�~��]�B�Q���ŧ��I�:��f����M�_^8&���~�4ih�|\�k�:cN�^U�<����G�^�k\���{�=�����h��P;-�:�'�OF�H&]ע���o��n]/�Tn�m"O�wS����V���1��j�K����u��/�{z��3�$���� 8�
[��ۘ�O�>���$�Q����x��ўȂE�.e'P�1�&���|;��	�B�;��J���~|�&�0_�1��GfHeJsB�,eY��#�����Ig��f:���Ԭ�~S'��^Rf}���y��y/ë��_��j=)����3I-��j���P$�j;+���;�yZ���4/��GC˝�Bw�{Qz�2����n�+�hD��\J���<x&u0�#H�"O���Bj��)�?�����)h�w�fQ<��G�YF����l��j>�����/�^�k�L~�����i�Y�%���X�
�c0�N]݀Bƀa�},�\�?q��S2�/H�0���&��dj��v��$�Q����D zjPhx�~n�iOcO�..��U�R�e�T�8�В��x�+�k�4���3��Bq�{�\���_�S��-�+`En$v�?�7�dP��gs��68�_�|E�e�3~���X.��g�S����f�%l��W�h�Sysk��q���p�1�$к�4?s���Y6�w��������x3���3-���'Tq���8R�uo׊ځ9��(�����9��J��&%�,�J����H��&�_#�EF���V"����F��*,?�ܓ;Թ�QG1CD�����/�43�9~��Y<2G�n��[�=h���y>�
���D�,��z<�xv!~�X�g����ǖ�0-����g�")���+�Bʓ!EOHZ�ۇ�~����X� ԇ-B��4����//�o��+k��Єq�����iǴ�?/|$�g��R��R�ڢ%"�����f`��Y���$p.�S��sLY�z�1[�e��c�U�H{��/��jb_?����X��&� �`k���^3$�����$ݓJ��tO͈̓{�Q������a�r��}�;�x�4�	�CWT��VX�"�62H0�B�э=5�p���(O�"c�N��RⱲ$E@���`���e7I���ٷ���i����y!��igǃO7T}�)��|H85'�Q�\��rSн�O9�~���X⇨�y��U�E�q���֭��I��Ί���Ζ=}S
�_�(~��j�U.!��Np�i�ֶ1��h��Ԏ�,��b>!���fIQ��_W��Ё��FA�6�f~�1k\�WZ�*��:��%��G�|E��bxY_�3Nn�OKx����d^쉧oV6��!��8�U/J�V����	G��̧�~�#Ml�
��T�9o�6����4�.&�Cq�Wf���c3L���`kOcG���x�h�X �� ).^\�����n%}6��}�*|�d�����In���c�)J�}���K8U��++�!�ns[2z$[�ikG����oІ.�D����G�uM��(^Q������)��d����W��]��:�^��ԿY�����N�\|hJ��.���)�o�֨ϐ�g\l2����9�����(&,�_ĵy�#ay:t�z�z�{�e1�¡�|���Y�do��Jgŉ�N_^!d
�\�}�um~_l�.3��_�q���u;���p	U�q�+�hd�;�0�%��{ڪ��}Ÿ��Hg��ZH_J�f����5v_�UKu��
>Bv���2���<��(�p���	�{o8�Ў��4���q��i2Q��6 ����v
��/�e���9���'_΋�Ar�l�x�v��J�:^���.kL��P�㜪ٕ������`l��/�;��n{z�CF���0=���V��e
���;��Z���K#E)����s�����G��Pe�hk�>���LCԬ2��#�p~���$p��P�݂#���>���Х
�$�U ,ܜtQ�ʋ��w�5�s�~�ɧ�l{�XZ�\u!���HgJ��v���M$o)eR#�Nɢ�,�D�f0X� ��%�Hq�ay�����O��f �k�׶�t��N�=Ц\hs�p6��$���_�JO@�����a yӭ����6�R>��&c��>$4ս�����
�ߠ�U8~K��Amb�Ϡj/���9�S��FS����Qi":R4�Ssjgϯ��?`<�S��A�`�U��M�MR��t�_~�n�a�h ������Ʊ�9e�P� �>�9�S,�8��đ���ަ	T��G�t���Vz*A�2M%v���Br�8M_�E��-8�p���=�$a�f����lo�j���^�Fc����o;p��J��"��p�iӎf+f�~�s)���\�S�A�i�Nt%��l0���U�޲�Io�c�b"��Y댃~�j�d��In�D?:��o\_
�x>Z��y�qf���]�,��c����[����v�zg�+JZK�B�}�D9��@2�"Vfw��D�%�Y�T&�a��M�&�=U�ͮ�������(�EJ�p�w([���������k��1�B����#�@fd]�`����}���3t��ű����E��D|�y�O�� ��N�{=PW&XM��S��v�*rm�S��9���?���s?��u#S�������-�(�J������?pIۮ#���8�n|}:�ɼ�zCy��Ʊj�x�����G$��ި�T��x
x��F�+�
.3���g!9p %�=۝��V;�Aї��g��7��:��ۄ��*���5�>f��"
뽩h�G�H,�y��9�-��7O���P����\�Š�L:�N�Z��Yՙj�L��ة@=�ݸ�hִ}�`��|ߌ��ăK�D��M.�4�H��ɽ:�.Ε��O��Iu���
Au�b�Å�M~��?�}��7h=#����2ul��`�#4�j�,��:[�&-��w2��`�2xg��K��?��
c2��=/6%���B��bs)R`���da7��ZN� v$'�E�����=PR7<{>���j�3�Ⱜ���T��'}˚��G֌*����H�.���M�֖Rvʃ���dP���s���ɝ>�M
,������#~m`X���>�mޡr�&է�w*����u��~�5BU"���`�,�^=�m��pԃ�9��U%���$P���gQ�fL'�M�_�+�&���<��]V$67�S��Lo,v2k6���3Ԉ�",a��q ����g+�I��}�,���VT8���Z��/��0�C�L��i�_�����:=���vj��i'�<���<*lr;+�ON���������nK�
+I�E�����E�����bQ���q�GG�������13�Z۟�w5��`����_��>D�'�~w~çt�?x>�T�8)�*Pj�󉌽��a��V�cІ1��jm��G�t@����vQқ�K���i���:����� /�G~�S|�39{��e ���sHC�6�h7FC�$za�t� q5H|7ҍD���WI��,�$韢���!T�0}�_�I�^<�����*�T�r���4fk�Ys���͠f�	�S^�V"���o5n�?A1[��AD�(r�"�~�W.[�%���ϱ���+����N��ձ��6B~.�|�9Ub�#;�5�n�\����ɮ[��M+2m����g���4�t;H�L�E?����Sm�c�|�����P���ӧ!z�+t��I ߵ���dS���[]�)���.C���j#���~Jt�_��
�(�w$eUd�.0�-z��휛�a1�G��~�S��]�a�K飚FM���6_����|�]�����k0����v�������`�~�$xOx7
ݱ����>~T5��8�=p�����c��e�ʼ2*W�P�ynO 1}�#N�{ք�elTB�M1v����8>�R$W\!ɲ�k�@�% �ֈ2�=6ma��'^��8os�b�Hp�呱��7#��&��ýQ�����X�i�8/����7�PY��̓�0�Qj ����Ψ(��c���+�[�%�־��Hd��2�uЧ��cKN��9��R�)�
LQB>;ʷk��5���"I��o�����6&"�]���s;��{Q0	������"��dEصAS���	��>��,�E)�]�N�b��1���nO�#2eEDJ��(��,<��W�ic
U��U@�7����w>�Uq����[kZ(�LL�#�����F/0[��Y�dA�����iP� ��-؇)X��3�U�O:"�����(s�R��>�r�C��>Jp?��0Q2���ll&C�� )��|�o�u�
cF�'�A��a�K��
�6{(�-1M BR,�>�3
5�%����d"�}�w���H��6���%C����c2r}ѐmN_��I��Ň8#֊F���¦r��%�.���K�FpK׭�����Z�XzY
.^��wKj�n���������lF� +-��ô����% ���@|����Gg�@��D�\��)&�n�&M�u��p�-ԡ�: ���$2���Ar΄9�ث�q�*�aJ�M3D� �n{�>؏b���j �~8���C>�BXr_�s���	�z�5	ԕ��d����H����+�i-\��l����t�d%�l\�'���~�̟q�`���_�|����[ȷO����}sX���زK#T=�赀@�r�,�r��?�Ӝ<"�j<k�H���y�{�P~#��ev������� �W%#g��A?d�i{no����yIy��u�*��Rg���?����`(k�d��=l�����>��l�Q��c��Y^��p��ЕZrc�JW�~�ˀ=�o3���?IQ���T��Җg��S!�eh���dܣ�Р6�c}v"��W�5Y�Q�,�xI���YN��'��o O��ii�����:}����(���oA�����[�QD
�E&��͆@��A����A�`�d�kQ��j��X"x����?/��n����Qf�o�C���H�9�5Kw ʔx$��Vt2�qg�]&lj�xhU�����h�Ǎd�6�/����ȉP�v�H1���My)���Ϳ�ۅ���c�c�"��F�?��Ĩ��c��� "�h���д�kF0��iջP�&�**_�u���?[P^��<M�������)�,����&�?�ɭ��A�.7؏��,��]�s��	�t*OTav�����6�n��ul�Nh3C D�ϴ�0ݶk@G�M'n�I���4q%lhqL?|�F��=��|ߒ�l�x�tsX����%��Q�W3kY:
3½�����!���������u΍S$cz9o#h!ޯ.bY�}��Ź5���[�,[��+���0����F�H8����z9Ń���e�|�VƂ}3��h۾ /FؽQ������{e������0ϋ�"T����JB�m.>A�NG@��W׮]���q�IL�`F�<|!����Ȃ�t74{?�:�&G�9)Ĥx�����;��"p��Ӵ�x��x8*���M?q��e!몁Q-��
~Ќo���i�wvhMY�����ҳ/���Z˃諊�	%ؙ�Ś�)�����nf��lU�W���~O�������6�e��ZPP��b�EkĤ�	.��e
���|�EQ���g�a���9� ���0�|P�1�&&1�(�Q�~>'����X�8F�3_P���&K�E��P��6�5\S�@��"�D�h1�ފ軍���4%����7H�yQ�$��U�Sxc����9Nv�>F��_CG��[�ҧ�h>-���J4��&!P�Ao���C�@��~y�!�ڑ>�В)�雺�^��K�(T���Є�XA�rp����ё#��z2����^��B��܂�P�馝yS7�l6�#O�Y� �6��#,{'M��Yݡ���o	�/�z�/*���3��d0a���_ԧ8�a 4J�W8Y�Y86ĶJMኁ[¯[�9�0p+�r�����x�(�Q���~� �]]�&@�f0O��!D���3�\�%:�;ھ�vV�H=�
t���ƹ߄��u=vW����E
 �!|�. ��/hyR2l���Zi�د�� ��7Y��5`�=�q]~�T@p�H\K��f�x@�e-���ey�DVY4��vhdՍ���QQ��ǣ�֟H���	����%�q7[%� pw�ݯ(�&����0]Kf⳪F ��A�&6�.�ių��<6V���ɛ��r�~;�i��
����U����)��ȟ���%�����FZs r��ZƠ ��X@`�Ґ���<%�����V����h�=<-}m ��?�z���w̽��0�� ȫс.޸�s2p�s��K���y�������]S�Ϣ��J��"Vr�*�Q?�2�x�R<��\��L�SiC��#��^N��2n���M��+���=p)'�J�<�X����w49��a&UR�6���)��_0:IP/{�
���@�|`.��9�kH8��~#,���^,rT�K,�k�m�0�q%�u���k�S��ާb|��g���;Yr�w<��ܥJ�/m�WT]�����~b�鏣�D���|~|;[���������?�b���&��5���i�_�F���z��cm���RG�}ʴ ���۰cfS�gE�_9����H��-ǎLft�<�ٳs���c�Z��� 5�#�$b�o�K��'�s�$+����ysL���.�O�J�$�0�7������*��ͥ���Q���'ef��2n��6.�����M�1���r��?�)D\�@j� � ��X{5�HD �٘�{�1�ɠ�p6Զ��"�aUHʹ��u��?���\�r�ZIRܿR��b7�͠F��F��e��tIpy�<�G��8���i�`S+�V�ť����g�Է��=َ�,�A�we��(�R�d�V���I���0�Sq��~�|�	<1�G�?����6A�#��T�f��o�ZJ���ѝ�R��x�tU�a>��Ӽ�?.��a6.^����8)��6�%uC��rYm��������@� !f�,~,he�������n��<�ZP�Fmn�vf�<�J��4s�� |{>� �>z��3ʇg�kUβ��<��Q�0d����@H I�>f��s��$Qw����p�nV۟��#
�h�̈́�dj%&KD�f��P��%����j=���tr��^���4���[�>vEd�J��2���u�G��{e�'��Q��r��ex�aE�#���J,�	ތ���/c�Z�E����( ,�ae����$�b�����;���F��gYIAZ�]}edLR3��q�j8S��kw-^1�k5�v�ꦉ� !X�9��fN�6�!2�q�e�4�.I��/I�3�[G�/�"���	e�X��X�j�3��h�2�e99S��9:���#��0І�!�g`��2���9a��\�Q(�uE��{m�Cɔ��v�Z[\�]���w��ǳ��B��Qu���d�G �#d��VK~e�ۧ.>Q�qCB�e�+�v�t:�}\��E��:�����%�t�z:���t��@T�a��]գCة��l|��~��y��Ӧ߱���D@���P$�v=J����j�bO�N�Z��)�#��B�,��!�f���QQ~o��<h\u*v��"�_�[n��Sy�(�
��eJ5V���$O�B�X���a�(�٦�T�-�>�qX ���}��������R,�x=?�#�O�����l�55:#D����A�\�-����],�%�ʦ
K�|`0X���HƗu ]w�6�u��\��I*����G��m�c}���$H/�u6\ t�x�������:S:�2v	�޻���e�v�n)�֣�B�8yJ�O��0��D�Y�	��`��&�ҹ{v̬�9+K;B�����k[��M��8���G	�t���2�Q+(ox�pm��vBg�����Fq#�(���N�����c�	��R�n�]L=w	,ґ��(�F	V�/�X �#K���f��~BH��w�M��u�� �߻�o�+�al�*	J���. �?�3k��B�[�{�'�\�n���BE0)Z�{�b��S�-}>3S���&2%�'�&�%/(I0s�+g;�NB���o�%�i}m��S��Lܶ�N	���U�w��n=6ۭv偦�� ���� �1�jc������vH��B繵�����ȜT��ټ���a�E enB����Cm�ޘq�8U���7ϟ�:���.^����t��ˢ�#w���;��* ��CA#�m��cs�"�1*��Z�>�}Q�s��u�'-+���PA��nΚJ��يct������a<Dw��:'Va��ݥ��F�����A�a�*��=L��� �KQ�Kt�?j����6�I�%F2��!I���c*�eoOW��{	����'EALf�B/�f���������>P~�1�L�d��G��^�{/c��A��$*��ۃޭ���=7��q�������M�Ka>��"s�݂�o`����w����(`��+F����7l�"	v`?� �D�E-b�Ǫ���!���W4�Byp=�bߩ�O7V\�[��2sI ���@@�����aKJ������;QC!������k�w�MC�_�Zvo(�$�Rj�쵒�7Л[#c�-���4��r2?_��sː�U滜m���ǣ�m���o�R��/̈́�la����� 7P[�f5ݢ'���a}�������s���ۜ�&(��6�8.ۈ�u�N��4����x�	@u脮��]�*946{9Ӆ�M��F�l����1���+�>�`1 f����������ձ�h�47�(���?ng�XN�y���D����{`�s�$t�n�M� ?5�>S�pg�h"�	���[ \�g_��h�x;M*[������!�6���c�|�<�h��Ix��w���<���C�
��襡+7�
��5h�GR�?�)�E�7B�����9�k���(3��M���ή����(e�0�����E��A>������Aߤ@>�;?��ѽl�8�D�O�>dADa��̦zw)�w��]WO��I�}��Љ!�ëX���*�ǄK��/��K}|�7����P<#�[���Z���&���,����1�p��yԼ���s���l[���ɟ��ٳ�ռ�����]+_���^\<�RBVo�O�դ��&Z��'kɩVP�ԕ�$C����YC��(ġgq�Y�R��g��Л��h����0S@�T�J@JGs�-֞ɇ�I%OZ ��/�y?9F|���C7�ʆ�1a[\=5)KmDW�����|� �I�� �ѫ#�'KS�I,��xz�0{X[��/M����z����&�r,HC��r��BkSŮ
xZQ��+ړe��>����wK�l~���<-L��{0��Yj��P��R�U�L��M��I|���Cϸ�-�ˎ�%8�<�;�u_�8]�޹b�nP����>3U|�a�����B��L��>�U�q �B�&�rāt�x�	������`L�@��U(�q�{�1�*{G����g~U�~, ��Z�! N�_yp̖�|B�{�:��_���{?�Ԥ}tŌ�P��%56�B�lT�� ������GqNs$֢���H٩\���Qɳ�ٮ71�����9�VY�wӍ�NA!��}��}������f���p�Wc֢z��'�3��U
����w�P��9!�,���ɤ�ڊ��m|G�%�p�mx�8��]x����/ʒ��)ڴ휏1kI�!�i�l��I�b���do���Ö�Q�%��W�!��Ӎp{�g�-@0�;�A0��P.�ie`.1B���H�}�B������q�z��(C!qUEΛD_��^���޳�����;�J��WA�[Ɏ�t>x��� �+��T8AGFEm؉l^�G���_��(ħ`�k��R���[`�l*t�,�}�����ڜ���m�2����3�I�T=9m��Y�Ghۇ�c�d���:���e%q��JQsM�KG�kV���_x��O��xY;Q���
S�cӊ���(.*Zke�W�_�e�I7�"1 0,�Y��R����3�\������@a-��¶��X���4휡��4I>�ޜ`hABaT����f�_�	�P���$�9[�O���!�7�����rex���N(�{ކ�)��Uh m��QTU��&�\�ipr}�R]>,�z�{��h�F�͘��"��j�����$�[�pُ�ICc�{<������>":�x<�	C��\t��Y1�9��ބC="`��'Y�b��#��'%�5�=j��a�:p0���`�.z���k�A��v�����v�1.��>��©!/$��\����툖�9u�A�j�6�a�w-�1��KW��p������ܪ�`N��H��4�BFLZ;�q~���t���H�Q����7� �(1�-�*�AQZ_��9|�[<����nKZ�?"�^J��k�(���|��`�\ͤ$�Լv���kK*u��t1h���cf��;�E�����GA�*A7/X	��2j22n���--�~D�LM���P��$.+6v�0�S�&xeƫ����z��0��𼶗�������#�]+K!�� �Y���^�8 bn�=�������d��F-ӵ�<}<�+߻����1ʛX5�:�x��W!h|u���M�J�f��w�&h�����9���}��O*��W:��5�$�<>Gݗd�|�\��4G�J;l��w��J��c�
h&���V1B"ו�V�������/�sԏ>�&�cO��%(��'D�(|0n>��M�1����4Z;������Zy(�� ���0?��B������Iu�J7�������E�urS�E-��d\љ�P�C1|$�֘~�eg���Blǐ�ގ�!����2�� ��O�{��2w�c��'j�P��f�ԫ��C�y��b�%3��b䴩�򵤆U�:���̳������9'kx�L�B����r�X�Rq����E`4��|��A<�hd���	�;���w��w)#}~(9AnrG��nI@
�>r'��C���o����i2
���|���H�� �F��Iٯ�|�#��6�	x�fb�iG����m1'�;)h����=��d�-=I���76d�37��_�-J��X�g���V�r8�T�8?�G<zw�UE������+t�&�Q��y���.>A��@��s� �ˌ�~I><Ь$À_�"ܳ-���B^��V��2Ǚ�M���~�ˋt.��UQ@=�9��&9[D#w2ߜhgX	��3K��A47F󁊄Ig~-��}oM��YY�Y�.���(��X-(�\�+ps������Q��tT"ț�m��A��? 0�ۃ��A��PH�%��6�
��,�/B�V�JB(�Zv�����h7�R�F8��<T#j�LӒ��0&���y^e
x��1%��ʎY.\_��@�"�r}+�E�#�,����?	���Ëw�!��_o2�'#wb$L������� ��;���@���w22�%BS��`���[���.BAaYP���ll��>!Y�p`Kq�q�F%"g��0��B�8��_'�ql� ,п�&5������Nr�G���������-�2��`�K���yA�.�K��)�i�#��U];NU{��J����1f(����:KР��=1�ܾ�e0��HU~����PKB��|Bǘ��?��*�.38qn$�q���F�����}���rb��_�B�ϒh_���DX�&1k��P�j"��0e����7�-G�ȾN�O�:��A��%=�Z�.�<��}vJ���I�[O"����$4q] .��X	�ܬ�*G�fei>-�q��[�
x<X?�|u޴�{�ōl��Y���C��9D�]3��R�����g��	51V�)�G�.
�$�z�%^��W-#azb6pҺ�L���υ<k~�>�ř��5ĳa���	C�Fʊ�V�B24�s�{z
��I��pǠ��
4ι8L2�ཥU���,��i����V,M�wMP�1��r	q:Hh�D	� ��h7��)���P5uB������V�Z9���h`{,�����o��v�ۍطx����̫%tFiǾQeae�{y�|=���ð��6�=F�C*�6�\ͭ�@��M2�]fb��J�+vxR� ��gS�Y���*�E9��ny��n态�ѥ ����v��_�����P�}]�[�MV@u��N.Ԓ�����da�<M���bQ R?�iw3�D-��r����7�� ��JJ,,�Q��B��{����
Q3=�T�W>��R��>�HRv�}�5q�˃��K�{1�@�T�C��Nn|ͤ����@o�7 ���Y�r�:� �~l�=5\����i�'G�S�xx�+��]�W���]� �������>�S'�)����xZ����Q���餒�8�:ü�3�S����@�_q���(�,8�-���"������pL��0\qqД�R�G{r���FO�,ǃ!x���ɲ��_�"�`Í����~�H3��,#y�q��mI�ވt2aa��ǻ8D���,]x�*���*B��-�rJɓ���l牊 5޸��P&�U �{ձ�lH�p2�L�s'����׈�k8ZV���頝:��3#����D�l�;$�h�:��_��'�L�(E�^�bo[��ny��2P��\h�v���q�v��
�ǊA��:8�8qe`�i�5a��s���\�=���`�|s������+����M�q+D��ղғ����i�S#��)VD�!�P�Fu��R(�2l'�������4�!�Ӥ� S��Oj�UT_�t���&�4l�B1	�hC�U�ng`��+���XO��^��VgN?)��W3i+����R���h|c_� ��@c��"�4!�����P��m
T�#��Gȹo8�̼o���^N��4��=P�Y'sG��-d=��rW��g+�w�)�׺W�Ӓ%@>�u�5��x�Ͱt��7�%�&)R�,�N�Pe���.i�͕��6��<Or�op,�f�7��1��O,oY�v��J�'�].v�Ĭ�t�AWf����c��lV=T��.�T\(�W�u���K�M��}��\�?�PB'�^P
\10�]���艂�A��Gk0��@dm���V<���i���,:��L�Z�N�B�W�c��aO�[��6e��Ǔq���.�˽���f�R�S�����.9�u�mr�R�0��R:?u޶X$P4A��K����Y��o��z�!F�o+�����d(*k�2]����c]�iY���u��HZ7*뫕��qǧai�7A�-�,����)YYE��tZ֬��S�=i�A/ҧ���n�A�T#g��\:v%����T�Yh	�����f���¥Wߊ;�ݵ���;���V�ŗc�����fDy#�<7����s�U�%��	S���r�� �*�����
3�ޞ���s$���<�ͨ  g1J㧸�^pb��`������Bol{��َJ�zBa�_n�{q�x}W��;�k���?sy��zC(/��5��H5��e�B�cFf�)�o,�M�-����2MQ���o�a8�N�c8*f6���oz�-�d��v<��j���[Q�_�9��.��IP4�^��5(q'�b�7T�]���y�K�(��ׅ��#��%��iKq*�(��Ŗ�f��-	��}�1RJ]��1B.�'`�Y�o�:�,��xN�X�����m�:�� ⃡���<�U#��|�ay�@/�k,�L��e^���@�+@#�v=�\��X���R7>@�	�����ЗB�q��	�1J�8��0]]!�>��.t h������ I�-������AӤ���X�7�8�;8=τ����GqvsY@�{��Ę��S"]�ʄ��uJ���<�����(U�|Y��pk&�Z��G<)��T�$d�18H���d��A58ki���.?d�c�K�2mA�d��thg�oe.7S�H�V�E[�>�W|���~��N>�J�,�Q����N$fE�����0��''�Vt�xW�iA�~��Ӗ�Z��i��SS�[XQ��Sq}n�Bh�9���]���ah�&�sQc7iA�e���3af��L����lҲ��W-y睨ʰ�e�5��dX�m����m����̅�J6��.%d"���;X�����	ό��g���#�6WVIR�J������=��F�mJ�}W���>r�%�ka2J�>A�H�t�UuuW�,*��
h�K��p���Nc����cPm�h�{����z�k�(�K��B��+FA��]8�\3<g~��&�{m��=�$U�����{e�ݵm<P^P-��/p�]x�6_�k���9��M����|P�e2Fi��\��`�L���'L��r�E|:'����u�`0׊����D�z�:���eŕ�Q�=gx̽��	�1#�u�l ����qV=O<�9�\G<���@�u�>j*v=������[��	~c򽢹���XE�5 ����÷&�$��D�'�BO�=5a�rNE��{��vy=��z>����-E��mP��lS�my鮯	�vi�	���3�iO�^�Ij���R(YW��[���+���Z�9Mؐ�^����$�x�Q���U��d����6�P�f�$^z��\�F�����,:T"���xR�gI0�	�
$a%�g�F��%�ˢ�e7 ���3�����[U������D�#�!�'y4�:���+���� ��i���e��	l�E*
��M��O�h#N�s��'l�����L)�z��L�A�Ҫ�*�/[� g������a���t�6���L�޵�g(燩՞��G�+_�t�p�~A[��P6��1c�rIJ����Yε�a�eK��5ٗtׯ�΂�؂��s�ݯ@s.��W߳���|BߴeHBbvb�
�ިz��ß$� q���h�t'D>�V��ct��XeI �fq&��q��]O�E��@:O{���������7LN�4*܇Jb��/�Id� ru��$6�-N�f��a+9W�~S�z����7a@+��1����V]W��Uܲ4�w��T}:8�%42T��6�Mϣ����2R��G(WxM�.%�ns�؆�� ��ڀg��[�2y8寓�6�0-��@Ɏ� ���	�F�]�J.W�W9�n��S�ł�01ҺZCHY�o�C�.A,�K*3�~�����Vp/���p�O�'QB/9�I�MB��g#�4�>��ik:��I���H~�<���>w��B@�G��5�4��l(z���MXy��Ѭ\�&\�Au����هY'��/�	�-Ugƨ%<��eR��Ώd��$�q�d#��FB���6&�!o�ϋ�b.j�X�v�τ��g~d�}*�F��O��C��1�ڀvOЎ�;3� �����cy[_���o������)8�N)��v*�|�I�޻[r��2B���(�]4s+}f���oğa�t��6�Z	�DPj/���J�58�j��-~���Ӭ��<P(��Ͳ�!'�	'��"e���-/
����I��JEWv��@�����ꨕr �?Ku�Lq��� ^�]�\�^�dz�0�KOB�
�o������h�tk#���*�W�ju�l�b��\\M�f�臨K�.���DYt��2����m^�^�J�7F�
g	7hu���~_��2�){��3�1�D�?�Z�:Ehʀۙ9e��.#����Q�
Д�$�y0(n �����'-�9{t�����G��{pK�H�ϓ>�����9Mg͢�+=��,��=0&���J���|�~�rx=�9U&�'� �;��0�(������d��3��+9S�N���92/������[Kp!~�I��=Rf8�xW�$,蟽�h[�vR �8b���o�=�H�ռ�(�A7��JT'��KLE�>��9�#�nT��VW4Y���h�]s ����T}�Pw��Y��\���cį����B$+�&x����jF]�%B�:~�ӧjg����j Q��y9�g�K�o~�&��F�W ���R9��0����?IVϰ�rȜ4.�Z�M�2�@ߕ�+�r��̶H��*�����`��d��d�o ID=�M�,W���J�%K��*��"�q������Yz���Kgu���k�_S�e��94��䊓A��D5`����m��P=�ӰF���@��f$�������F+�q��Q׼��vU��H�^a�t��n���`-�������jx�&����l<��R�\>�D�I<���`�~� c^R��{zg*"�����i�.j����׳��)�$�Ǭ��޻�p����Ά���@Ŧ_�9�uy�G�"s��|��H�%F�?R�@%�a�VJU���1�����]��Y�D���L�r�]���g�6�UR\`����!��&��	���v�TqȲ_Έ/��L����pɱP`ѽ�� �'崚���-8w��1��=}i��+�����^�kNo\҄�ß�]���2�t9z�O\"u�8�X��1��V^�_[V��Q�ޅ�g�3S0 �;���>,e_��ZRO�%���.#s��?���}B�Ħ$x0�� �x?�I�E�k�0�B��/��x��on��#3lk2v�Z0 �rꓺ.� j"L����y�۫�>{�Z {�r&~aD����9AkH��!��k-g7���y�8��I����,i�
Y�^�@��"�no<J^E<.w�h'�]���j��d�g�ie���&���Ie�Ϸӯ�*`�+{Q���vS�8���G+���;�I\w�=G�0ctN|��r�)!�Z<���O��l�1ӫ,�7�+��� �zzB�?��B�	�0~�$@�}�,���X{��Ȯ��*�)�ԪH��P2 J��`^�;p�}�o�3�1�{���>�jq-iU���L;���>L���R�#<�E�p�N�k&v�Jό:�;���FU�,'��5�?b2&K����6,��%�D�e"�g��Q��-yϊmz����B$�} �R���4|,�@t�&B�F6�t�v�O_y��*�IH�u$"~���[W%�������y��w�A����i�ލ�j���h5z�
�\��a����CӃ��nn$��w?To;=iأJR�Z$��E����m�D
�F��R.�泱�26���@�Q����;|U�7��&5e ���h��-K�]c0Wh�F�*턭��M���l]4ԃ3�C8���M��c��S�u�?.�!j��� F�
�q�TUӶ����w�?,��ia�����(d�r�<�u�׭R�v�O0x�������)�ة���4�ɽ��	r�8�/�v�,���c�e����

��\{,9�l)�1	x����NNtH�4 =��������A)��E����K�v�>u�q{	�v&o�����2����E����I-0�?�2`3X���L��gkm�W^����a(��ʨ���X��(����Q/�4f5�O���i�Hء��I�`2������o�~��6�*�2���������������gQX����|'�⥔��b����n���(��[�|l4�Ӻc���I0"y���}ؿ�F,�u^M�l1���W Ė)��`f�OّJe�ڨQ6�� F�G�_9	�z�:���9�'�S�h�
J&�2�����3�|A�e\��>s�y�{�����X����"�j��cD輸(X�7��_�z�lwΆK��9�?���0^:q�ч"E��j`[N���x_��C��*jg�ҌH���������{Nx�k=�,OT̮�!,��$�D�fN�h�;e֌�\#x	N�P@G�eJc�<��;�v	�3	�I���*�to��IQ;�,���b��xm���{�%j��̳��<h����پLwln��96)�Pyǣn\0�x��n���7s� u�35���6KZ�� ��h��D<,W?�;�gaC?���@M0���#��LD�;`%�5��]mYV�ĺ��~.���~❫�x�,���(�����*��a7��6�yy��sKR[�o�n��~ƈ
�A�aRz�q|�8M^�v��)C����[k�W�$*���쬸�՚C�;=s�"
{TҌ$&ďO��N�5��F�B����Y`�7�Jr>�ǳs���uE	N��:���*f.S{L|V���8��Bsi��Mp��߈�J�Mu��Sh�A91
�u��-��2�A�K��r�	L8��l^��,˶gj~��μ��@���N�c�-{��^��H'�J�]����P��㸤U�#GP�����^+�v+���/�t�����PLX΃���@�?�O�[#�D��SW-������o7Ƚ!��?i��
�me�}���V|���g�P��N��E�ej��(�i��_;κJ�k% ��<����+�Kv���u�9����9k�m�'Ф�-���y�}u]0!s�L=��[�e�5eTeA�j���,+as�3�k�8/2�ݶ�c��n(�s-r>93�S	3X lb�nh/�c&.~�7�����/k�D��;b)�$��w�CΜ*�B�w`Y�K�F� a�"�n���Q^���x���u^R쒁�B0w���6��W�[#3��	 ��MF�zƅ�����W=)��u |K~��Y�D_�?-������+�;�FP�?��	ޚn���8�K�S^e����<����2x]�F��V� 
�$�e��`�,!G���X�$9��=lO����N�YZ'pv�H>s�W	/�mk�A�V�7��C�*��@��#�x9!�Y�W;��ij��v=XJ��r�,R7jӜ�bx�� �4���E�������Th�U\��U��.�4��<	Ȭ/�S�=��*���R=_��Ҙ8�%VZ޳�������RaU��)v�)\8n�|��7�A׹���>Bf�ᯣOt�:f6�������=b$Q�����dd"�/�-��A�R�ib-!TD��vN^4n�9*c%?�u1��L�˃Bo�1!���m�E�Ω�e�~c��H�����Z.B=L�.
{,s����a!�\�x����Z���c��{0�ӆ�P(ȟ�y��Sτ�{W!%��Ѵ�#�!�k�f9t6	��%fj�3��s����.�Q%���c.�0|DgV<T1���Z�^�u~�H�3pF��=A٨8�k1�V�.l|�4³��"N];s���>ĸ��ѽ�ts�|��3!���d��S/�?jG��@a��c��;pNG�X�>P2w���R�3�`v��o�~[x��!�����Pהt�N?�q��<3�)�e�/�Z�s���'�&q�6����:���x4�I��O=�1���svo�|B��'Tjm��s�8i�!�t+���0R�<z�}[���k�U��2z�:66_��ʝֹ�&p�oDhsq��K�&`֗Q������QkJc�wXYk��Up\��
 �S�����Jx�>���["���&�A�.��G��*�BD�͛-������/�� չz�;jM,���G!�T%W�O��C��I�ʦ��o*	j5+��gyke��P���	JS�f������?T��m��_ @~u���|�z,=��h�˥]��)����)���������{f�fh�e}��t
��x�7V�)��;v�vq1fV���;����Q6��Mwy�P�]G1y]yZm�U)f<l�N�a�kL���� �f�x3ə|��}�H�,/�+H�"���I���@�4�+ĠV� ��;rdv�]���D�){��!�o#���GY3�Xs�p�N���݂%�ª	��b	Tq��A; 4��b}nC�E����,��Vqa�A��HE%`��Md�t�za��!��7�U^U��h�u�K�Ij��H(�����웃��S;(8�jp�d	ƪD�
vg�2���s�ջǞN$�l������;���r2bG�\g�!^8=��`{����"	��.����!;��Z��o��C��{_�+*��?�W�J#��Gm��֦�@#�?Ae��o�eC0�
�w��vE���J>�
��b�J�Y{`����u�t������[�cMR>��g��7( Q� �^�9 ����8(Ϸ���&��?(��3jDЕ����Ʊ�[�;p�*l��.g>��^r!��W�.Z��3�á#�@�%�T�>������9Q����X�q���V��]�� �h�p�8}�y�NlCϺ�W��;���;���1�=J		짟s���o�]U&�ֵ�RU�B(ZPcMy�Pp�NΑ���?D=��#]�G��[s�,^���uPo��b�qAzG6�mױ,���*3��:����$b��.j�3�ࡩ�q,���T����	����>��m݀CJ�06;R=�(��e��ۑ���s��h��t�P�8�K�d�PZ N��j�\	Ȩ�����ˋϹ%w�i� �)�6/K�v�V]L_*[�7q�#��_���)j،���=�Ĳ[J��u9�>���!�G����s%��@�K��\r!���Zo�]p�����D�^���\� ���e�2����bH3��+��)�z���S��I[�K�CιI�'i�?�*K`(4H��1a�O'���wʋ�1�S�Ά��4gV��3�8�d������U���\S��p�Y5o��qM�3I��'pZ�~o�ɚ���OU��1H(�tn+�C~���d,�m����2N����Qy?P}.��)WKC9W�xVƈj`W�:�(�j�s]u��������9�ք��z�o�-B\���%Z���Z��]D������  ���EV�#"�����*�i��7˃۷�|Z?ڗ!U�E�~�v�jg�)I�.�JJi�� Q]W�n���|�١�X�ܐ~�o3_6�lҿ��Z��=L;��arr1,����5Fӎ��k$�c���Ԭ�/�P���u����q���x9��\������Wa�m<����D�6OYBY��)�:|`-��`�C'�u�=���t($:H`����I��f���@ao���m����Q?G}��9���AOn¢Rr�>,cI�� �j	���;Sm �;
�vg�'���0���"&J��h�A)@t�'#�s"�+Ι<J�̠Rccy6g8�Z�25�WyB�6�0�-l�L��,F$.&�I���l�y��^�}>�����V���h���2�9 �8(�D`ֈ<a�Qi	a�BF\�F)�Lv:p%//�޷��۰�C�7.8d��mpg����t�E�E��6�@��SA�r4�]��d�
=��]��Ɖ^nA�[ٔ���W<�ښ\d��JR*�~O��S� JJ��YѻyA��9�n7Q�
c|�j�"�)`	��J�X.��ƾ�<Wgy+Æf���O��,�1g��}H<����Z?�*檵�F��
|��)o���!�b��p<u�k�}��_�p�4�#op�=����M���2�*7 ����!������7�vׂ�L��֡p����wD�7H�ԧU�L�m0��mf�7�I��:�q��류�J�@�YRc���<��ot�"#,��� ��{�0�or��GƫY�M1�.�f$�k�R:�b��N?�<���10�7��MuK���VRAC���I��z[�ܴ&��c`����0���?8��GD�aH��.��nU�l����9�p~���������ͩ��ǁp��<YS�N;e��(H�$o�hȟ���ݢ:�_���d�	d́�c����'�!U���^s}�qE����|�-{����d���\�`�5�"1��b�Hؒ�?y���V7���A5���Ob�Gt#�Vt%<k�j�L����Z{E�d�����}�f�u���oÙ�-�V�z�cG�Aw��2��[��4����!���<J��A�C�O��fFL��yE"ڕh/���#gV�r⦩�x�>U`�	��q坌A�O���o�L��<ߝُW,��{ul���oA'W���Ǒ��U=�D��Y�xj$S�dD����,\�5�6p�}�|�k�[Ө�f�T��p4�`B��B�j�f��BGh���Aެ��S���*`���X�;�\{�ϝ5�h���'1�A�T�M�@�X�����=άhc.��RΨ�b.Zzv�4��R��� �Y��A~?�Vz�oU�܃�H�����ezrMG#PAMO����>1�iVi`S�+�D�Ӎ[��K�ݞq^� �'�="&�$f�ވf0c��3>nf<�|����;��K��B��p�zL�ډ���;Y��eC(�N�'�K@����]�F�d{��m�- mΒ���*4:��-�ח�]V�'���{�O��´r���q6+�`0pʗ��� AG��G�	e��_e���OCPw	�./U1 �(�	�ޮy��Q��?U�x�Σ��]Yt�y�o�h��g<P��#�a��1�{Z ���9ѶAf�=��4�Ы�{��(��!�2�7c����`Y��)�"5��S->ou~�Ž̍ZY�W;\gxbﺚ����K�c�	Ka6�����Ǵ�`o�=���K����ΐ�>�qKC$g�̡�Pu9��*E-�Q-~<
Ң�MN \A�P��;��]_�r�� վ:�Ռ�:]G���=S��5��=zZ_Ƶ��w�^P���D��ll@1�9 )�kx�No䛦�!�Y�G�E3�&�fB�J}�l���4�S�$���=�e���6>�p�L]X(��P"�A���)]@���I��#�����T�B���+��41�ת���J1��#�Lq'�J�t����R �-�Fkn��5rW�Q�v�L�� ]��8�3Z�Î����ćǺ�^�ٳ�����w�sea�=�<V�n������';[|�V�` X���R/PLe�ʅ;rD׳��wK�1���R-H3�{�MzϦ�� �V=�d���k�s���/ܟ��C�t���~W�x���3�}�[,
��"���~9�f'3�c��~*����\�*��Avd�����:1r�=�G`��I��"^�fx����J.E�I�/��q+(!��+�0��,�%g�c�Pm�BJ�7���1� �~U��m:�ۏ��C��d:�-����W��y�U��#�h�U�QŌ2���zX�h��khŋ2�����`� ���˥�}���ۼ���M���%����0I��c�h��DW c�,p���ʲ0x�K{���nzR1vA�g��Z^����u"�`�s�bf��;�a`�s����7#��%���m�i�rA�sMyVނ�>Q�̀C�ŭ7f��'ع�yE�bw��b1��eI��mR���ɨ�7���5���(z��\޸�H�?X`Q��"�o����Cn���
$���W-D2�X7���GY�7�S�n�y/D{����r@*@��������,����.�����\�_��DA.
���8�-�EM"��}c�Z���X�	a�/�e�!�Q &�1�.
w-�Ay�z�,���-���1�M��ݹ_ެ؁ū�`�?)J��	�(��ӋC������?�l��'����¬(�Ty����D���Y�	^��彺�j�+�;�*eH��E�f \�[Un�����g���y_��ʖ�nl�.��6�;d_�Y�p1��kT���V2���k~�>E�T��4��î���?|}zw>�B9��#fUe V�B&�i��9��A��&��O�څ���nh����x�܍ռ�T���7�9nF�ׁ*i��sز&���7�e����q�ڻd��:qNkN~��-5�]E�;Q�B~�m��v�I������):1�wP�R�U���� ����^3'�z�t/�6\���A�ի��`������yfGf	ģAEwkPz:\8z:ӎ�~+�<�B��ʫ��|�ID����la
���b h��?.��F?O�N��u�11���4����]��@���r��Fn��3i!�W�o"�x���S�ڴ��G�g�W�ѕ�c㦷ꬪ�_�3�#������m&U3�p����C���s�
dU`�qb�ˣ	���7&G�4�i�\��^HS>j�"�e��U�' �\�޾%���6|k�U����Ç\��`�CuȜ�h�,H�C�!�������r$+_��(6�ZY���>�:8',���p���L�!�W���zc�$Шn���D���k�׊	�X��,�����.�YCha�cJb8t�	��%��>D���� Q�X:�
�.�ߔ��S����������c(� w��bA�;O��|6)�^�,�b�|��J�IF���q��(�D��rd��˽op7��1��k�	Q����y��%���U)^���7N�'��"�� ��M�ow=@P��M�&��J%�bY�(-��m9Y����SD����j���,J����v�1,�S�d4�Dq!�Q�U���Fg<��X��Q*-��J.�
�,J6v3�(��T���GPZ�A=�h�}�+�4S�`�P�����"�K,��G6�p��sމ�����A`��r��a%��0���0΃����նW�sXo�Iz�c��'�o�bD��}�ዼ����?�p��m��[�΅D��_��P�@��I��z��O�9��gh�}(k���P�jK���r�_��N�.���7:ۖR`M�w��h��s�|cUNK�:4/�G���/^��R�1�֧	�se�����7kf��0�]�C�Pvu�etQ�u�m
�6�ģs���{I������\ b{�G��L�Kš�J���䧆	�&Qo��1ӕ��jE�	�Qr�C&���p���8C�s�+畳!*QkW�O�8�$��x?B��um�ᬘSŻ !��	�P�o�g��u�sn����9����/��
�ޝq�����&��d�_��^���p� l�4l��8av�5����,��������5��cJ�XO?jEO���>�#&c|՚#	v����Q2��	�W"H;��]aE��Z	�P_�g*FKD���E����^ەz�@��[]�7��#���p�C$s/�#l���m��)>��On�(�tȡerGMqvF(�����Sb��O�̩M��mڙ� eB�CM�88��ix�?w����1�d���/㍞#��7���@����Z����׶��6�9�辀/���זPV̙xX�
�M���+{}��t�w��h���O2	\�������D�%^��+=� 9�I���D�׺ZބxFϼ����z���,X�ɓ��V��.D��Q.µ1F���6!�� g��R �z5Iz��W�6xR�M��Dz����f��*v�9��9����s1`Pf&�,���K��p������x�C~v$�3q5�6�d�W'5��˂�{̒�}z�o�_��?��}��~s��~�I˅eQ�(Yf�M�6/�r��
��{U�ML�ya:��#MQj��~l\E#-�i���k�$���M3�[?i��4���o��zf/�9��1@�	*C[��c#X�Ԃ"8F���֔2���p��P�11�D���nK�6k����3�	T���6�T���;��x��=
}U���b�*�ѳ���C	���l)�vC<���w�_A�,?����_�{�.Y�����}�|���h`�-oQG��!{|�J;�NM� .�g��'/>-:�!�[R���u�@��/7c*��~2�.��4}�<�������U�$�4��M�[���s��~-������q��>-�]�p�2	a���^B��Tc����c�(���D���C3k�ث�Ӫ�߹�t�ǝ�p��^�y������+g=�O�U��ONa�&qY���x�Q`�g�ھ1B�ݾ���x�N�9?@�eA��_�a���'�#���kZmޥW��܍�)�>P�W�1�����k���#vVø��]M�H`P����'D:�K�7�H��y�c)�E�]����	LbU��x�k�/zYU�[Z���p����(�q#��iq;�^o`�֭%�R8�BE�DuG��d�Q�=������J!vШVO�����=@����u�<`���[N�t	!b��X�i����h�)d�C��ǧ���^��G��^8)�w6�Bv0ɢE� �v��G��s��u��z�u�_�h�Z�cN��KJҸi�jǣ�`��!�����c0���֐��� S��2�;V�xD:��r=�&��ق���9(>��������k�r͏�_�9,&�'�Ս��p+Ų7�z��T��-O:�:B�2�ջ�)�iK5����I���7Q�{�OܡO#��2Ί�	1�Rw�8˚�]ΰ�C�A�˚|�v�|Z��8﷯�)ӁD��
SG~x�
���ՐD��|�mq&Ӕ|S�U�j�h��"�,��!
[�]��>z�Yd��b��j�Z;S��,��TG2�D7�lu;#�u�xvNK�����KY��d��A�B�Jj���8:W ���4>WD���Չ�����Á�n��6�7]���Y� �$��g��҅���M��C�ř�0UU(s3�cl1) �V	Fix�@�Y�o��Z薵�qՎ�.����˕��,ܸXs��ۡT��n�k�G�΀~Y<�'��R�F
1��]�R�~��)s)d��9���&��u��ԭ^�d�����^�`��:��6��X�e-v�@>�&��P]��֌sH�0���ds�G�xj�T��#�<\��>e7������4��v%���r�I^ ��x�]�׍=�ݙ�+3A�W�����s"�3C��H�z�Z��B:�F������{U*_ 9�/��*p��+Hf���04u�	��c�8]�%�&�Pv�a-�X��׸�v6/����@�pbyb9�bi�D�!�3��O���,�aY��ߓ���);�U��~��^�G��Z,�H���<�1v܁���	VZ�4�bόaBȿC��z
d;�~q�}2%��P���6X!������� s�{bv����J\4L�X�[�;�=��n�1YBW8-��H���:��p��_����T������P�1��5���;�f��;@?_�|����u�Jp�q^̭}�a����PNl�7������<Ǒ��\P��T��7�Qq5�P4��L$���^��:�b���c�R��1��L~f�;���e�i��@"���ww������Z>�4��h�����{
�`7vA����m��;�X=k��p��6����|rc�h�'���F��Zg��f��R�2�e<��#?b�AΛX��
�M�m��<+K��q����.���M㉧�/��m��L���va6�d&dj�-ڢoY;��iIE��(�Sy"��-�紿��vي;��.�KLF���:����;�Y}�ڼ��j;7� �b��e������{��r�+Fqlq��o��S��35(��^l 64��Y(���lR �P�L�6_��-��3��K��?�LYZ����μr]{.��S�F ���gH^֘�6gm3(I�c��RZxD�y�������`'Ii�e�6|r�_E%Ko�?����r�z�ĩ�b[��GU҃��Fӛ�E��,]aP�a���+ө{�����g�t�'S�k��U=���l�
�
��3�iUQ8�V���d��\��Şb9^Ϛ[��7.��� )R&������%]1�8�Β	M!��6򑗆t��%~��v�.��v�*��=>I�:�#ډ�b[�~)�Mcv���	A�໬ox�^$�|��l��(h���m��y���W��TL	�!̇���������CzS��(�ɫ���}r��]�F���.��|����z�h.�T�	�t��k�Vbܱ��ua[Dw��ELݽ�hT�u8�s�"�� ٪<�:Q��sh�@!*����ߩ e��<�?=���M���V+�'-tخL�z��x{?J�������OYyl�A��$��gd�ڙ3��[i���RKP��Q�h��a���lH&/U4vMfʲY�%ʦ^1�Y(�鋢����f�����l��l���5uL��v��k�hH�h�J��;P�n�a#��8�J7��폔���O<��덭��jp��l�{�s�߿Ӡ*|n7��m�5��W���E�A�h�����Y��F�7%9���\#���(t����I��a�%n#u<[x��ɷ�tW;䭛��8e���6cD��~�`;q���nN�o��
�'i�z�c����gхi��U�����M����	8N�����q�.{$:��|ݨrè��@�;<�!��v��:���~��h�ׄ������v�s�RN8���o/��ѐ�u�+��v���m�N�F�F�j}>���z�&�����D��[�e�"��5v����O'�����{�)'U�E�&Ά��dLq#�M��&�]�������_����ϴJ�	���/^!��{���{v6���C������Sn!��A'���1Q�1��S���}���O��Ӌ�T N���<��sqw`��g
�_G�����L&����Dä�Z4�n��0zZ�	��.�]�h���}49�X���l��a1gf|�f���{���Ly0���6���8��L�y�����*��5v��cΦ�S�X����N{U���<5���e�h��G����A�q���*[�i�9�+*A��҅ ���W�5�d���,�)p_ky,\&����K m���>=���g�G�%����{�
 ��)��	��q���rx`�h�C�=ؠ��2��y�3�4��Π)�ZmvтҼ[1�/V�^��Q�l
��eA;�C���:���j��>��(Z�M�'�7����}��L�
��A�U�%Ӌ~��(oS���'U��������U�D	���5�`�ݸ7l3�1���2ĉ�����#F�׈\���@#�� �ë+�]'��v�ܸ<��I-E��F����CS<����� �Q�$���W��C��(W�\�4���N�`R��i-"�O���0��H,�����g@&����jնR7U� �
RaE��W\�7��9��_� �)�{9�ܺ��E

�`	������M�)�ʭ*�����r���_�;3���  ՈPE�H���ȭ�?�u 0Dg�$���:�[�]�;��KĻt eTd����V��}�?�j�8
;'Vx�;U�1��}����$��@ȟ��]��D��X%����mf���(�x 폎��ʂ�5��,��OM�����S��J�ߓ��9�7����ԫ4A� /r��U>�^'z�<X��u��E��Jd����u�:��]ڴ�~��:�?���o㾡B�D�;�_���8�L�n ����J�[b����ޙ�P>��U�էo�GK@���y/���ƍ���,��*x��r�D��|a��I;���٘�C��;H�u"Q���*N�_��y~<���
l���	��툀�~�SA�\㛂���j�흩��&�����Lzr�'7eg��<�uTlp1�2&�䛳r��v�R��5+"����d�yn���|�!ӹ��s�Dd&ݨ�i�
C�XD=����}�:��L��$Q-���L�M��~x/���6E2n��0����OM ,7�h׍T��@j��6���
y�MN�G�8�B� �m'j���m� |��Ä�|�0gSRF�9@��GhZ��΂7f�cL�{W.~����}L{�cb����Z���N_��������,wQ��+t9w��E�?��|���[��Y�3�
Z�y���� j�V��������Q�y %j.�)X$%W6i]:��"=��H6�KtͷR�� <�����
` Da��6��J
��|��;�c�_�&H���KA92�F:.�����t�����5�s���E���O]��y�Y��z.�;��p9����=i�HT����� %���[���#�����vP�e�YwQ��*��#�՗ݮu~K��w�	�>��K�H�V0���_� z���A�T�)(V<e{bjmO>�����I�plNW���ѐJ8Ϧo��2N���K0r�����{X�r�T���g6��b3J�M�W3�ْW��l
:�p>��g)����Zک&�p�7�tV���i w�����LZ������,HDɐĻ�{H{�!�`<L���	�����@��F��=r����N�]�<��$������[�V�HY���*[�ʰ<6>Җ�n���؊�=�zb�}Qg'���?{����ځ��� �r8W �5=���Z���0�6=Pۜ�wֺ��G��qqg� �D�B��mO��ǚ�$�A9 k��7���3"�;S���#:!'����"�e=�+�^b��8o��q?2�?�\(��:=���p�4�]H�>��e�|�#�e-G:k,�w��W�*J��_	�,� j�v��ŗ%�:��Xp�3L���ޅ�.�M����Zȗ)+Q4~���t�]Z��`�wŵOPf*Ӳ�z㮔(���?'|�~�N�h�5c����Sk?�r^ �L�Kb�ij������*� ڨd�^�Px�?|��H����V�[�r�y^��R0&y�=e�:���Y.~k$��M��� �\����|&�= �-T/�=ؘ���opB���K���o0 �>��Z՗�'e���n���iy̮7�b��.^��'`��������,m,�\Ѝ;��U���@���MZE� �|�Z����Y���j�C2h�=iC!�Rxv�*S)��4|L.I��d��V�yfH]f]�l�\:�G���c�hsz�}��H,�@��F3@��%叔3���\0'+�Zcu�� �1�nF2� ��� qdEgm�g&tv�g-�5��q7-�T�:���-'S@�Q��8B�#uѸ[�kd��gPhpH�<���D2�ptY�TO��:�nc�o�Q�Ű��2+�|a	L|�R.�+���i�@����N.���W
y���|KB�.�-����п3�j�e��SB2ю��RA�s�MTd���wł�����7�3"�H(�F�f?5�!�xQS� yY�Ts=f�/I�S���֞�����y������,T�D8��I�t)Ӌ���E=���y��LV.K��N.�<����I/|\:��X�������"��>֦�Õk�wM��7P�pv bk�<z�bX�.j�G,�i+�/.�sT;m�]��ZqK!~#A��A� ��]���0@Y_ǡ�Z��گ6��п���*)� ,�@K�I��V V-X������M4�3�"!�^�#�:�ط6�$�:�i/oU�[&k��;P�K����������V�.֓��R�j�y�����QV@��A@ >���l0y���T�_ ���`�A���t·�$f(�1�f����:�d���@�!sb�<�
�BR����\���%޵, �YN��B���Ե/����/���������Mi�5�u�Yr�`���G��½�c�A�Ճ<󹠛 �.�1�q�>��ˣ�o�WЅ�(xA'��4i������/�����,L���3��F2q_�J��L���;�h5
X$�8fD$��	�te�S-��6! �@�(3O���-�AO"5��d)&{�S���'�)�CQ�yz�^+��f?^���#��a0{W��E�F�i!ּP&�*0��|�Q�"���5��fn�Z�$O�@�Hx�� o�1�5ۭo,�t��˔�)�+�=s$b��=Ua��O���2MU��4�����J�?�MՃ��}"u�^��
������Q���P�G,V��o���&L��zJD�}�����Xʚ�rT)5�5S�!%8�2`��D8��Oҥ���*�c:R��!�-x�!^�`$�@������0kˈ&rg���1�)�MA?`����m����!S�"���U�@=-����+�������=��?�V �O���V7�a~N~�����[����+}��E����"F�3��s/�٦a��k�3�6fP��ߵ��d��R޹0ȣ��=ު�;���D�����P������g6�8�d���R�_�·�%^�*�\<���;퀸q�PD���cq�G�]n��[p�O^�&i�WvHk�.x�[���|�jrw�[�����C�ks��"�̒��M�Q�EK�@eP������5���PNaGS��F���ʪ�-ANhޟZʨ�6�^n���pPb�l����[�Yo�,0��vULb��,��"XW�aĪ�^yV<=@jr��f����a�'�i�����% ���4d%E���ն�g�Lo�$������r=���� �Җ�	�����=|�崙C����"
xHw�R�R�07���`�p�ȗ�֍6ۣM^eʌM�K�9-�Aў�5�S0�gb9�^ɲj�q�Ro��z��6J�;%V�
5KZ��@�dR���cvB�j'XI�/һA�ZΙ��28p�,_����8�q��"��M_��2�x?���LM��{S���1��S�e�Y�r�sM����-&l�M�1���j� x�=��pt[@�=u��<~���=.�{���0���	����g	�c�����ķ��K1>��]+�P��	*y��F�4���"�"�����aش��h���L��M�A��G�U���+����w�R��Ap��u1�C�`A�t?�
�A+e���.K}���8-!Me� �k�آ�f��MBc���v3#�"������$㿬12�1h�n�dA1l�Wr&Rs�g!+�XM~�N���M�ݬ��4j��	z�mOQ�k�v�?O���P�9y���w�x8���_+z� '�r �:`J�w>O�~����P�Ѡd���"y�T��z��y��I�|��!]/��-�io p��	�v^��V�_S/j��W��0��Z���r#�(��wOH�6�홣�6&�!
;P���>��k�;���>�����Y�{t��=�ڒ���`����Dxx�cO8�@0o���or����f]\���H[YǜQ;��SR+ Z�X���4�=��9DY�,�Tt��.u�����l¼I���4):�G'�&Xr����DB=n}�9^��ҕ�t+B�n 
�Q����.%?�R�Η�QZ-+���5����cy��h�& �j)C\�e�@p��+�1s��".�0|d3s�hÑy��Xb6~�p(s񵦌w'���;�-:l��eM!@�s&Œ�7Ҙ�����(A;�z�v����rԸ��o��d�=6��3�l��Q�@����Z�����w�(9�Tk�W�@��Kebq��7temaD�^_��ގ&*�P$(�m��M���7��Yl�仪v�V���+�;]���օেK��:}�7���V�&k ��i驟6�@���EG����fڿ�p�i�>�J�y�f���<�E�U������P.�>�_)�]�W,�g��;*E�)��>-H�ҽXJ؄3B��ƎѢrjL��<ף�,��N~�9u��Xl8ʋ�9���
�2O���U��y�"͒��{��>�o͌��x([���T]eF���8���S+�OM��Ň�f�*�V��*_yl�f��;f�D\s.�݋�Yu����Y������!�G��
�[Vb�����HeJ��I,�~�o~5[�m�U��Ʃ%�
��kD�r}DS��ˑ@�6;O���};��d��j���؃�15I�����w!�x�˚x�k�͞X0��$��J�`��A7-�;���$=��Ij��9�u
ն�c� ����q��*&)s#�-�Z�����p�A. ^����i��/n4H��A ��X�'�@E��q�5��t"]T����xa�Ј�~x@'oK�z��D@�m`o�jG���{�+8��WOgP�0�&vb��9��Jy[cV��J���5o%^
�7z�u9�{F���s�Y�@���/�5t(�@/E.�w�ʜh��������X�ɲ�Â�9Y�![�P}QY���*�}y*x����cB:�ċ����hv�PV=�U&z�c-_��S�����G"3ް%��j��	�c!��9���(5�]���{�K�8�k'��"���-�+�J��b4�\/7GO,L�{lT���#jH ! ��FCŮu�o�{��L��չI��`�A�#�* �Bf�{���Hn����k��6�Tݗ%�e5q`ǭ�Է4Ko�RL���m���&q�I%�?��s�a��(�h����53)C�@��@�%[`�/�l�F��V��O�bI��W/��j���'{?� �޾ �1\�8$��[������pP����b����sE����g~�l�W�!�ʹ�Y�
��S<�x�ד�q.�[C<{��k���W�l�W��絙�@�^)R�݅0=�g���WJ9�5��������A���H�g�p�����Sv��#� ��]!�z�zDӃ���JX0qG���w�G�$������I�Q)�.'C4��jY?Q�eZ�������Ӄl�j�-�=�x~|����l�V�"^�I�mp��"��W��x
�͙�.r�Z9��4���?�"�9W�nQtR2,�O`���z��� $����OGh�]p�^�����`�J��
LYm��5FB��)
����^�6F�M�����\귽*75�����*,*��0��o$��^A����2aS�6^�P�z[�x<kÜ�A���67�����Yj��j���)R�H�S��懴/)/����yb
��\���)tx�h�C�_�0��*�J3���o�})���<��Q�Y��[H��'��w��_����	�:�v�q)̸��
�R�N^T�(���WUDiZ��֎7�9!`�7���<��W��2���7��>��1dw^d�7����:�U�3L�Jr�λ9�tz�����
Ee��UAD�[�T=�����鈐`/�=+c.%�hQ-O�|�J	u�vj�>Ǿ8��0Ab��U���V�F.l�'���� 1�◠�[D���VU�������1�,<`7����@V�5B�d��,}s�ͣ��x]�3~�z��gi�\�(��Se��	�+�6@st}%k'Β���QA-9}1�`;�ΜFm4u'�"�򊖄�0VE.�|����s}�g�DyP����P���y�\(@��C�&��E>˧-k��:S�Ϗ��5�2	�W5����G�)������8ـ6��r�t8x�cs��>J]FV	7�6���v%�@<;,�!>St�X���<slC�7Y�ֳIh�D�+��G�T�$�?�08�_D�%}P�w[#m֟V��OA�X��[�ﻒ)!�8e�
�pǌ��={��zi@�u�ܢ��h������FD!XtF	�l�_%��L2�8�`B�i?�����*�e����J��%D�6E�� ���
��*d��cR"��e�0J�Є1'�|�kB\K:{��lZލ�gjM԰�7
�m�!:��*�?=g?
5
p����G���w��JB�	S�z\9�2 ��7�ʁǝ��1��y ��:I��
�͹'���ս�� ��q[V5������C��D0ף����G��	�(�g=�(�|ӧD::[�f���� ��-��	zEj���㠭�Xm׺w�^F�[39ͧ�(O�K��4P��q- sDn�)j�!:�a֥�7�9������G��f��qvc�2�',$�(��P�G���^�4�#�N�J�����G<%�����T��c�dK���v�RPQ��+�>��m$���)��Q[[ҿs�����B�a�M���"��u�!���vqiެ��Uv�w�Ӈk�i�Zd /�����V�V>�0fw:��-�_T�ڱ�{�AJ+O������X�A,��HL� �L�π6-ˬs�X��?6��a�f�7����On���l^a��_�x�;V0��h�W�VRY�*筃㚮�o2�!�Hg��l��?O`�|���4A�]ʺ��<�����@�eH��-w�d��d/��8�䍶F#2m�,^�����`|S��X+P��o  �6���1ꩺe�ڮ�qF�<��Ć&��MI�N����jW��Zce�@Z�6.g��)@�����N̰��2}I{�i��#C�)�8U'Gs}�����q��9xv
�#5 u��S3�4��&yR�J��������C��p�Yס�c'hY��ܣ2Z�w�*U돷�'c�O���z%>l�;TW�?�N6�E����V��Rh��
�^�j�c��M��-x��"�+�]�o5Ej��(x�r�(��m�H��IYOe���i�K���u�����9ǝ�Aa<EE�q8%6x�gN;���5�
�
C���	�^�f$v��c]W���r��9��Qg����WQj�r�l��ԓ ������6_[�%E�?���r��y���4KI,�c�:j+0�n����~��4�s�7MTiGw�YՠT�ي�Z*M�~Й4<�$��h�a�#�Į��|T���������59�n�nC�~�G��[���Xw�4� ������m�Y��m�Ƥ��+h;�.t��?���н��Pu��~��&��nf3�F��XSG����*�r��r��b���C�|���'�넽&�Ԍ����4��0u�:0�)=��pJ�����X�1�\�`���)����*ݻ���\G�����>1@~F�3��8�٘t	�6�gc�1%� Kx��ח�%O���hI�=�fԹ{�n2 �l�<�
wΝᘙ�h�qYT	q��:c�'��E��|��Ŕ�h\u�Z���Xk�27ʬ�A�cj��fSf0�6���V�/��M�jp�}a�6�ZH۵@iCm��.��ո�,=��@w�83�Vhk���\�l[��$��"��	�B9��ҷ[X�L�l<���@���Q#�Uv:�?�У�v�3���x�z��;��^G��%����n�Ϻ�D_c�u�FW;���4س��2���g5�x�D�xWR%w�7H+I�0�/�x<y�M?@f���	�?���� ��� �)��`C/0��I��Y�3u�P�wJf�>�R�����C;W����iw�.�88\� {���a�Ϧ�=���R�@��x=�|V*F�PHY���|�� 0	X���z��VO�TF�a�D{�����������42R��\J��{��f��{Lr!�n&���I"R���8���"�����'S̮ZG����OG���4���hw7�q���-+~(P��Ok���BO�Y(?'�i-G
l��h��Pu��p��/��=+Q�Q�5�(<X��@ ���K7<t`���RΎ?���)�w#җ�uK�ǀ���[.���Sro�^P)
m�{?��?&J ��5�xP4[��:u�67>_���P©��g�B}v)����L¯6'�_�]��V���働�=m�J���,[�Q�cҒQ�"��*�Ԥ�F������;�tw����Ʈ�@��6��2�������L:�S�t�ޏ�O�)tK��~�����ٗ�s&
��?�9��.�����o�l����U?܉n��+��|;bNm���s�4 
KU��!V�nr����: 8��gr���K�~צ�9���-@Լޠ)U��WB|�]���KZ	��4$�C6�ڳ��,(��C�iҮ�n��_oG��H��YT7�v|{z��}�	��9��t\��tש�i�1iQ�G����O���3#�^Nv��nT��Z�$�Z�Qm�b��쾄��O��J��ʗhj�<H�W	-�۩�6�
������c��i���UU��{ew�X�D�+�>(@Fk%����_����8�l���@\�K�a� ?Z�����ہ7�z�0�e'�(�0fGGȮPu�ӟQ�8�j]#�]Q�0R0%r)�'(���#B��u�Ѹ�[1r0dC)R ,Wg�����%����w�w�L-J�-�)����6�����;�w��ɺiz��'Y~u�+����������I!��	U� �i�ڭ^�e�5��"��{܅����3����;�D�$��
ZT�|���RMV PnJ��4�mpS�h��|�M��C���V�`o�a)s�:�ޏ�K�M+��Q^T� ���r�V���S4�LR4m2F.=\�'�4:��J�(C�>��buS%�T.��+���t^*3�5��I�}�=3.�\��vȬ��0'?�i�t����(�L�z#��|�E���|f�qT����]�,2K"P�!�a`�u��馘���F���#��䐲�z��P�+ JU�ue%̃\ƨ�)2���{��h|�Ģ���T�4h�M�FL�i*����S��|$n�vB��֘Go�P���v9���蕚%a�?���1����*�\C�l��HK�Q�/���@�J�N��DÏ�F�ȓm�(�J-g-������T�m����9u�������^ �Sw�.�b �t��h�U��Z���)�P�z�l���PFwn��	ٮ떅�'��HY*sgt Q��繕=��BF�ߜZoq�nl�KR~O`M��1��r(�zۮcv�w��A-���ǊhJ���b���9��7|-T�s�w����#���=^LX�]R��	[KP�?s�� ����ܒ�Nپ)0��h>��5l&��XJU4� �y�Gm���D2p��dr^5������Tv�ִ�1��6<����
�����7(�	V�O�چ��2[ڂ�U�c%��g �I�I�M�λ��B�<�| �$+ْ054�{\�yȴ ا���xy��UB���O>f��$�_Rn��e�!�+����ά��^� ���]��CZ=/ѐ��*������<#���Q+���F��¢��9��4�#ߕ���\���D[i�(在��(��ڔ��9z��yd�0�� �5+��T��^���3�r騊<�x��4�>&��r\aN0s��IZ��V/g���vw�����y�����X.��v��D�B�0�T���#�E�`�	��a�^�۰����Ab�}�i�=t��ܑs��]+���ϰM�GW����� ��1ry�_:�S�hw���A+:�1ZE2�e-�T$b������g��Q��B"�ٻu$�8�=ڱ��s?������I`���Ue�	���Rc3h����_掞#7Ę�٣��l��,�im�(��ù��}�����=��ȶcD`��E0��@��-Q����6%ND7%i1�{�0o�H=.[%y�e;f��[
zT#ҧ�2ŵ��=��XPKL�j�]N�Z�N�#>�蠚Q�99�w*ح�����A�^�Q9�V���$Rb�����4�s�<\)N� N��k�m#���9��>mg��M��ah��;}U
I����}�h�G��)q����a���ϡ��J���.���e6h`�� ���L�A��E��+����/�	Y0p��;-'�c�`����g�eZ������zl�X��墘q�� ��t!9�W��Qv��?�e�|u�s�v;,��o�П�3zB��2K��{� ����A��$���*�<T��,�}9J�D�YZmgN���D�o�x�ګ��&�e&Y��{=jA�2�!��\�,�����ib�|S~	^vDb�*5Xѱ�7��n��N4�M]����W�(��2����#:M�>D��)�ʱ"��q{3SqWwb�	�/>��i��E~�5;�E&�������t8&��aQZ�ٝ9����
C"V���pw v����^�����
�;�dX4�)������6�h���i��ђL�y/� )����]�dD�ی�)��׏>�95P�!�UmK��k�P�W��t_�񯻯I�nc��_��!uH���ۖ��%�BI?��D�5��r�%4�gowu#��dz�fߩ�b�*�!����?D͵�E?ȉ)�.�êhE:�奻��ʍ't��T����?�S�c����8;ؽު4r�Tځb�RX���_��&��+���@8�}7��a���y�4+q,��o������ȯ/E��0�3��d��(���w�v�����+�sX�Q���r���0�d��hD�l<X�H�φ!��#�-��D�l)[E_O!E�_�t�!L�*0�J
�w�sO�H#�6��f�sK����
K���0�Eu��E�$��F���7(�$��t&�V�x��E�������؎��~F�\�!`;q��/�-�6��{��|��6�;l�a��i����oT��3%�~+V��+������/Z͔V"}��4����BNrKG�l_�^��gN(����S޺���s�9�2_��d��+Hf����m(��pj������D��������e��qGH�ӯ,����ά��Ƚ�y��;A/)C�R:0���{�-\��Y��z2䭽���z�o��>�ֳIKg�թ��<虀�B��:�!�?��)��-�o�r��wƂQS`�.�����U��НG��ò�JT<��)��#@�mn� Þ~:�r2������p����P�v�^�4p,QЯ�8_��g���F.|��B^��s�B�ҎBLr7#��灚�N����^����{Y����\ZgDӶ�O�F7��F��3��++���0����W/1E�SI��������w�f��q9*��	Nו})ȩ/�N��~=�
)���h�?�d̍�ULu���`���Hh8MN9߳�&&��Y�"������p����,��MT�@@�ґ4��.-nb�@Q���{��U��J�d����ÔZ�~N��Z��%!�5� �k�H�����d�-��2^4@)�쏆]����y:AS�����̓Z�'�K�ӂ���M`���B�(ΪY9�?��W:촭>�
3i�}9n�MJbܭe���n�7~�ț{���ۥ^�Î��f��K�#�EA5�<�fr(������Z��YZ���d�1��~�;��q&�$!���J��6��� ��7�Xf/�^#��UL�

i39��嶺��T?�,�KA�ƾyFl��0���M��O�`�ʴ,	M�[�K�\9��?��7C���wUGEn�'�uck�)Ȳ@��țz�*ܸ�I��0�+�w�-&F�����P͘��)n��������5h�����j�:�#�`?eܡ�JI�w������_!Y��U���`m�����%]�kCwS%��e��|M-���#�S�ʧ��}�����o�.}5��4�yY����boԫ�	?B>�:��L��a*Ǥ �5�.�С�4s�ͼ�M�pu�(����{�{��%�P���-�0�����-珄�٭�q�����Q�5���ҝ-[H�y��ӷ���2'��qC$d\�u��P��i�\{8�wd#�<e%K�q�UAw�$��W�:�̨$�kE*)�䷏�졹�svy�QF��n��.�(��m���7�	2V��,�.��$0[��Et��ņ�^9�)F)��h��!v"�˄xJ�a`��1d��^�H&������{0���)�4��;YS��	������2Z�@��9�9ez��_�TH��I7z�#(�]��V��\�U�. �te�X��v�Q�����AXr�!�?�YrqR�B� �"��?K$S'��T��⺺F�,�L�����W��U�:�������*pd�5;�5����������|���v��o,D�������V�<�0�{YL���j2��1Y����<܆،)?�޼_v�YD�C�3g6���������,Bޅ��j�[h@P������Q�p�	�黪�1��'����tQ! ~��u������K�=�<O�Q���[~v��j�6j��j0f�H�@�!�T�_v�ܦD�6�b���{��\ͫ���J#S�@�c��K	M�+ B���G��R{���&�n�%8L�Q�2�m�J$��h�mXNH��>x�+j�����l_d�f�ٝ�.�l���5�DM��]Α����g1X���A�e��$�+��M����L���_�<�>�;GE0'���|<K�����'6/�Z&���ȿ����h���8($d]v�AoЂT�H�;V�Rh�(�i��(�q�F�V��7J¡Җ{�ż����p�@���,��Ғq�.[-2lqH����Oq�'��Ф=�������]c�ȵ-Т�M_�n��z}�pШ�y�����6�h���x�8<�ՑD�7Ȭ�@'�+S�,�f��)Է�1���BaA����l��)��@r�ָL���C���έ�Y��{����+��(9ե�����·��˹kISm]s�Z��9njxmp���&f�l<u��E��������c1�Ii���wҹ$�2��吔�*P�Xz�[]� ���/�^���2#�cJI�} M�gi�ho�N�8�(�Ȗ �i� �y���@�O�,��\��f��<h���],p�����S{�P�'�j�8�h��Z��u~$!���
汯������MC�K��8@�LO�udB�"\�)l �@���Ő)Ϲ4*��U��(5���l��l�sV^jt;ޏq������)��!�a��8�(9�v7�\�v��=�a�l���FAR��Տphh�z&��+R.
ê�2���~�y��v����Ȝ'�vF��U�qI@��Woח���������&m����&}@/�Q�
�L�Z ��;�p��E�5��v2E���9P�þQ����f���o��b�{61��=���6���>zr佬rPj*��q��\k?s$�G�3+%?��(JC���!7�DA3�oP$�_� $�h��g>�P���Ԛ�۽�Vh��;����գK|,8h�H�Щ�T0�Sy�ً֍1���)H���
.�W��g���G�*D�c	Ua8���I�mޜj���d��pv�o6[]`�}�,�Z?�����C��OJ�R�?Bs����� �K�"�+���!�L�� 9�UL�0�7�q��4a��d3w��K8<�NUꘄ�@Ж���T�`q����"�㭲�����w�]C
`�:�Ʒt��:?-Fif�:ܖ9�4-=�a[)��a��hA�Ǒs딪j��	-�a������X�����'4�����H1A�%����Q������W8V���M9��̩o(��q�p{o;W��!ob����ʞ�
uɖ&��ٿ'I�.,���0�GԠ���.���h?�1������,��K�x���hD�Xj���+\|��>Q�GA���]N���V���������2��a�S�F'0�}0J�R������	�9�1���YR��r�X`; �v+���w�:�`�Y�l����n����ziL�,��~�gQ�6)��9����R������?�h�P�8\����|�,䀘{�|�/�0~]�7v˕DR9"L���ڸ���_Y�b�pΐ\S��8L�R���^6y����h��I������H2G�8��:q^�ܯ�D����20��@YF��.Ʀ�j�f���������\�Ӛ9��@c�V�Va��a���؟�G�{�	al#��]��.?0|`�Q�]&�5:�l����WH���5D���L��f$�C�}����s�R$�9��H�+�����Ue�}�G�I��yH��$AJ���7{qTi�26�J�#y�G襭�e���n�]2h[��^�2i,�@ʰ@��,р'RY`5�=7!�Rr�z�|�-�R��+)�MRn�)��7T@�� �>�C����@���ЬS��"�{��Ki��.�M^���Cy��rzd0P���>jZb&�l|ԟ�p�M����r4�W.g���[����i���k.p▣Xh�n�x�8FV!�(��܋B�4+�9B��1,g5	�����+QF���\Y�:4� �\($�NI�L&Ԣ$a~�ƝzV�r|�`#y�yC�>�p�O�9���\;�:ۂΰq��>Ê�ǜcG��!�=��g��2���ǧ	I�&���G�*�?��#q$:/K�t��>[;����S��'���ɷ@��j����� ���OH���c!��Af��/�� f���KV=c�\�E6[8⩢H�ݎ�)~�^��d�GUp�xm��U�謁n+��ՍK̇]��q�RKͯ%�F�'�w���3o�n�9� Ob���i����E�D�2����ʤ�x����Z~�P�L[)*���v�F-N�LY cm�@Ù��I�i�r�H>���j⿾���cbJ���W�+���깅_`/N*E� ������WR����e�=<�ل���Ť���i�ƺ�H� C��Ǜl�����������6��x�e��\\����$�4y�o����`ʿ�֖A��Dk!�����E�N�S �:��x�r3"���}͂qۂ��8��Ϗ�C�#�>��X�j]T��\!��3��-��B��1VqB�:���h�H��Z}����׶`ang��ұl>���|~ɪ��|����]�ְ>��i݆'��6�٪�weŭq���H��ck$�T`3s \
����Q��y�%��nw���$�\~war�� �6ALw1��1�w�Κ�+O��b�)�:�K�fO�:�沒���w�=-y��fϽ/7c�|�l����-�}R�t;>��iٱ76��K�@P���=>yK���U�	�&lJ�P���N�I�������V��U)BQ,K�1�S4��TE�N���cY*�(��u�
�)�?j|��Y�M��]%�Pu���)�z�Ɓ��ޔ���X�>G� �(���@��E�E|r���)HbνmJl/
ڃ�g?2��/�`�_5OfR��fǓn���v��	H�*� �j��痧�J���p_:h-p��'����ó	�07�"3G�A��~��9��i����r�y����&�����c\0A��wh}ٚF�Ѳ��qY��~�uPo�m[�%�H����A��G\��bsJG|)�6Qb����͗T���t�Ub�l>�:}w�gl9I�U-.�|\�y���Q�Z��i�/��/B�P}�76|��P����Fm�,�T�
S����~~����<�-�E��ȫwJ��Y�� s���䘧�Z����[�텚0(�$�X�������ddΛ/����y 7P��X�oaω��A��e�d�пYU�P��A2� �RM��<�|����c���;p��x�H_�����'h�<�W�bc�X�a��:�(����OP��I��H�:p�(w���[��0�C���C*��5�����Ȕǯ��X�U���O���o{�Q{�Em�L�R�=��� ��2~�n!���>�
��ڊɁ��X��	xJخ�^ �m<�I�|�9���k�1�亿ޣ���;w�c���iV��k�M`t���aB���b�.~-!0g�v6`�?U�Z��/b�CUks�o	PM����W���U8�u� (c�rQ?&�m]�8�$βn7��F�/I���r�>������(T>Л��k���i-@P�Q�ab�j��)�'�lG�:]^+-��݄N�|%�l�je�K��7�|�J�3���U�A���¶o��i�oB� ����{�I~A�����E!��%�y,V��OIyo����$d���[��X��yd�@���U�?s��x��ü��u~������g wM�X����W&?o�4�]%����3���pg4J�e�����RU\�48�䉷���`q	�^�e(����*d�U�cA��bSK[g�x���H�^�#*
���[S�]m��N����K�g~��/1��&�A��$Cre��tS
�~��0f7
VEJ�6�h��'��*U�3�\y�gjѮ���*զ�r��3�D�S w�����4 Y��K9fL�D�a+�f�͟�7�,� ��vK%ȑ����������-�w���h S�"��}��T��{u�u���$�����)������~�2�1�ZTp�^?L�>1���*2CA�-��d��5x"�(�p҃
�k�0ʶ��C��ʀ1[�D���y��EH#g�Ӯt��2�g^�%�s>C�9 �J��R�س���է>v����-3�o6Àu�*���X�v�s�F�F�->��3��;J�2���)��d�Y͂�$�"��K���F��L|��_e��3�χ���z)�
���r���:��z��b@lYy)C���8�MQ����#�t�X��
ɞd ��˕=.�_%#�����O,�A,@����қVJ�	ܿ���av}�^ai��u��B����� h���[5��5��yn*����4��~=Sݠ�Q��[Ϙ�\v��>�V8����޻o��uꞠ�.X.�i��a��{�yf�W�#f�tw��@�aDc�l�g�x�?���%-�+�w��=O>����-�!-�WS)�:��!	G�b��.�w��������ױ���m2b=J>�q|0���ߕ}G�6�\����Y��s�<f�A����ؚ{v���*��Ӣ5yG�2v�t]l�?z�H��83�n���������?�F4ʙ�P��.���
M�E���Y�oզ� ��*�K�!�*f�3�5{�)������L�5:�V�c��h��m.�3}7��_X� �B�\��_^�n�����X�%�tkY6�ˢ��x���N��'�1�9�Ϻܑ���"0z��v�����>cPRځ[���2�Ԥ���o㗖����ՠ�����V,D�#,	�潛�gV^A�h�g�� =�������a�\��,�Iz�w�ٛ����Bj��"?Kp��0���>�v���O��)U�Uf�%"-�qP��ơI"�I\�4�"j���D�f�&�ͨo�k�!r� �|��셢���[^L�����´���Ν�q��b�L�Te������7QFpӚ�	k�u�rs���Q�l��]~���K���Ң�<�*�L;H�4JCf1���C�� 2�K1�'����U���|-� ��' ��'��b�	(d--AX�C�i�(�|򁫏[%�B�,`�m��Y֎��AF��A�&�H�� ��Zw������(5��=`�m� ;��%f� �V/y%��N�P�H�|�~��YXwn��ʉ���q��}Z�$i��_��J��ڰ6��c��w	�����e�����ҁ-h�Xa�#�w
#<��n��m"7��搶�B���L}ļ��2ӿ�e�c����n�`.\�`<�D5�K�6@q�J	�[�P���A�Wˠ2�N�����J�DL�+O���Q?Y�9*����~�}5ٸ�z���/���>�v�{;^����Jދ�-#*��B�,�41+�k�JȘ/���Hb��iTP��|�9BV���sMu~Y:/��P��CQx �%@�����:wS��*���2�=�7�Ye�m�ϳ�5i�#ت\4硫�8���u��[�I�����W���w	ߴ-ݯ��:�+f�2��ot#N�6SEӇ�z"��*���p[)��]1����� sߗ�>�<sC$/�}�kdu	h���{�V,���6@$�����Υ��$��_�/?ǸH�6����x����á@���AS�Y4]�;����6���ܜ#��Ņh�q�e����Iﮂ��\(ۧ7Ȳ_'��~3�U���U���x��	�^C�،�K���n��֏��^����˒rjY��7�7�y��&4?�ɕ�Ň�݆g_�g����#�3��iO!��?c�b���W�H.<���u�ߕ��c�6�\"�Pœ>!bJ	�y�|�����r�V,Y	�32�iъ+��/횴�ӱkE�o���#�\����1�̖�~�]����6��Xv��~�ٞJ��]|�	nvD�Z=W&$�n��\\mf��6I��y�m��X%�/#�V.��	&�ه2��J���w�a4��1���+�~k��žyG��۫��[K���u0g{2)��V���q�����df�!��}eސ'_VpX�̘��f� �D��o\ǝ��nv�(�FT�*��'�JCf�dO���������gG~]֦� <D�(��r����b4��+hg��E�K�������]kNDm��ɳ8؆�����M�li��g�>̤�%��G���#d&]�43�X���@��m�����h��&�~�c��/�m�&�X"��Xfn
�A��w⁐w6�֨up4:m6Ruv}���5]J�kX���N2����$(g���%6��tc�D��cɹ���~�J�RE��н���I�z@[�T�٦��wh�J�8EO�"�=�{�ޞ�Г���`�yH�.̇N���E��i3Xj��,�w��
���ԡ`�
<�&=�ް�ц:��w�����S���*�&�Ҹ�P8�d���� %͓�,D�$\��d�6	rE�#O
�\�����GnL�`d?0��;b���SR�6�7Lg��g���wb!㬯���T[Y�{�M�Y�,��C�Ru�F��V���N��ȞG
�.=�: ��un̄狙����S�إ���lT(>�^�{�z[1O���ݷ���Y���o��A,*�H�ê+�4��V颿��ky���dx�e��k��a��P;�A6�-#�~��#UǬ�<0N�'4�Nɷ,Y?�O^��|�3x-��]A��BRg3[�=L-�wqՄ�A��[4iR��/�F��D�|d2��ѡ$P����+�K!�Sí^�e6�8��b��? ��T�$����$�X1�p��,����~�� t�8�Y�l�JZ�N��yh���G1�+CR�=4����X�����#�l`h�x��^��E�� �|Ѡω»u,�K����A��M�L��1:��E䉔tJ������JZU��]ޠ�����47Ȩo�ˆ��F��o���p��r�}�Lc{1��Jlڇ�
]p�܏rG��)�|�L���΀� %������\�����1ƾ:�lYI~��J��%䟛��c�0N����׈�\�]UVQ!<�����E�G�o��U����M��k���$�]e ��~oiz��$v�D"MX�}t�E���{�aA�[�M�pi��Q	J�	4��?���'��Yo�фݠV�込j'DTa��b��w�]1��U#�TkK��G�ݍiFϵ�Ǯ\�g,���FAȺj����i��/?Ñ88��B%S
)ȫ}��$&9�1W-��s(�>H���Pй+�����y���rY��V5�M�����~|�I�5��)DU�%ޕ�U�M�J�I;0!�0.*2�ىp�C�J=3�y�'��^�_�#Z��܀(
��e���:��,TL�a�����s@�1��7R���S�Z����	���	���}��_%�f�(S�����؛�r^�ۤ���cz����8J�Y{�;e�Qd��M!��Z��H��$�7�А�~�M����(��а�>M���O�徲]TpF��p)�O� �@�`��ꡡ�iVʂP{<���:�/�� B�ϬʑZ���R≯Kҋ&�dœ���G��";��?U��}�l�c	����Qa��>��e�Y�}`"%��<v�k|�#����E�+;�vb��b���H��!C�e&JzK5ԏ�� �oT`(hs1����we@�c,L��DT_����~�c������(���m�)�f�۠f��U�ҙ����*,��:|�N��A��`�UEV��u̱�'k6fb��ܡ!6��d����V]���|����X��d"�~>E3��@�qE����H�`�?P;:^���?8�*�"|�c4!�	��t<�����1i;ݦ�TlMw2v���
6��Zs�h`�Tx/��L�%��|~>�],��PP9#�K�߸ds��I� �W�%��"&�J�UIDQ&����!E�w\�\�d��Ɣ%���E*N�\��4�	��Z9����Q6�$�7��2+�f�x�a�,�[V���U����1�]"�s�Уt������@H���s�%Te�%�^))�H�?Z�/������N��Z����Yh_!�,m����T*7�����>a�
������6o���.{'0�<�;�wN����a�BXkmJ�vF�٥*l^�Tm���\z�v���/�U>��Q�f����1�7�K��P|���(�Ŋ����m@w�N�9��f���P
�M�;r�c��j=aRY�^�U0��Zp��f�/��ȄR�|��lUq�ԯ.�|�K�&,(��C�A��K���&BE�-:��ro��$����K�E�B��:q+((�|�vN����2��~7�$�`��t+$�����Sڷ��_�2����i��a�/jKq3t&N�����������i���}1��E�:�@�{��@��(��?'���Re�wCZ�
@a]�Ə��C�86!O����O�I'_��>��*��Mb@	�4ę,�o�)�a�y4q�5�L��y�b�r�W��ݻ�s�
rƕ�Y���*�����{�2D-����f3ӵp�l�����@��K -5S� r�{�l��Pa��,�_���-#˲��އ��)�2�v١�<]s�<G�=<hFc��ETg3�~�	�MB>XPgB���uS+:�k�g�gJ�]��{:r��}`a<��1b�aK���!<_��e�K������I� ���e���~�;.�o:rby�*�nŋ��q��'�!�����ɩG]����
�C?i�n�W���H�^F{S;!;طb��+Q_*+}lu��VХ\r�Q @P� ��u F-�h��)1��C�OP�w��'��ђ��H>�|T"��>fr��!Űt\�)��zbj)�9�iQURd�#�e���ưvr�Ltr��
���#Nb
�E�R��֫��F�<]Q*Z�(^1�PQ�P�KR���̇���j�^�.
BX�'�h��[��6������Ԝ��B`�]���!]~ڪsO�'��S��@M��|������&	&k�yb-�`�V���/Xp�B��m���+����jQLa?A��O~j�Nf�Ob�Vz�K"(�,��$����(���p�uv�"A[?߃��z퓴Ue���[�9�Plav�ՠ
�p{#d����X{�f].��*P�K"7>ϮE��臘l��4����
�l�t������e��AGVt���k��X~7�Q���S���h� '��؜�q�����gV+6!��,��0w��l:%�q��+"��P�'2��dkVy��/cv��4�!������&�c��>����Z�;�du����_S�
�G9�.>l����yǗ˭W�;��춽��n.�(����7�Smĵ���X��N�0�T�MnWA�d+#]���6,H�k�9�����rÙU�Ӹ����O��rs�cۀ^�ډ&D�@zSF��r}>���1���=)�/%#�ڭ��ki��޸�
�
�����f�U�;A��h�U8m��o��6�)�SAO�c>I���T��%5/��z��R�F-�[�N�]g�Qf���.[M��6�I&�7�'�,ȧx�T��ܳ �s��pX&!��e�4\�-�΅]��[~��'ͱĨ�3X���v�]7z9�4��U�u�ҜO9�;G�i�!����ٿ���X��V}�Pk�\.i�K%U�r�8��Z%�(���#/�gu�|j�O��U�@��db�EW���Z�ˀM���g������0��*�u�����{�Sfr4�z��l9��RQ6/P"w[���hq�Φ�$\��^�A�������k�����uڏ� Vk�q���M�LjWH�ߝS�?Bz:B���� 1sy��S��>_!\\���i�����i+��ȥ���-w��(�{���� z\���������Ng��V��S4�1�;"��Q��j����Vܹ�b+NH��^�!�:X��` �͖�
�p��q�{��L ��~��Q�!P{)�?�����IH�֪������ζ�ېd|���V�vx�v>�գd�*RA���q,�d΄����1"nk�� �<�Y� ���݇����x�8��Sy��
B��$�+���L��@���fxl��?6	�6i���'T���$�<��yq�=�����z��?�8%�W*��iT=�G��J'%���:H7���"@�
��'�P�hl�x+�̀��T�O&����YW�Tm�H�9;���ogvMF�ŋa<�Xaa&���%��="��o��4G?��Ԕo���n���뙣��Qu�s����դ����l��)����"̨vAF?���>��k��GZ�-7��S�1�J�k5Cb�}����s�;M���T���lV%=;����b'��f�^�+��V�ʭ"��焏�P���k$�Q�i�+-���H���!l�J$�O���FY�&�f}��몾u�-�X�:M�3�4���ͽ^�Kj��������֯����h�i�8geٴRJ�I5�dG��5r�7����M�����L�����v�N���aXyp�����[�	�g�z֟�o�;YFZ"򟰖?�4uW;3�M��G�@�������A����v�2�iZ:s�c��7������^ m��^>F� �;���`�u�a1;W旵�i]�(�i��=kh���K��5Oe��rb�=�kʖ��m����3�Ӫ����Խ��#X�.$�Ȣ�l{By����w�4-ec
^-�)����D��$������2DN���P`�ץ�:(Փ�X���P�4{+��8���r@#@ez�Xc��3w�iM��g����~��#d�l���+���&�E�`|�yEe0ޚ�(nC�PJ����b��Zsk��ς���,ӭډx����;y��h^Z>\��������
Si.�А���G-�Kc���-��!V�ӏEs�qX���C
�-fr�O\���3`ol��'��^��=�:�	���� ��}F���7?�� �]���z`)0	fD�Y��T�1�Bh��R�vAH�7*��S��	�ܪ��J�	N2�M�2q�����������w�����I�Y���:)g��-��@��Y�'dr�":q/��U�Υ��Ȣ�/�=t����������*l?c��G��^cա��D�.n�#
ih���f���"r�c�7���Bb�;���g^�w�s<�"K2Q2F�k�~7��V��]�����0���oTT�[��j�6V��}L�?��9���B��'5�y�Ȃm%��<醞�����'�҃� x%�7���'9}D�Y���(O�B(�^�H�rE�X����3fު�n��n=�R�y�@�4d�Y�+/���1��=�������Ks9��]!_t�2��`�+�=(����W��S�)���8{��׆� j�@��-6�{v�����I���K'J�?�6�u��q(�6^B�����ν�<��4��u)��=��8�-T9�r�s��XɎ�du��$P67��� �3���k��b�9��eQ�-w��@�$`4!�BJB40F�7���+��%F�e�AՑ���������a�OA�ׄ$寨%f��C���-̆�M1�:�p޸��'�F��j���߳�x��甖��  s��H^(jD�p��@x��< T�>?��%��Fj����Y�V᦭�<1�c������g(���1`s����SCHq��_.B[�S�!
���?�A�ͬM���Ў�q8���=�&�ݓ��׌а4�1���Qpb���uG*`kÛ	�1�9��]iKln�U׊1�������M���0]6�BTxJ�sp*�'��N�k�#�'|���� X5��W�J���9�� �E,�"G�~#�0��J�47�3�.���af-e�&�
DM�g�Rr�^=+�ҒmD<z�F���EnNJ��I���.l��1]�o7jF(�M�~��t����p�}O��,��\�Dс�t��2��+�v������V���78TK��~�>�1wC�gi�u��j:j<Z7?=���VJ0I_�u.�9X��:��sB�)���"���O���%c�aW�� �떞Oܞ�ِ����S��d(��D"���K�_F�;��8%�O���P�Cd�
#^)�2�P��k�u� ������|��&.U�z{<sC�J�
T@d�F�B�V����} v-�$W�v}�󆃲�'@,�t���˽�Ԝ��ss��p�J�ѳ\�!�G�b�; �(W�96�7�AEp�����P���pD�Lt��R�~R�;�I(Đ�ft� ѿۍ��	jȒ�N�0G}�d�Nπ�-\}�ʫ�m�Q��J9ʰp���߻���.>�D�?r��`#�HuP���s}���bK����H�U��+��8��`�h�Q�^��ouv�O�-��	B������)*h��9|�t�I8�"�T(l�3��.j5ڿ}(�Z7�WI�3ŢlpO�1`*��S���}]��G3�`�����K��������sz|ݱ������.�.��ǧ&4�ӥ4��4z+�{~-�\C���o=��ǭخ]���%@��I3�bÝ	&jR�1w��9@	����3&�VeQ&Z.��2��Q�k�{ 7�����Ȱ˘r���RU�O�:�H!��.�r����'�T�߇��b��H��zȨ�\l��7�X y�v/eg�Ot�M���6�}~�UM�`�Fv�1[��=D0������{�Ba@�kW`��*,��4'c߃U�5���!n��m��`l�C�w[�u�=��PB��a��-�y����,�8��������a֪r��� �b\��m�
?�:M�)	��F���i�s91Q����hJ=�M��g8O�{���:_��[�Rb�~m���E�����x|����7*3�p,=Ѡ 89�.��l�Z}P.V�ЪVT������"��m��D�[�Ah	�Z�{"�����R�Ŏ�	���&t7�܊��s+Z�<����~Ym�E�oK��H�ªi��>!��=�v$,�R�t@�\�{.�pX��P;�$��r��,���Ja6˭�O� J<θ��E�2������B��W�Z��J+�̗P�mU��} ��'V��T�8����I?�r��eE��h�J[��N�B,�\�[�O)y�mM���I�6B6W?<(�)���P_���d^jb��܊�-s>"$5VSdP��ݺ/G}����6B�X!@9h�,J�POubP]��R�p\�9~f�3@$F���=�(��sQ)�ѥ�[���3����.;�j�gL�t��c10�����wVY$А�����*�ْ_�J��H��-���;��v�8}�W	�3_@����L8����n��,���t�J754�9CZ|T�*�G���\�v�+W���)�_�pD��@�d�:O?Z��_VVz����j�\v�&�M����A�E|4��%���] T��D*��E��y�8Z"��ߌ�����qm!t����$t<�L����$��������_=��Y��[6���a]��	�S��!F�C(�����QYG���)�⬦�U����2=�H9A^vJ�p��r&�##�vt���F��0�(5�DHq?��.�VoN��m����ʄ;����r���[�����z��|��\;�o���0��)�p�4},�Q^[׉�ݦ��/����tm! �D+�gjY�%��MN��D���{���I�@(UM��q8�G���P���;:�]�����1����Ѫ��֖|�Wu7����{���
���g 3��>�!�����L.����H��@t��l~������ᯝ"�:`G�V9���1�Y����n�%�m1h��z��\�� ���d*���ʇbV���ˏn��,�h���C�{ �J&��Ds�62P��gf�_.���muH@P��_Yϖ�$ı���#���bU'��k�2_��\�I�>zQ�2xY-��#;I�QHP(�9V����A�����W{�A���'m��j�ɬ��Y
���Z��vj����-� wո���s��ݨ���oô�/b���Tj�P��=3�B�W��p�������-�?W�§0���M�s��IǦL�u�ߎ{��v3F{��S�����꛰��y^��ݔ�������*4k�u�?�]཯Tv4Qg+'��̰�K�S���"Y�/.g@�<rI�8_s����8fG�_l��:��D�t��ݑO݀��S�������	
����ZJ�}�t�۝ɤ��"&��8b3���9{7,Sϡ��~g�wUo�}�&�L�:�ƕ���������Wt	L�G��J��k� o����A� ���³��VR�s[#)��`{9�P�h����ёXdϹ|��'���ʉ��laީg�|�hCw���Ն�N5P�p=���M�?Xɻ�d� $^Dd��dv�_��{1.�8h�eM]a��$;�� �P��AyFփϿ": =iMC�#z��`������L���B��4�;�N�am��2�����{Z�椸>�ޏ�za�XZ.�_��������9���>��柾��]I��A��zgQ�l9UgMclK�\��Ɵ9�k��A��K�}�;|���"�>4t�`3�! l��m���x#դn�a�K�ԥ_��$�|1��l��bHZĈ���-�p1�$FNQ��
pLg {��}�n4/�J���Q�M	�cD�d��J�i�fm`�*�B뇹��!�WE !,z�C�{ٯ�����\�	�7��kzm5���!9����+��%-�S7�c\����)����C��5qT�L�ۤ+j�\��q�,�4ڳ��f���lK��B���9��h�����׉b$��L�
���C��|p�.������[\װ`�S�����E�ڎ�+�{�~��Q��&�^f�$�� �[b"��I�(�G����hFN�;�pW?T)��A���	x��7� ��a���s���  ?�9�n��Z�� ��ߛ���&���93
4�l�s�/:�'Tv΅t��fy�&6q�+�`c��Π[���_h�_Ka�A��~�Q���[���w�+
_��4���d�s�I��kF���oXZ��K�����r�"@{r�����sX򓅗ճ��!Wc*40�"�U�uR����Ӹ��0�T����K�O=0�8�^'(0�}0���a3�8b�3Z�z��؛b����8�L��~��i������:en�q]�����|�a�k������S.�T���A��~1?��!��+����:Yc7^*������f���bcx� �E�ϟ��-+IZPS0���D���5<���k?�Jiﺹ]�Fm����X�?ܿ�b��8>���R��l�dC�� ��K�
����m!t�6�K-���)��d�W���������o\�>��l��U]�U��c8����e�d�����n+
ctL��[�{�f�����U!՛���~�Gˎ���B�Ym�%����ux�$�(s7��x�Qn��}�jw)R̄`GΣ��0m��|G��!�"r����%D�X)��r��*��9������#9^5���vڥ!|?�n�;k�f@�Q&�Yd��øc����ސ�C�w�h �_�0�}��A�X�wqUj�,l��b_W+k��F'�b���)��8|r���̂3�1���`.���n4�-�4�����j~�\�}In��o��-����e��u����;�H�������c��A��J��TTx��|�B߽w�E���R�����9�^s�m�/'�y��HH1��u�b�-氟���
���FA��?5`��g����{I
����2�AsتHI/�T���I��� @��C��=��!�i�>�$�a΋A��4Nm��e宀f~ I
�Y�9�zÁz(��&A�UQ��I#E_��X������� X�pn�K�����b�W�l��?�r�z�/�� /�QῘT`_�|?�q3S�_z�(�����2�����O>��J�J\�d/Ï#/�m�̜;��.���2�_�#�؀)�Bs�:�U��`�e��G��IL�I��
�9��9(m�*_�s
�4�yd��d�9�R�jNȞ��ރS��f	MrqP6'�9Ů��F�6u�m��:��ޝ;v�>��y���J_C�r7<F̢]�t6�2yp_zо!B�a�JV���<�k,۔A,���i���8q%�t	BՈ0lP��;���2�%��� �s�}-�7>����;�9S�u�L�4��?��~mʞUJhؘ�?g��{'=����3������i��p�1��$>�C>�d��N&��0�R~K�#�ʭ=��7�&NDZU�{�J�>�֊��PпF�Ĺ�x/!Ů�1j�WaU� �=��+�/N���#<S5�Q�����1�U`�����G��'�o��5>e�\�$$�䈼T�	r��-���/��%v"M���m�F�V6����H�J4��ڊ�j
�Z+S��(�K��J�������?5����D���A{�PT�=�"�}����� <�\sR9��=�RS<�%�0���y/e@�1F��d��L���!���⌞��g6^���k�54ڡ֫�)[gZ�K6Ìv���'&.�&b��v�� ?� �3º�ytSɄ��5k��P)��_Uβ}�VVoQX#s�ҀzK��x�V�@C�=��k��	�D�l/��^a'�@W��PX�y�[�j�� ��U_��<r�����w����7I Ϻ�y7�X��_�nʌ�˝�X�Ǿ��/@�8(���xv]�$V\Gu��;�1�
�y��h$�.H̃��7D���ׇ�,���I�G�1�c�p���{7|w�$V�n8�a��0�&�3�:��Hm{�� 3�JJ���0�i���2{
��&:��o�Ylw�nC��C��&��_�u
�!�3'�:�*V���=9Atǭp˵o�ں�h|�÷��'S(���6���L����u�@���s7wws��1zoXUo���%kP2��t�<cC�3��a8��c�`NCq?��l�î�/������#��t즐��Q�%�2���m����!����1 M�6�ݽ�Ʈ+,nzYaATL���\���z}>�>�!�����ͦ�]�B%e+f5�5@�25�ţ�0��5}!�ԗ��,W����ϭ!�45D��M����]vb;�-��i��a�Er\^Ԥ
b!�~��N����zĻ�4�We�|�a?���+-W�<Q_K���@8 �S��^����w��0�'�EO��G{�JW�N7�ˑ�x���c#�*Ц��]c��;���;���%��2Ɇ,{��I\��*y!����+���shtT��V$�'I6s	h�]fx�m��qLP�Ξ���&Y)��\��f3�J�#|�I�?���/�M��+�lJW�Gm�F�Uw�WG����V2P����,��i�%�ze��D]��F�tb���{)�WMP����o�x���Gt��V2��j���g�V+�]��DD�@��$�c�;�J���{�]���ő^��D���eN����?�# y��$�H��W�/!Rk_i��@z�m��ʧ�H�Q�r�;��$��e�ӌ�d��%8;��PHg����*o�|�ə�m5>�ʺ�C�D!*�S9M?�K!��(���~@#mn=�N\��
��ή�׳�I�C��;ũ��G��w�W�q&�_U���2\M�;}�G�0�&!|.{�v�/'r�a�SNC9P��i4�jߋ���I�²w��� �y�Z;[>S6W>��՝ #!������n�?�h��}A�=��V�,��|���i	'�l����5?��̍-��.����gs�Q��W��&�'��iP"��&��xєA�2i
���)�9��r/�����<�D�v�k�j���*��y�7�������3o�Rd�@�[�'t[�
�u��	����7��[��27�]� ��x�,@|�Z�~|�jn6�F���� �׼G��&ɜ����UJ� �Tϗ�_�|�O[���w�"��;j�F��:�u��c5��_�����o9(�	�g�(�k���6O��4�5���mu����H3��f;��smXpϳd��8�J5��ɔ'��yx������+;���G���8��3Gu����F:^>����n}��A��0���}�_y(:̈�]�F5?[�Ɩ��3(6�cJ�S�(��	W2�n�;\�KX@�M��t��Fts�_��~�#-:x�G��1������|X��瓌l�Q���6fi=GM����n��P#=^*T�����%��x�J�_�0X�07��#�����<�Ӳ��&��Ҁ�n��z��,۾E~Z?��������"}M'�$��x���4{RԼ4H�UꙂ)=�E�����m.�]�"I��\����t�*q���}���%<��6���ECmQ:n���"X}����(�Q{��W(���=xS�4|D�ۖ��G[z��m�`���t�\�B̽�ԱB�) F�GAq��m�oGYę��\��H�!��P祃f��j93>��i5�٤��=��#�x]���	�<�@sq{�΃�Y;W0c�F��,�Ά�'�#'�+�"��@�� �n���tv	��L8�w�������)�����K?�����U�!��@���Y!���&�� ��i�\��+�('lCuv}��ʑI�{({OC�/%/�-Յ���V�O�%`��?7���]��>�y�ǴD��/z�v�*��2_�Z�	���IN��M
!\L�܊�X��jg{�~40��{3��S�4��u1�Ձ<c,){Dq�a�w�6/��3������X=�f�x��ɻe:'�>�hfr׋XM>�HEi0xQ5ƚѢ�`�S��������H'k��*5'�NR��	���� �)�,ϼ.�:�-T�.b:H����2N%F��B�}������Pz	�	 �@��Ne�N�y�y�"ì�y�����y���G�`��k�x��r��!M���ϓF�Teh�7�<e�U��u��_{�F��QL�t~��1x!`�c���t��������h������u���̎�(�?R�y�GJ�/�c�(J�����YѳN��m�<[�=�^:�պ:/c�`;���+SN��H>���T��h>�����IE�6�W6Uh�bW�#CT
�%�](�/ ��H ��^�&���^�6�$��dǊ龠
OB}����0�4褼S�^�n���`2/\d�-~�\Ňiy�y"}���(�\�-oك����3��o͙�]�u��h���olJ6�Y�J��$mY�8h���P�Vibzs*2�����ѹLOА�(�^�4����A=�o��rU�^o������2<�y���0⓴�3^3ɡ����GK�|��Χ��{1T.��S�/��=�aw`PxUгc?�`�W+;���
X�V�j*��@f93�
�f��O��)>#�`�d~�y&Z{�y04�:��tTNm�.�Q��x�O:-�<�sK���%:�%��u��.%O��e��X�<[������(�.�-�U&���_2j��LK�iB5�$�ELG;L�b&��4��6NnFό'�|뾃w����w��ɵ�{-4� ���������d�-�s��9�i�򺫌Ʌ���P �qX���e 5���K;p�}�\�V�ƚ`��2t�M��ǥ�A����~���s��b�s<��o�ڼ?I�2��5{�[.�hZ��y,��h�2�U-~lg#�%�'�f,�L�y�L��FHRow��<t��jޙ�`���@���@��(�Q�=�p����&]�rʖ��j�*��a~�r�<�H��s�H�~�p�v�ӣ��Eʩ�-g1N!�v�
�;N�ɐ��ؔ���G��������#���6r�+G.�7�Τ5Hm8��#�8HH���|�龀�Mw��s��Yx5IJ�P�л�?}��"li�Y�hc��p<]XJ8�XǼ|-2�b8��$N���<iD�.�����b4����1����	�Z^�U��bu�6F�#)�G,�U9�B�)-/��7�Vdu)������5I�����B��L!G�����8��j��P�������K^�x��G«G��&�M|���[(�LDB�U
s��r�~7�t�|`@i��� ΂[$�7r� ׾��fo�g���+j#L��F�=�p���	�߸����E��������J������dw
Pwg�+&���ɱ������5�� S:���$��Rz�-�&�����f�n�D�Ԋ�BBQ:yP���d'��H�Y\�*���������i�a��2�1ϩZv5K5c���M.��,�4��E��<1<��S"��r#�Ē��8�ܜ���;��>o���|,Vm�L�srxT��Ğ�����ƺi��2����SFh:uw�-d�iһTZ�2�l�
>��?Jޗ� }�1��o�D��wŰ�����\��B���yW�R��IJʗ`��\�-�BPߑ�_e���z�S�҇i&�+���<yQ-���/^�ei�õ.X�N����	W��N6K�[� ���?X�Fk��Dm�i��"� ���d/��Y��[�����7���k�L䷱km3�7�i< �B2=G�6�������@~�5%l)9���S[���F �H�E�X;$��D<�Ȫ���0Gx1�20�ǅB�������{@�ClB���Iz�v�������s�"��a��{ ��9h�L�� �亠������7��:$_�-��Fl�	6)�_���]�Uw:�7G��qul�s�`*ų1���6@���1�W��L�VCbkj�*��oʀ���X�s0C(���x� psU�-�J�,�r�6�<3 q����5�Gj���9��fsZB��Z�'^ � w�n���i[aV�lO������YD���b��!�_��{����{���xI�[�i^s�ܪ=l�0F��	̗֦��#6ƈ���OD;|慢�ۥ�%4$ն�:��5A��]��?c^Vٺ�݃�y�������Ёb]�ѕ������I�q��+:���+ZLlS��q{+r�..`�TyuWܷ���!bx�PQ��ٟ1:��c�&L�g@q�Ib�D;���S֓my��X�b�����/]Ql[���QL���,�f�-~�[�>��q��i�����ZJ������$��aO��߁�z����>��/R&�dI����b�xQ'�3K5&C��=�������=�Y��3ͬİ�r��J?�Z��3K�^j�p,DI��I9����Lw�G��':���sp*R��`=n䟲i/�m�`����$$������V�I��d��c��^�(5�d�_~2��w�g�2k���,	���!��*�|$̷1<~�r�	����_���X���)a�#�7���/�<�HM4���ث����IIH�����v�T�!��vB%�͹m  K�H8�N�脕��"��5e<^��h��-ZB�C�ewb�?>A!��!��N�6*.l���d{���n��C�`i�Ж�=��Aa������`>f��،v髭�!Ue@T$�uO�����qg(q[��J�)krt;y��7��)��o�BmƎ/�'>?7�n(�����%�oB:p�?4� �DoK�9�K�.��u@>wC��g�y}7�L/o���q�S���p��)+k��.[���j]�>��y+�Z��������[��0D\-8Z�/�I(#�9�#$��R����"��%��Q���x�.�� ؚa`�ΑC�-#A�`XP�ȵbR��[M
����c�#�j��4�H��Hv��4Ͷ���}���X�V���9��9��ma��V�#��NɎ�����Q�o� ��=w��~y�}t�\��H`+N���·�f�az��Ŋ3X�W!�q~zł=�����-������7���3�C=.���$�mQ�C�Ȟi$\��W��<��V�u፱�
�	�����Pc"Y|X�#����Ep���t{*� ~!�ۥ�E���2K:�r����!�D�tU�����KU��h�0��-���/2e��7rQZ�/��ǰ`,����&�?�-^�̍���Pkt��@�W���X���66��<��t��mc�;�4�W��Q�9��C��0&�g🖤XM�A9�7Y2yۋ*���,1���\"I�G�����ij�B�:��4�+^]�2�C-�u��pI���V0Ϗo���<uz��_�O�W��jzsnL�j@x��|eN�+}�,t"޹���*D��b�rm���(���ߤ�M� ���H{�w��3�/I�O��	3��B�\�4�n�7Ew�t�YR�ˋ�Y�S��7�1���&/0{N�qÅ�Ԓ��VdQ��o0{�����V��`L:�ֿ���٤��k�1��c9y;���H�����õ�1�rs ����[2�IDN��R�1�6�*uϻ��rk��`OIKO��.�`i��Ќτ"t+�!�����#�n_Q��f$���er��C�O�T�ב�2MPHU�38M�?���"WE��l���XJ2��T�&���oDt��tx`*p֏: 1-s+�!Q���+�5��Q���ȏ7˗�k$��}��"{LA���6K[V^�q���z�ڵ��!��+O�T���U��2�핒m��ː3C��i�r�3T�VM|�,:���.�� ���`yec&W���6DgN4�qR�q��:���<����N.o�_�FM?'A?v�҅�;�#��5!46Y��U����e;*P�&;�B6C��'14����gA�_����xR(b|�S
�|s�Ό�U����ϙ
���[��>�l�S��hart����u���#��B���f���J�O��z6� H�b
B�ס� �C�v��\��-~�M����3<נ3��>
�y��_'�)��t����J�8`љq��D�2��+^�Jk��T�V�@��V������q����;��yQ��iA��~M�L̯O�~�q��2�s��i�=���ޞP�Z?�Z��40�����靴
\���gyR}�sm��8��4�ɒ�ǛO*�����9�c���������;���V4��ؽ�J��8��������1e�E�A\A�GOA��L9�e.�)�@�"�h�f�Ţx�<���.o�Ż��"��͗Dӑm�,Gc�����P��T#xǬ����o[�S�
�`�t��)��@�J�����u��F�b���-`��0��Њ��	Fb4��D�wp>��kc�旅���f�=�2��y!�����ߠ�gQj�������iB�c2\�15h���S���k6�V�_]Y?�6�rzٰUY�i*�A���Fk��9�US�O ��tM�4R~K�S;I������
�Ca�~v6�o�4�0V��Aj��g+�
hIr�漣�h���	�߱��
���Ʈr��_�؜�Z9� t�7���гc׍4�E�P���<-���b�{#H�&,�u���+	��RX�\D�tU���Q�x�6�D�"5O�p�}Q׹��Y�z .^A!���/{R���B�����&#�_�����)S쳳a��>t�EC���!r���6�,���1�#N�������.��>�1��5��읻՜@jn�C�d�L������[m��Z�qE;!���'��iĸ]��DݥPw���b�u�(�~͆���Ôo���.�`��~��b�#`��qja�_��K/(���Vf�'�i�1��J�aG�cW`+�Cq
���G�U��s_�W/0��r��z���Z���'o� ���ݨ��O��Ln��$����a$��Z��Qҏ���8�!\�a�7~��Hm��{���gY<WXje�*'�5��ᶤ'M'��H��ЏH�~���:V��zڔ�i,��~�-9���x> .��VV J�ʤd���fz�Ϫl��A�G���}�z"~��t��K�v*��k�#�,1#�[�S�f�xi���4��(��s�8��Z�_�m��1>rb������ݚ3,�s]��͛���)y����&O	?!M�}��>4:lk�C���{0�P�|��~�5��]�/��y���Y��-7�7$%�Z/�V�)�z�G�m�e�"�1��w9�q�'\��w����K�}V�)������%�4��LJ>�c�I���w�d�yY,��;��?fu^+�"$�>�6?���U:@M/����1&�J2�Ggd����蘢�@C�,�\5wj3*qO�z6�JA�t>�G
��d��w�M����ݪ�U'�@ܕ�^ �ZQkX!G�`v�;L���O-�����	���A���!vd� �I\���3 q
i��l��/�; ��"v�D}�� 1-��ݙЏ<`\9�4U�a�;ua��>O�$bC2�l��g�9e����Ms��)�m���	NA���tF�c���z2Tl#1�|��㤮�!Ĕ�v_4^��s�1���.�D�����t�B�F���s�����W�j�C!Kr�8��{��ӣ.��L=�EqrI�|�6��및�`=�iV�E���V��OhT9@Yz'u�!_�:Nn*Wؔ�db� ���:	��qZ��$&Lל�83�T<�T��\�
W�Pl�e�~���_ j:?D"�����g��?�C��{��Nٙv'MBM�g����f�D�f���YROTZ�E�4�4+�����OD��-KT^���Ǔ"X:LPJ�ݛy��=�R֣���ILW
������D�������d��g��fRi��������;�4P8�8��x;G�f����k%q���s�8eɶ��-:������qc�s|,Y#9�ĸn=��D�ap��M��2����,d�on�뙶H��t�
N�P���Q��Gf�炃��cs��Q}r#��{j�:�/�Q�E~�-����(0W^ձN���2萈y�cO"�>5�l���j����&/��jF;m�mC�2bHThe^�8��[a�P���K�F�X�nJu=�7�ƈ�7�y2� �^�F�}g���3)�m(��?�C����7��*�?�̥���cpXQ�1�)�����d5{�*lQ}����rfV��b�s�O�r�R�MR7y�|�Lh�Ju��-Ð{QX���[$s%mwP�A�52:C�ͻ�]sO�Ǝ��+Ǡ���|~t&�L-gQlol���"���̨�m�b<���)ޚ�͓�)��C��],I6$�;����[���w��o�iu������R�yG����b���T6���9�mE�10��H��K�F�eG�,�V�-�Y��Y}�rX���>hP)��Ү�{H�?2Zyo^��$�U�>|��7-_ݺԤn?�V�����i)HǞU�&G�"B��X�A{�Q�bv�bMܮ�X���aG�L����E5j�Ss����΄Xkߓ�yx�I1NC�i�[f-�J?�%�	�m�kLJ.���jz6��P0�̃O?P��-n;=U�������Vq� �A���Sg�N�aA�3��-)�%j_"��%�Y�s7�DD �+��y�����C
_��*K~h��`�zCY�PQ�W�&G�
z��p�N��c�i���&���^��C{{3y���NDdf+1���I|�v8{�ł䕫}[ˊ���5��)�� �	 L��ޝ0������G���!�
PX�삡2	`�5[l�~l8�DK��O-�0�&��#�����]r<��sV���CI�o\U垬E�ZȪ�(��}���}n'�%�+�L6�[��1��Ū"'����}č!��`X�ef5�{��]�6�M�se��IB\� ^P݇�#R��:�L�b*�˒��)�%W���}[È���)CG���:�k-�Uad��f��zW�~�='�c�A�Iɛ��?jW�K#2�wjBʢ�ϥ�
���(���8ZK2N@<,D�rWu�R��b��s`_i�O��>&���@����
���"�c���;�+�3ğ�� ��;��Ov���؍z�l]��az���:ɓ͚t;Za6�;�c_�Hfm�����}N�!w��ս�`|�\t��(���_wԜ��mv������t/N�{ ��C(8˳@���Q}H��&��G����Ye$*�*�Rh��k��w�Fn��6�~�- c�y�ݪz���?��h���x��l�e��W��|���h�3�d��T0{�d(6��-����R�d�ހ��������K���,{D�b�����P=X����Y���Ǉ3�Vh!"�RI��R��Mv�U0�*�C��?��36YI�2 )�� 5�e��`|���'O1�SNl�� 뉥���K ya_7ę
I�:����e��3,5�����%G��J�KvK{	\	s��S��/��,jg�/�R�=^HZ�o��[?�8r�;��KN�Fx��g8����6�ؠ!x]���h!��@5e�S���e�m;�n�9I�G��3*=�`a������V0����kU��,��v�n��@�E`}S��y�O��{�}�K|<�J����<��b֝�l��u/����c�E�5HN�	/K�n9�Es|X:��*0$�6�	�x�b��˯���"%q	��܇0< � �)<}O�a�4箟�G�%
F�A�������D�(8/)^Osްl�"�4&W�ˁͲ=��|�4ꈫB���~�γµ���������H�4��B�,��������J��zD�
�`����ډ{��`��M
��_T&���t����1Ie���*�Lt5:��n	xV�ة$H�k��]��(���M6X�#b�<e�A1�$�� H�WwV����gA�WabF�؊�Է,V���_^�����7답��'�x�~f�e���{�uWn�� ���+���EH�!�W�/*=e�� ���Ja�x�^V��D���Э|J����A^�@`�o������nfc?����) ~qOJ2�*=�L���p~l;�a��6�,r]^0�A?���G��kncs�E�b��.��x<���l�(h'!��qj�'J�v��$b�N��n��:�w �:^?C`X_�b1Y/Z��������nz?�*��dG�u�?P�Ь~�6r(��n�M$\c� #�ݸ�y��b�ӗ_[�KeȼE99��s����q�"�[�F�PޢtM����Ǚ�K�б�yg�k��N-1? O�Kx�<%���S8��1��{_UXi��J���H���y�N^�=;�{G#�EZ��␶:��?|���D.�,�)�I�PǷ���Ȏ��r���A�cg�祝�7�劯�����uD\��rV��1������#�8��Z{L���-��G�������>��e�r��C�
U�Gy)#V��~�z����݀�w���M����~/d�ك��祐�Y���XJ1.3���8�	��
G]8��v�����t�:s7��e˶��$�j6�����3V��\�4L�t��w`�=�
�JǗP��)�Aa�����M~'=H$P\}�V�#� ��Ly�ؤQ�}�#����T`L����A@��	��o�Կ���ѝ�q��D������O�aP8��$�������zH)D�[/I�o��)P@�-F�B� ;ޔN��p|�r9�O���ll��$���6`2fE��}���JqҳD!��@ԙ�wfX���6U�Ql����p�i�.��c�Ⱒ��ؤ��j��O��4��Q�����h
wLh���N�[2�˰�ʭ��A��J�+���
���
.A��>���+��*g�-�;�]����hBR����N���Q��*������GH%Մ�Ճ%�2��~ͼAE<��F��q���P���mn��l�ʓ���`�R=gk�?3@q����w�(fp��dȰX'�Zӯ5,��W�2M�}��1㸼�\��Z�����t���1��o����;��-X�4Y�1�C��7@���e��#AK�Z9T��ً��00P�$5�C��E��z柛Z��V%!GݔM��_�6�5c���V��^_0f|Uҽ��h��6�3�M�^�h_�{h�lZ}��������\�Ȯ
 m�g/�BӃ+憩4�n����[���:?\q�a�u֋I�PU2�0�F��Q�^�cn?��&xOt�x~�d�YB��gp�9$��9,�����"4h�D��]��*�س��+}��*,��O�"��SvS��m}��<t�z��lC�(��>�&�s��]�E�`��s��'>@�[t��c����d6;��͊����Aĸ�	kՈ�},L����f�~� ڎ:�q�S���I�b"�w�PO4.�����n�� ���;�p>�N@��f⠂1x8��F��/�z�&�9$&I�y2	��9;g!��Z6\��Hl䯩�9�~�%.K���@�q%�1U�h��*;L���(SJN��łS)"W3�!s[8#���0إTp�"��-H'�@�2@�e���lߩ{n6!��\+�� �C�|�$��1`/d!�w-�O�[cWW��@�"�K���ns��5��';���jnb�?]D&l��J��y[������YDD�T]�Mx����i-{ҽ���P��?�}а���3%��^��gy�Z 򿙻w��n�u�;����s��;!6_n�?��Wv�8��"��jK;_��>�&�"�O��82U �h/��p�����Jibʚ��=��ҩ���W�S�ڟ�PDw	�XкXL���N0�ۙ-7?�����A-�oh�\h��ϒ|��6�}X�����ֹ�m	њ)�������K�ϒ��e��������8(��&�N����iԙ|��j��XJ$AH�E�k���S��zx 9gt�C����O#���y�]�"��u��NГ��p�z	� �s�����!�@Avy�D��
��V��'���_��,$���,��<K^�G��n� ���`�5��L�Vfw�0�F�Ɇ���7����*{�So=-8@����Vث
�ɺ$56���gj?�1I4OT��K�Oy3E�G��⬡uzx[hj�+�i���J��}G8��@k��w-�1�A�N�������E�|i�
�rFP�����O�� �WL��]<淧����^���T���+���a{7�}�����G�d��RG�@�!�BFbp#���0��w����e57����PoN^'<��M{@���@�+&ziO}����>\"���#��������t�)���~Tw�N_MڄE�r�󐶍?��s|���R��Q��J̉��5���Q��M�nG��D�W@:�>�� )���+n�j�Z��V +G��Z)ɷ���2���4-�I�!0P+!:�s�ݧ���QN/��@���ffH�l�Ν��{����!��+��1�X*X��!ѩ0�4���	ݭZ���j*�����d4~�qY	�ǌ:vtO�SvT��d��H%ol_�@�&�����j��,�_@�}+�.P�W��3'���L+�ɡ$�A���Q�4�c-F2���L&���k���R3$���Q���C�):utʃ�:����S��dס:־��o	y��F&�Ec������JN�l2���k�"ӛ�<���Cc�g᏾zG��ј��|pͻ���yϗ�	Ӌ��s�Q��]ܽ
%��ݣs:#�� �$T9����H����+f�Bؖ��^7ǹ�UG[X��L����z��\((��yu!ޙ�?�������5̂�;B�4�t8��qˑ!�[Ѵ�"�F2��Fn�I��qcl�??.�E<�g���5H�-6K"A��O� W�L_�f�_�����3k/ELn^kXlY��x�h�
vTg�~�?xd��f��l7>����9�VL���+�]y��6cm��(�С�D�:aD�^�p҇��&M��Z��F��!���s���ç-��F�������|x'��0��K�� ��@��H����*��xn�� ������D_�#2�ۥ�"�N1�*8��'��eV� �;���ہ ��K@���a�*��GJ[^��V2�ƇD3K��`,�'6B^�M\����x��yKU1�]�X-�Ρ��e>(�J�n&�{%�L����D�@=����9�C��X�/k.o������Tw52�R�M딽�8N떆3���9,(v˗�=���[�y#���9������5�%�%9�!�P`��\�D��r��ޒ��>�����k(oz�Cԏ{�*�\����G�ph[C>l�!��G��_��q:��=�uB�N®O���b����b�$>�v��~��c�&���B�sdk���aPIL^cY���>`*�X���QWV�2q �2S��%��~�k␋�40����p��`���k��4Q�Es\���P/��WI4"�����{0T��!�'��.ݲ ��[I�
�v�	({9>b2G�x~{�cΐ;��DNO��3�c�Vh��LU�N9[�0l*�ǿ`g����Y]������D`G��.�ǰᾪOUÜ<C�d��h�W��/������a6e�帥�e{�{1��DS<��Q��_�������h���m�l_ �ŨN���?�y������_���1C�Wqwf �>�ʑ������)%�V!�|b�S�S���1�[�y\oc?8 �A�)�k�<gq"^�J'԰ـ�ŶV��y�=H�D?8��_C�˻d�r�D�,��9��F��)��K�?���&�.�8�DF�Z�bN�+������B���]�l��g����������:@!E��;��h8�R�Vҋø�^~�xԈn���V�Уao@�NԽR�Y��'	��a4������A`e����e����Vb��甥���4(�=�a"pS�E�L�����=����Ah:�.���YèO��9̺�:�1��d�4�fTW�W��a�	Q'�6.{>�	� .}���%F��UE��7���f��8HS���7=̶�{�c����j�%f׆%���yR3���(�R���z���8�`F�C�V�K��p�Qx�;��|�4H��`[Z�T�Ha�"=�_��۩�'�j6O�u��?�2
#&;�cz���v��4���]�̕C�#��>u�U��8�xp7�d�~h��B�N�L���9�3�o�J:�רu����L�"��#�3���	9�{V3y΂���q�{���`J�E#_}��=�=p�mc�������e:p�a<�6ۈ{{��Y�$����E�a�;7nO6���T@����p��ļ��I߸T%x�B� b�}��c�hФT^� D�^Mu"�P"6���x��̫H�6c'ž���Z;aT�5��M0��0����>�w�h����:-�G��-m��xm����������̀��I�Q�rMo�w�,}�tu�6ڸ���F��ĸ{��/n1��d�� ϭ)�տ��x�Xn�`��7)?5�z�����+{-��m|��}�J��卒*(ΟM%x�`���5�0G��QZ��h�9[���me��?d�zz��^z^>}H�:nI-���K��O�N�6���2�`�(>mX铔�45`����ν/Rh��[j�4䩎�U���T�Fr
?:6fAxw�_��u�Cpmw.��CШ�6'~˚��!�v�9w���p�[_ԬX�v��2B��^%�.��N�vYN�ݚS�ή�&~����b����?e�?�����n�x�G�T��!����Mׄ�g; ����z,��yv��{6�+�C���6������UJ$5H�_�X6��E�Tn��$���7�_"�X�C��}!`Mj4�+��eZ��~�֒�A��|�J*��@*��sȩV�F�g�P�1|�[�Q�7��M���VԺ�0^~�G't��J�jN��חӬ�aw2������N���vWAP52����d&'����ym�>_S�/k���\��C���䯤��L�"7� x48s#��f��Z�AiǜW@���K�tI����Q�K�1'���U�L�#k�,q*��k3L��~	���x�d��z�"�1�0<���Y���T�ٵ<d�&IBQ��0�
i?Atpt�o<�3�S���[b�����v�3�^�� -Mb� "jlE�im��pW ��- ��	C!H�{cn�2C�� �R��ު�"K�=���sK���� ؽU[��<�ϙ��qO?{%��q]� ��3`�3
9�wM��`qnВ�����ZVT`����枊>vf��Gw��R�b=a��
�V�{-6�i^�[�-;�D�����p�yk{���QL}��_�cô�X"M�i�g��H�Uݩ̙�����bAcr�bz�VH�'�dFG�ȫFR�l�ؒ_�T�q���8
��gq����r����S*��+3���1+�T�ꖐ���`��@�~�.��DX�k��%��Ag�d�4z�)�$6��;P%�@�ݮ��+��-���P��'Lf�a�b���֩F@����92x�޴%�߃����~���Bߖe� + ���4CCr��'a�*���BW;��B.vX�����J�͍<7!��nbC��0�+���A������䊐�8�C�2����G�iN�p��cvXCg{�[�\����(gK#�^sogZ*�YДw�qqXn¯Q�-ٌ��S���X�>%3��1��~\03j���Wř��s�dx�^�t�?����F�FX0��,���6"�v����_� ��='�"���ܸ�%)acFI�����vkBR�������f��*��`����W�eqhu �*R7� ��ţ��a�'#�[%�k�h�5Aʈ�ک��prc�b��<�9	l�2��J�X��g�p��]U���k�H�Q<\��o+��p�V#Y5�z��|�9�3e��rPC���5�Z�+��iZn<U<�5�&zt�?ԑ=��}��
��"��n�Ixk]+�$�i���mTA����<�;'S����l��Y� �l_�i�'/,�0��J��z@��g�E�ij%^g���/<q�V=�G
���]`�uTI�VU�ߣ�eڬi`���:�aσ�-��%"���O���9�	fn�]�ԁ��z=��}��#�n��ɱ�_%J	4�P�	8��Oڊ0��  P����,�����Βɢ
M��ܾ&Ol���/�?�;���5��@�֝�_��u�
�95�ir-V��mV�s9�=�O�`��mT"��'}Yԋ�v��Uj�Ŕ#���(YZ�Rby�6�Vr�˙��I������y'�W��މ�ke�,@�*NW�-�p���C��Yz�Q�>O�s��#%�؇�����He���/	{S#��`��r�{G��R����(��l	�'��do�R�}����s5&�Jj���1���YV�dHt���w�q`��>J��;�=�m���V���06o���z���ڞ%���ț;s�h���c ��^���̲��G(�R0/��st�s8R����6�$jJ�خ�����8�v!�fV|�B=	�m�u�#�&��؁(��;5b��W.fkm�F��!����쐿o��ɡ�ѡ3�,��Q�.`V�>x3�5ÿ�Av������\�@~PW����4��gIfۦ�b�[�����b ��2��ZC;��"">��vb;HvFϙ`���ɖ�_BE�����=�%���6��=Iڲ��H����p�����Q�2��&�=a� ��z
�sK�8�ӟ?qB߾�b��7ƞ�9��Z/8����c��<���A�\nW��6���s��܄'����^1#�v �宱j�9�^�k��r�Sa4���P/�����7����KS��N�����ax��=��uMRҐ��W����w�>�7"�	&�U=�C�^ڤڃ�K�Bn��O����&4�����M������3-����F���a�����n��Ɇ7@��׹RŻ��ż��3��Am@�<S1��⇊��d�P#
����Og\a�$Ҍ~3<�x����H�o/��R�Q+���}�c�G���oD7͹g)�'��ه��h�ֹW�$�N�k蛀5�DxYZf�,و��� ��J�y"\m*	�7� ��x<���lԂ��F��4*'k���v���������\���3�+S�&���5��U�扚������u�L��hwV�2qEeLXi�]����1w����u#�ܦ>��b�-��͑��q�S����~(�YA���.�%��*Ģ�y�r����w�E���ii�J�Cק�R�2���?�w#�f�ʐ��m��������=��F��U�L��s�حw
`N�mv��s[껊꿥ֱ�C�F4�*��颇�vUkvH�� �]�c@��t))��+*��k�(�0x~c7N:�!GR/,s��
u1y*�Zc:��>��pĩb���C��:������2a�2�K�-�:!�������,6vB��4C��M�C��O*d��S�5@�G獓�à��.D�tS�sP5��?������JP5W��Wb�(%^�<��Rx|u�4��&��W���*9�����Fic�^�^���u�6�$�XѮ�Y�C<�1��,��ڄE�cz�d:�r?��J�!J'.���<k�)"���5&E�+aY��g��EI8��M�Ѻim��]�<G���	v{c]묍y��u��(u=�ws	�G���2b�� ~�[�C,=�>W��p�&�=�����,D��7�r��Q?0���O�&F��$�~"�ڑC/e����հg~L��w$:��n" �2�S�����l�Sʓ�pN��4�'�ΰv���j����9�|ƀCr�zHRu�����_t�N�q�Rn���]�����n�BE�׈5�R���{;:��md�ܙ_L�wa.78t}x��[Y~�S�o��l���b(Q
1��9{���+U��2���U��7���:̜2{N�G*v�T�9Σ��1v�����I��Փ2�L��d��q2�vU.����F�6�SF	k�{�GsQ��l^y�(ĸ��,�<[g�BT�̉ε:#�!�l�� ���t�]lU������c�s�*�:��#�7�hӶ
P�G?�)o�j�h����V�PГx��u�=1D4ZKU���Q��SV�K�"��2�zkllR�����%Ǔ��w��ٟ^��1o�bCqq�[��thȤ�\����G�=SxWd��يi7$j�4;�sYɉ�l��K	�-�Z�?��qw1�f��-X�~��	���T���C�B�H�Q#����!����n�p{�P�CO��c�YRU(�`��J~?�"
)����i��MV���LB2�-�B������\��eSXT�/O~�&Ɲ_���� :ꗖת��!��rv4��� {�4�
��7�wل��kbA%����I'"�-�p����+�����|vu�l*հ�6% �>�50Y
���Pfa����ԏVJ�T�	�W���Z!O�=�����S���i�ܭ��ğĻ	���wyXj��� VD}<*�M`n��v�m9c��f�������O-YdQ鳱I�}�����!D$9h�+|�,m��yl#Ǿ���KΣ�t]�4	��`e_\�I�2x�eS�	�\��#�#��k�d�im����]:g�HHg����Av��u���&j�9�ݫ3y�6�R�B9��m.�$��v`��0����D<)ܥF��)76{�`i�LN���v0_�Ӷ˙�9�)AC[���]��
�3�L����5�+ޖt�wv(�ow���+��\5�k\judc(g��H-P.�!0ǻwq�P��;��9a��s��v��aק@
A
��w�;�#�j�Ӟi~��,�7��q��6���(ʏ�3V�Lt4�V ��B�FW�B�쮉^ �=��/ִ$<~������8�J�G�K��NYE3�!�� -�����4��;7l`��	��+d��}�"�]�a���A+�DF�]�~F?���ek���A�b��F�p^�Q��%�(G���\��\�24t��ӳC�Cm=|.�J}��bs�����<���uWT�Dqc���=��X�+趟ބ���0�̙��P�\DS����l5�������Ջx��n��{�2l/N�y��mE7��嗎7^����������h���-��}�`���zT. zs(0(�����=�r�����
5�~�c��[�"vtk�q�%��ʧ��1f�!;X���e�O�Λ�ni"r��Z�1y({_%��}�e�~�����X1^��$�(w��}��d�pO}X5(q�g��U<��R~�K~Ӛ��4�ܑ0^�i���y��qC��#��N�j���g�f�ȱM���@�6��U�k��&XB��䏟���ҷ�p�iK�HANM7�}hhWds0�;d�*Ti�\!��������	���L$C%�#�*�ف�"SJ�˶�f,�|��fBQ������.8@��Y�L\�R	�4����r��);�f��g0ç�Q��@��m7��I��y�i+v/-b�p&uT���11���0$�u}��{{R��$��V%9����]��tGz�x����D����u��T�lQ�L-��/��p��b��w	6��d|'6�����7PM�\� ��%��
z- �����m �����r]*J�j�<�,�H�Y�,��`�$���|cvL+�a�M�8���$�������M�����vɤ&�&����q�.�F���_5QpV���1@�]�_�l�gz^w��-�>���@uʆ��"˃��ޱ<?B�#!JWG�%1�j�kol!�j{#e��b��w� U��R�W��|f�2�V���C�9�ݻo��U���8��:"�Ľ'-��F�f�48�db���4�F��9�gƓ�Z� ��m4M�ϝN���h�e��/m�F*�2��r�N�+�؉�P���6� �8JD��e�}t}�M��f�鬩<�7��G��F����T����t㑃#㿍;�f�=vR9<�ʌ�����Yn��-<V��k�(��sJsK���k�9�4�����w�^_"D���Jf/���X�, i���.ɍ��lSƯ����AB�و�V�r��:ӥހ��ף]M�"� �;�	��Rz�9^�I�J"R�sM��*A��'Tg+�6�礭��t�V�I�ն�F�^$:&��]C���dʍE�0|�?��Ŧ ���c�L&C��|A�|��1>����O���x��%hu<p�-���T�w?���Y"F�\Ǉ�#�$$�!0i�N^i�l~�)�$6�x�~�`׈�A����ј�Z���ah��Ve�Ј�%�sH����-�86 �+� �j{�Dʕ������~�^B�wt,8�#�=�·�!��!�3�&�1�S9�dq�Ɏ~�qӫ�u�Oa��������v�y ��uY�e���p��}�>�a<}�	���*�7MlB�n��Q3k�C���lb���||������^5-N@*ڼ��/�Q�=D9�����X�`���+��s_����N]�f�X\�]�s�D�	�mL��E�ᾝ(���ձ��'�� ȕiyG�QCh4\�e[S���9IJ$����0�:<�*d�b 8k��è�(�8	 �]��p�EI���I�G$D�b�]T�ASـ�E+���ގ�=w���џDs^���:��S�R�y`� R	��,Cx�"�tdY1X���.X�le�s�֜�i��C��x(��t�~Ĝ���ύW9����~
�ArJvX ����:e�=������ Bh&�R����Z�B�p.�l��j�l{Ө��\x��aRFeT����6alU�'���2��; �S��1���귣y��(�JX��
�Ƥk�r(/b���+��@�	��E�;z��ld��G�^z�,��k�1� �t'�r V�^>��c;�βUM�ړC���M�����������>h�/�K=�i#H9_b�S'�.�)�Ck~�*#"b}b@O�� �б�:� �V��Ұ�O���NM�F��P�������&��v��L��+@�o�?C	1��X����A��FƐ��K��W���9�#�q7�����{#��ҫ���� �g	�_�N���T��,���u���������N����SD�f¯��?a���SQ�%��9.�K@�+P��L{���/
7�|`bj��H����`�' 5r0�j�d���|;;���08%hun�R~��ʳj2��S���">rff;���-���^�̀��u���S<���Y�|:�$|g�f�1=���3	F*�FFi���8T2�ؤ�9 $���f ��?(�cht��Pk�J�9�5�2h�:y�z��<:�=�t��7N�fޠ�UCLe ����D(���X
�u��c��OQ�GZLI�i�C&�j�2�^�3��_�z��J'�$��1�r��a�ӊ���YfQt���M��"�eΨ�V���0�R� �r����f�I/_G�|��C%��k���y�B�V�����m�P��ɨA�\Wȭ;���<\�VL0<Xw����P�P	�9f���],[�.B�l_ J�	�+�U	�{�&p4�i�q> U2����+��X�:�Zz�Ou�v��n/�eb�g�<��XҪ*��?0��뫖v���ש�n��2J�4�ڷ�:MzWJv!�Ud�KB���f�AM�� ����Z�-���h��Ƒ; �y�>�>6���jӸhs�fZ�Ѿj�{jO���}��F���Ii�b[�L77Ei4/�.&TFJ~���G��=���p�Z`/�!�B�:�e1gC�J,�}v<���r1�Vl>yK#��r�}ʪ�ſ%��w��l�v��YW(��h�+�09��fZ�H1�_����/���S9|S+�cϙ�ح[�'��x�y�!ۿ��0=�]k_��C�(�,,��c�|+E7	�qLKc���PV��L�z\�F(��m����|0�r���#��Kt�A��f<���c;���zۅҢ�3���
��M.P�[�kp��q��8��.=El�i��t�N���wbX�<�Z��������}��+JE�������Gvk_�a�@V�M��B�Ԟ��.�sA�}���pF�qO-�A�X�W;�g/X>�_w��?c�J�謌s�Hc���cʃyK����d]�L��SY	�#�af��6�f�CO)����{��m��t!��U�R�7{�X4�^
��L0��m�����J�4h�e2k����x�f� ��Rk-�
4�~����%3�|=��ȉ��j�D1�_K�P|�8���௤+(م�Fo�a�V�/6��YL_��PMf�Nݺ��X�F�䯣t�1�t��9I���L��QJ�`#�X��-.;=��J��X�I�ߊ--�t+Fr�Hʝ����t����2KJ��)������_���N�ť̍~�G9M���