-- megafunction wizard: %LPM_DIVIDE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_DIVIDE

-- ============================================================
-- File Name: Divide_32Bit.vhd
-- Megafunction Name(s):
--                      LPM_DIVIDE
--
-- Simulation Library Files(s):
--                      lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 23.1std.1 Build 993 05/14/2024 SC Lite Edition
-- ************************************************************


--Copyright (C) 2024  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions
--and other software and tools, and any partner logic
--functions, and any output files from any of the foregoing
--(including device programming or simulation files), and any
--associated documentation or information are expressly subject
--to the terms and conditions of the Intel Program License
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.


LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

LIBRARY lpm;
USE lpm.ALL;

ENTITY Divide_32Bit IS
  PORT
    (
      clock    : IN  std_logic;
      denom    : IN  std_logic_vector (31 DOWNTO 0);
      numer    : IN  std_logic_vector (31 DOWNTO 0);
      quotient : OUT std_logic_vector (31 DOWNTO 0);
      remain   : OUT std_logic_vector (31 DOWNTO 0)
      );
END Divide_32Bit;


ARCHITECTURE SYN OF divide_32bit IS

  SIGNAL sub_wire0 : std_logic_vector (31 DOWNTO 0);
  SIGNAL sub_wire1 : std_logic_vector (31 DOWNTO 0);



  COMPONENT lpm_divide
    GENERIC (
      lpm_drepresentation : string;
      lpm_hint            : string;
      lpm_nrepresentation : string;
      lpm_pipeline        : natural;
      lpm_type            : string;
      lpm_widthd          : natural;
      lpm_widthn          : natural
      );
    PORT (
      clock    : IN  std_logic;
      denom    : IN  std_logic_vector (31 DOWNTO 0);
      numer    : IN  std_logic_vector (31 DOWNTO 0);
      quotient : OUT std_logic_vector (31 DOWNTO 0);
      remain   : OUT std_logic_vector (31 DOWNTO 0)
      );
  END COMPONENT;

BEGIN
  quotient <= sub_wire0(31 DOWNTO 0);
  remain   <= sub_wire1(31 DOWNTO 0);

  LPM_DIVIDE_component : LPM_DIVIDE
    GENERIC MAP (
      lpm_drepresentation => "UNSIGNED",
      lpm_hint            => "LPM_REMAINDERPOSITIVE=TRUE",
      lpm_nrepresentation => "UNSIGNED",
      lpm_pipeline        => 31,
      lpm_type            => "LPM_DIVIDE",
      lpm_widthd          => 32,
      lpm_widthn          => 32
      )
    PORT MAP (
      clock    => clock,
      denom    => denom,
      numer    => numer,
      quotient => sub_wire0,
      remain   => sub_wire1
      );



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
-- Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "-1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "1"
-- Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "LPM_REMAINDERPOSITIVE=TRUE"
-- Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "31"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
-- Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: denom 0 0 32 0 INPUT NODEFVAL "denom[31..0]"
-- Retrieval info: USED_PORT: numer 0 0 32 0 INPUT NODEFVAL "numer[31..0]"
-- Retrieval info: USED_PORT: quotient 0 0 32 0 OUTPUT NODEFVAL "quotient[31..0]"
-- Retrieval info: USED_PORT: remain 0 0 32 0 OUTPUT NODEFVAL "remain[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @denom 0 0 32 0 denom 0 0 32 0
-- Retrieval info: CONNECT: @numer 0 0 32 0 numer 0 0 32 0
-- Retrieval info: CONNECT: quotient 0 0 32 0 @quotient 0 0 32 0
-- Retrieval info: CONNECT: remain 0 0 32 0 @remain 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Divide_32Bit.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Divide_32Bit.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Divide_32Bit.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Divide_32Bit.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Divide_32Bit_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
